-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Oct 8 2025 23:18:15

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "MAIN" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of MAIN
entity MAIN is
port (
    s3_phy : out std_logic;
    il_min_comp2 : in std_logic;
    il_max_comp1 : in std_logic;
    s1_phy : out std_logic;
    reset : in std_logic;
    il_min_comp1 : in std_logic;
    delay_tr_input : in std_logic;
    s4_phy : out std_logic;
    rgb_g : out std_logic;
    start_stop : in std_logic;
    s2_phy : out std_logic;
    rgb_r : out std_logic;
    rgb_b : out std_logic;
    pwm_output : out std_logic;
    il_max_comp2 : in std_logic;
    delay_hc_input : in std_logic);
end MAIN;

-- Architecture of MAIN
-- View name is \INTERFACE\
architecture \INTERFACE\ of MAIN is

signal \N__48353\ : std_logic;
signal \N__48352\ : std_logic;
signal \N__48351\ : std_logic;
signal \N__48342\ : std_logic;
signal \N__48341\ : std_logic;
signal \N__48340\ : std_logic;
signal \N__48333\ : std_logic;
signal \N__48332\ : std_logic;
signal \N__48331\ : std_logic;
signal \N__48324\ : std_logic;
signal \N__48323\ : std_logic;
signal \N__48322\ : std_logic;
signal \N__48315\ : std_logic;
signal \N__48314\ : std_logic;
signal \N__48313\ : std_logic;
signal \N__48306\ : std_logic;
signal \N__48305\ : std_logic;
signal \N__48304\ : std_logic;
signal \N__48297\ : std_logic;
signal \N__48296\ : std_logic;
signal \N__48295\ : std_logic;
signal \N__48288\ : std_logic;
signal \N__48287\ : std_logic;
signal \N__48286\ : std_logic;
signal \N__48279\ : std_logic;
signal \N__48278\ : std_logic;
signal \N__48277\ : std_logic;
signal \N__48270\ : std_logic;
signal \N__48269\ : std_logic;
signal \N__48268\ : std_logic;
signal \N__48261\ : std_logic;
signal \N__48260\ : std_logic;
signal \N__48259\ : std_logic;
signal \N__48252\ : std_logic;
signal \N__48251\ : std_logic;
signal \N__48250\ : std_logic;
signal \N__48243\ : std_logic;
signal \N__48242\ : std_logic;
signal \N__48241\ : std_logic;
signal \N__48224\ : std_logic;
signal \N__48221\ : std_logic;
signal \N__48218\ : std_logic;
signal \N__48215\ : std_logic;
signal \N__48214\ : std_logic;
signal \N__48211\ : std_logic;
signal \N__48208\ : std_logic;
signal \N__48205\ : std_logic;
signal \N__48202\ : std_logic;
signal \N__48197\ : std_logic;
signal \N__48196\ : std_logic;
signal \N__48195\ : std_logic;
signal \N__48192\ : std_logic;
signal \N__48189\ : std_logic;
signal \N__48186\ : std_logic;
signal \N__48185\ : std_logic;
signal \N__48184\ : std_logic;
signal \N__48183\ : std_logic;
signal \N__48182\ : std_logic;
signal \N__48181\ : std_logic;
signal \N__48180\ : std_logic;
signal \N__48179\ : std_logic;
signal \N__48178\ : std_logic;
signal \N__48177\ : std_logic;
signal \N__48176\ : std_logic;
signal \N__48175\ : std_logic;
signal \N__48174\ : std_logic;
signal \N__48173\ : std_logic;
signal \N__48164\ : std_logic;
signal \N__48159\ : std_logic;
signal \N__48158\ : std_logic;
signal \N__48157\ : std_logic;
signal \N__48156\ : std_logic;
signal \N__48155\ : std_logic;
signal \N__48154\ : std_logic;
signal \N__48153\ : std_logic;
signal \N__48150\ : std_logic;
signal \N__48149\ : std_logic;
signal \N__48146\ : std_logic;
signal \N__48145\ : std_logic;
signal \N__48142\ : std_logic;
signal \N__48139\ : std_logic;
signal \N__48126\ : std_logic;
signal \N__48121\ : std_logic;
signal \N__48118\ : std_logic;
signal \N__48115\ : std_logic;
signal \N__48110\ : std_logic;
signal \N__48093\ : std_logic;
signal \N__48088\ : std_logic;
signal \N__48085\ : std_logic;
signal \N__48074\ : std_logic;
signal \N__48073\ : std_logic;
signal \N__48072\ : std_logic;
signal \N__48071\ : std_logic;
signal \N__48068\ : std_logic;
signal \N__48067\ : std_logic;
signal \N__48066\ : std_logic;
signal \N__48065\ : std_logic;
signal \N__48064\ : std_logic;
signal \N__48063\ : std_logic;
signal \N__48062\ : std_logic;
signal \N__48061\ : std_logic;
signal \N__48060\ : std_logic;
signal \N__48059\ : std_logic;
signal \N__48056\ : std_logic;
signal \N__48053\ : std_logic;
signal \N__48050\ : std_logic;
signal \N__48049\ : std_logic;
signal \N__48048\ : std_logic;
signal \N__48047\ : std_logic;
signal \N__48042\ : std_logic;
signal \N__48039\ : std_logic;
signal \N__48036\ : std_logic;
signal \N__48033\ : std_logic;
signal \N__48030\ : std_logic;
signal \N__48029\ : std_logic;
signal \N__48028\ : std_logic;
signal \N__48027\ : std_logic;
signal \N__48026\ : std_logic;
signal \N__48025\ : std_logic;
signal \N__48024\ : std_logic;
signal \N__48015\ : std_logic;
signal \N__48002\ : std_logic;
signal \N__47999\ : std_logic;
signal \N__47998\ : std_logic;
signal \N__47997\ : std_logic;
signal \N__47988\ : std_logic;
signal \N__47983\ : std_logic;
signal \N__47974\ : std_logic;
signal \N__47969\ : std_logic;
signal \N__47966\ : std_logic;
signal \N__47961\ : std_logic;
signal \N__47948\ : std_logic;
signal \N__47947\ : std_logic;
signal \N__47946\ : std_logic;
signal \N__47943\ : std_logic;
signal \N__47942\ : std_logic;
signal \N__47941\ : std_logic;
signal \N__47940\ : std_logic;
signal \N__47937\ : std_logic;
signal \N__47934\ : std_logic;
signal \N__47933\ : std_logic;
signal \N__47930\ : std_logic;
signal \N__47923\ : std_logic;
signal \N__47916\ : std_logic;
signal \N__47915\ : std_logic;
signal \N__47914\ : std_logic;
signal \N__47913\ : std_logic;
signal \N__47912\ : std_logic;
signal \N__47911\ : std_logic;
signal \N__47910\ : std_logic;
signal \N__47903\ : std_logic;
signal \N__47898\ : std_logic;
signal \N__47895\ : std_logic;
signal \N__47894\ : std_logic;
signal \N__47893\ : std_logic;
signal \N__47892\ : std_logic;
signal \N__47891\ : std_logic;
signal \N__47890\ : std_logic;
signal \N__47889\ : std_logic;
signal \N__47888\ : std_logic;
signal \N__47887\ : std_logic;
signal \N__47886\ : std_logic;
signal \N__47879\ : std_logic;
signal \N__47874\ : std_logic;
signal \N__47873\ : std_logic;
signal \N__47872\ : std_logic;
signal \N__47867\ : std_logic;
signal \N__47850\ : std_logic;
signal \N__47845\ : std_logic;
signal \N__47840\ : std_logic;
signal \N__47831\ : std_logic;
signal \N__47828\ : std_logic;
signal \N__47825\ : std_logic;
signal \N__47824\ : std_logic;
signal \N__47821\ : std_logic;
signal \N__47818\ : std_logic;
signal \N__47813\ : std_logic;
signal \N__47810\ : std_logic;
signal \N__47807\ : std_logic;
signal \N__47806\ : std_logic;
signal \N__47803\ : std_logic;
signal \N__47800\ : std_logic;
signal \N__47797\ : std_logic;
signal \N__47794\ : std_logic;
signal \N__47791\ : std_logic;
signal \N__47788\ : std_logic;
signal \N__47783\ : std_logic;
signal \N__47782\ : std_logic;
signal \N__47781\ : std_logic;
signal \N__47780\ : std_logic;
signal \N__47779\ : std_logic;
signal \N__47776\ : std_logic;
signal \N__47773\ : std_logic;
signal \N__47770\ : std_logic;
signal \N__47767\ : std_logic;
signal \N__47764\ : std_logic;
signal \N__47761\ : std_logic;
signal \N__47756\ : std_logic;
signal \N__47753\ : std_logic;
signal \N__47750\ : std_logic;
signal \N__47745\ : std_logic;
signal \N__47742\ : std_logic;
signal \N__47735\ : std_logic;
signal \N__47732\ : std_logic;
signal \N__47729\ : std_logic;
signal \N__47726\ : std_logic;
signal \N__47725\ : std_logic;
signal \N__47724\ : std_logic;
signal \N__47723\ : std_logic;
signal \N__47720\ : std_logic;
signal \N__47713\ : std_logic;
signal \N__47708\ : std_logic;
signal \N__47707\ : std_logic;
signal \N__47706\ : std_logic;
signal \N__47701\ : std_logic;
signal \N__47698\ : std_logic;
signal \N__47695\ : std_logic;
signal \N__47694\ : std_logic;
signal \N__47691\ : std_logic;
signal \N__47688\ : std_logic;
signal \N__47685\ : std_logic;
signal \N__47684\ : std_logic;
signal \N__47681\ : std_logic;
signal \N__47678\ : std_logic;
signal \N__47673\ : std_logic;
signal \N__47666\ : std_logic;
signal \N__47665\ : std_logic;
signal \N__47664\ : std_logic;
signal \N__47663\ : std_logic;
signal \N__47660\ : std_logic;
signal \N__47657\ : std_logic;
signal \N__47652\ : std_logic;
signal \N__47649\ : std_logic;
signal \N__47642\ : std_logic;
signal \N__47641\ : std_logic;
signal \N__47638\ : std_logic;
signal \N__47637\ : std_logic;
signal \N__47634\ : std_logic;
signal \N__47631\ : std_logic;
signal \N__47628\ : std_logic;
signal \N__47625\ : std_logic;
signal \N__47622\ : std_logic;
signal \N__47615\ : std_logic;
signal \N__47612\ : std_logic;
signal \N__47609\ : std_logic;
signal \N__47606\ : std_logic;
signal \N__47605\ : std_logic;
signal \N__47604\ : std_logic;
signal \N__47599\ : std_logic;
signal \N__47598\ : std_logic;
signal \N__47597\ : std_logic;
signal \N__47596\ : std_logic;
signal \N__47595\ : std_logic;
signal \N__47594\ : std_logic;
signal \N__47593\ : std_logic;
signal \N__47590\ : std_logic;
signal \N__47587\ : std_logic;
signal \N__47578\ : std_logic;
signal \N__47573\ : std_logic;
signal \N__47570\ : std_logic;
signal \N__47567\ : std_logic;
signal \N__47564\ : std_logic;
signal \N__47561\ : std_logic;
signal \N__47558\ : std_logic;
signal \N__47555\ : std_logic;
signal \N__47552\ : std_logic;
signal \N__47547\ : std_logic;
signal \N__47540\ : std_logic;
signal \N__47539\ : std_logic;
signal \N__47538\ : std_logic;
signal \N__47537\ : std_logic;
signal \N__47536\ : std_logic;
signal \N__47535\ : std_logic;
signal \N__47534\ : std_logic;
signal \N__47531\ : std_logic;
signal \N__47530\ : std_logic;
signal \N__47527\ : std_logic;
signal \N__47524\ : std_logic;
signal \N__47521\ : std_logic;
signal \N__47520\ : std_logic;
signal \N__47513\ : std_logic;
signal \N__47510\ : std_logic;
signal \N__47507\ : std_logic;
signal \N__47502\ : std_logic;
signal \N__47499\ : std_logic;
signal \N__47496\ : std_logic;
signal \N__47493\ : std_logic;
signal \N__47488\ : std_logic;
signal \N__47487\ : std_logic;
signal \N__47484\ : std_logic;
signal \N__47481\ : std_logic;
signal \N__47478\ : std_logic;
signal \N__47475\ : std_logic;
signal \N__47472\ : std_logic;
signal \N__47469\ : std_logic;
signal \N__47466\ : std_logic;
signal \N__47463\ : std_logic;
signal \N__47456\ : std_logic;
signal \N__47447\ : std_logic;
signal \N__47444\ : std_logic;
signal \N__47443\ : std_logic;
signal \N__47442\ : std_logic;
signal \N__47439\ : std_logic;
signal \N__47436\ : std_logic;
signal \N__47435\ : std_logic;
signal \N__47432\ : std_logic;
signal \N__47429\ : std_logic;
signal \N__47426\ : std_logic;
signal \N__47421\ : std_logic;
signal \N__47418\ : std_logic;
signal \N__47413\ : std_logic;
signal \N__47410\ : std_logic;
signal \N__47407\ : std_logic;
signal \N__47402\ : std_logic;
signal \N__47401\ : std_logic;
signal \N__47400\ : std_logic;
signal \N__47397\ : std_logic;
signal \N__47392\ : std_logic;
signal \N__47391\ : std_logic;
signal \N__47390\ : std_logic;
signal \N__47387\ : std_logic;
signal \N__47384\ : std_logic;
signal \N__47379\ : std_logic;
signal \N__47376\ : std_logic;
signal \N__47371\ : std_logic;
signal \N__47366\ : std_logic;
signal \N__47363\ : std_logic;
signal \N__47360\ : std_logic;
signal \N__47357\ : std_logic;
signal \N__47354\ : std_logic;
signal \N__47351\ : std_logic;
signal \N__47350\ : std_logic;
signal \N__47349\ : std_logic;
signal \N__47348\ : std_logic;
signal \N__47347\ : std_logic;
signal \N__47346\ : std_logic;
signal \N__47345\ : std_logic;
signal \N__47344\ : std_logic;
signal \N__47343\ : std_logic;
signal \N__47342\ : std_logic;
signal \N__47341\ : std_logic;
signal \N__47340\ : std_logic;
signal \N__47339\ : std_logic;
signal \N__47338\ : std_logic;
signal \N__47337\ : std_logic;
signal \N__47336\ : std_logic;
signal \N__47335\ : std_logic;
signal \N__47334\ : std_logic;
signal \N__47333\ : std_logic;
signal \N__47332\ : std_logic;
signal \N__47331\ : std_logic;
signal \N__47330\ : std_logic;
signal \N__47329\ : std_logic;
signal \N__47328\ : std_logic;
signal \N__47327\ : std_logic;
signal \N__47326\ : std_logic;
signal \N__47325\ : std_logic;
signal \N__47324\ : std_logic;
signal \N__47323\ : std_logic;
signal \N__47322\ : std_logic;
signal \N__47321\ : std_logic;
signal \N__47320\ : std_logic;
signal \N__47319\ : std_logic;
signal \N__47318\ : std_logic;
signal \N__47317\ : std_logic;
signal \N__47316\ : std_logic;
signal \N__47315\ : std_logic;
signal \N__47314\ : std_logic;
signal \N__47313\ : std_logic;
signal \N__47312\ : std_logic;
signal \N__47311\ : std_logic;
signal \N__47310\ : std_logic;
signal \N__47309\ : std_logic;
signal \N__47308\ : std_logic;
signal \N__47307\ : std_logic;
signal \N__47306\ : std_logic;
signal \N__47305\ : std_logic;
signal \N__47304\ : std_logic;
signal \N__47303\ : std_logic;
signal \N__47302\ : std_logic;
signal \N__47301\ : std_logic;
signal \N__47300\ : std_logic;
signal \N__47299\ : std_logic;
signal \N__47298\ : std_logic;
signal \N__47297\ : std_logic;
signal \N__47296\ : std_logic;
signal \N__47295\ : std_logic;
signal \N__47294\ : std_logic;
signal \N__47293\ : std_logic;
signal \N__47292\ : std_logic;
signal \N__47291\ : std_logic;
signal \N__47290\ : std_logic;
signal \N__47289\ : std_logic;
signal \N__47288\ : std_logic;
signal \N__47287\ : std_logic;
signal \N__47286\ : std_logic;
signal \N__47285\ : std_logic;
signal \N__47284\ : std_logic;
signal \N__47283\ : std_logic;
signal \N__47282\ : std_logic;
signal \N__47281\ : std_logic;
signal \N__47280\ : std_logic;
signal \N__47279\ : std_logic;
signal \N__47278\ : std_logic;
signal \N__47277\ : std_logic;
signal \N__47276\ : std_logic;
signal \N__47275\ : std_logic;
signal \N__47274\ : std_logic;
signal \N__47273\ : std_logic;
signal \N__47272\ : std_logic;
signal \N__47271\ : std_logic;
signal \N__47270\ : std_logic;
signal \N__47269\ : std_logic;
signal \N__47268\ : std_logic;
signal \N__47267\ : std_logic;
signal \N__47266\ : std_logic;
signal \N__47265\ : std_logic;
signal \N__47264\ : std_logic;
signal \N__47263\ : std_logic;
signal \N__47262\ : std_logic;
signal \N__47261\ : std_logic;
signal \N__47260\ : std_logic;
signal \N__47259\ : std_logic;
signal \N__47258\ : std_logic;
signal \N__47257\ : std_logic;
signal \N__47256\ : std_logic;
signal \N__47255\ : std_logic;
signal \N__47254\ : std_logic;
signal \N__47253\ : std_logic;
signal \N__47252\ : std_logic;
signal \N__47251\ : std_logic;
signal \N__47250\ : std_logic;
signal \N__47249\ : std_logic;
signal \N__47248\ : std_logic;
signal \N__47247\ : std_logic;
signal \N__47246\ : std_logic;
signal \N__47245\ : std_logic;
signal \N__47244\ : std_logic;
signal \N__47243\ : std_logic;
signal \N__47242\ : std_logic;
signal \N__47241\ : std_logic;
signal \N__47240\ : std_logic;
signal \N__47239\ : std_logic;
signal \N__47238\ : std_logic;
signal \N__47237\ : std_logic;
signal \N__47236\ : std_logic;
signal \N__47235\ : std_logic;
signal \N__47234\ : std_logic;
signal \N__47233\ : std_logic;
signal \N__47232\ : std_logic;
signal \N__47231\ : std_logic;
signal \N__47230\ : std_logic;
signal \N__47229\ : std_logic;
signal \N__47228\ : std_logic;
signal \N__47227\ : std_logic;
signal \N__47226\ : std_logic;
signal \N__47225\ : std_logic;
signal \N__47224\ : std_logic;
signal \N__47223\ : std_logic;
signal \N__47222\ : std_logic;
signal \N__47221\ : std_logic;
signal \N__47220\ : std_logic;
signal \N__47219\ : std_logic;
signal \N__47218\ : std_logic;
signal \N__47217\ : std_logic;
signal \N__47216\ : std_logic;
signal \N__47215\ : std_logic;
signal \N__47214\ : std_logic;
signal \N__47213\ : std_logic;
signal \N__47212\ : std_logic;
signal \N__47211\ : std_logic;
signal \N__47210\ : std_logic;
signal \N__47209\ : std_logic;
signal \N__47208\ : std_logic;
signal \N__47207\ : std_logic;
signal \N__47206\ : std_logic;
signal \N__47205\ : std_logic;
signal \N__47204\ : std_logic;
signal \N__47203\ : std_logic;
signal \N__47202\ : std_logic;
signal \N__47201\ : std_logic;
signal \N__47200\ : std_logic;
signal \N__47199\ : std_logic;
signal \N__47198\ : std_logic;
signal \N__47197\ : std_logic;
signal \N__47196\ : std_logic;
signal \N__47195\ : std_logic;
signal \N__47194\ : std_logic;
signal \N__47193\ : std_logic;
signal \N__47192\ : std_logic;
signal \N__47191\ : std_logic;
signal \N__47190\ : std_logic;
signal \N__47189\ : std_logic;
signal \N__46862\ : std_logic;
signal \N__46859\ : std_logic;
signal \N__46858\ : std_logic;
signal \N__46857\ : std_logic;
signal \N__46856\ : std_logic;
signal \N__46853\ : std_logic;
signal \N__46852\ : std_logic;
signal \N__46849\ : std_logic;
signal \N__46846\ : std_logic;
signal \N__46843\ : std_logic;
signal \N__46840\ : std_logic;
signal \N__46837\ : std_logic;
signal \N__46834\ : std_logic;
signal \N__46831\ : std_logic;
signal \N__46828\ : std_logic;
signal \N__46827\ : std_logic;
signal \N__46826\ : std_logic;
signal \N__46823\ : std_logic;
signal \N__46820\ : std_logic;
signal \N__46817\ : std_logic;
signal \N__46812\ : std_logic;
signal \N__46809\ : std_logic;
signal \N__46806\ : std_logic;
signal \N__46801\ : std_logic;
signal \N__46796\ : std_logic;
signal \N__46793\ : std_logic;
signal \N__46790\ : std_logic;
signal \N__46781\ : std_logic;
signal \N__46780\ : std_logic;
signal \N__46779\ : std_logic;
signal \N__46778\ : std_logic;
signal \N__46777\ : std_logic;
signal \N__46774\ : std_logic;
signal \N__46773\ : std_logic;
signal \N__46770\ : std_logic;
signal \N__46767\ : std_logic;
signal \N__46764\ : std_logic;
signal \N__46761\ : std_logic;
signal \N__46758\ : std_logic;
signal \N__46755\ : std_logic;
signal \N__46752\ : std_logic;
signal \N__46749\ : std_logic;
signal \N__46746\ : std_logic;
signal \N__46745\ : std_logic;
signal \N__46744\ : std_logic;
signal \N__46743\ : std_logic;
signal \N__46742\ : std_logic;
signal \N__46741\ : std_logic;
signal \N__46740\ : std_logic;
signal \N__46739\ : std_logic;
signal \N__46738\ : std_logic;
signal \N__46737\ : std_logic;
signal \N__46736\ : std_logic;
signal \N__46735\ : std_logic;
signal \N__46734\ : std_logic;
signal \N__46733\ : std_logic;
signal \N__46732\ : std_logic;
signal \N__46731\ : std_logic;
signal \N__46730\ : std_logic;
signal \N__46729\ : std_logic;
signal \N__46728\ : std_logic;
signal \N__46727\ : std_logic;
signal \N__46726\ : std_logic;
signal \N__46725\ : std_logic;
signal \N__46724\ : std_logic;
signal \N__46723\ : std_logic;
signal \N__46722\ : std_logic;
signal \N__46721\ : std_logic;
signal \N__46720\ : std_logic;
signal \N__46719\ : std_logic;
signal \N__46718\ : std_logic;
signal \N__46717\ : std_logic;
signal \N__46716\ : std_logic;
signal \N__46715\ : std_logic;
signal \N__46714\ : std_logic;
signal \N__46713\ : std_logic;
signal \N__46712\ : std_logic;
signal \N__46711\ : std_logic;
signal \N__46710\ : std_logic;
signal \N__46709\ : std_logic;
signal \N__46708\ : std_logic;
signal \N__46707\ : std_logic;
signal \N__46706\ : std_logic;
signal \N__46705\ : std_logic;
signal \N__46704\ : std_logic;
signal \N__46703\ : std_logic;
signal \N__46702\ : std_logic;
signal \N__46701\ : std_logic;
signal \N__46698\ : std_logic;
signal \N__46697\ : std_logic;
signal \N__46696\ : std_logic;
signal \N__46695\ : std_logic;
signal \N__46694\ : std_logic;
signal \N__46693\ : std_logic;
signal \N__46692\ : std_logic;
signal \N__46691\ : std_logic;
signal \N__46690\ : std_logic;
signal \N__46689\ : std_logic;
signal \N__46688\ : std_logic;
signal \N__46687\ : std_logic;
signal \N__46686\ : std_logic;
signal \N__46685\ : std_logic;
signal \N__46684\ : std_logic;
signal \N__46683\ : std_logic;
signal \N__46682\ : std_logic;
signal \N__46681\ : std_logic;
signal \N__46680\ : std_logic;
signal \N__46679\ : std_logic;
signal \N__46678\ : std_logic;
signal \N__46677\ : std_logic;
signal \N__46676\ : std_logic;
signal \N__46675\ : std_logic;
signal \N__46674\ : std_logic;
signal \N__46673\ : std_logic;
signal \N__46672\ : std_logic;
signal \N__46671\ : std_logic;
signal \N__46670\ : std_logic;
signal \N__46669\ : std_logic;
signal \N__46668\ : std_logic;
signal \N__46667\ : std_logic;
signal \N__46666\ : std_logic;
signal \N__46665\ : std_logic;
signal \N__46664\ : std_logic;
signal \N__46663\ : std_logic;
signal \N__46662\ : std_logic;
signal \N__46661\ : std_logic;
signal \N__46660\ : std_logic;
signal \N__46659\ : std_logic;
signal \N__46658\ : std_logic;
signal \N__46657\ : std_logic;
signal \N__46656\ : std_logic;
signal \N__46655\ : std_logic;
signal \N__46654\ : std_logic;
signal \N__46653\ : std_logic;
signal \N__46652\ : std_logic;
signal \N__46651\ : std_logic;
signal \N__46650\ : std_logic;
signal \N__46649\ : std_logic;
signal \N__46648\ : std_logic;
signal \N__46647\ : std_logic;
signal \N__46646\ : std_logic;
signal \N__46645\ : std_logic;
signal \N__46644\ : std_logic;
signal \N__46643\ : std_logic;
signal \N__46642\ : std_logic;
signal \N__46641\ : std_logic;
signal \N__46640\ : std_logic;
signal \N__46639\ : std_logic;
signal \N__46638\ : std_logic;
signal \N__46637\ : std_logic;
signal \N__46636\ : std_logic;
signal \N__46635\ : std_logic;
signal \N__46634\ : std_logic;
signal \N__46633\ : std_logic;
signal \N__46632\ : std_logic;
signal \N__46631\ : std_logic;
signal \N__46630\ : std_logic;
signal \N__46629\ : std_logic;
signal \N__46628\ : std_logic;
signal \N__46627\ : std_logic;
signal \N__46624\ : std_logic;
signal \N__46621\ : std_logic;
signal \N__46620\ : std_logic;
signal \N__46619\ : std_logic;
signal \N__46618\ : std_logic;
signal \N__46617\ : std_logic;
signal \N__46616\ : std_logic;
signal \N__46615\ : std_logic;
signal \N__46614\ : std_logic;
signal \N__46613\ : std_logic;
signal \N__46612\ : std_logic;
signal \N__46611\ : std_logic;
signal \N__46610\ : std_logic;
signal \N__46609\ : std_logic;
signal \N__46608\ : std_logic;
signal \N__46607\ : std_logic;
signal \N__46606\ : std_logic;
signal \N__46605\ : std_logic;
signal \N__46604\ : std_logic;
signal \N__46603\ : std_logic;
signal \N__46602\ : std_logic;
signal \N__46601\ : std_logic;
signal \N__46600\ : std_logic;
signal \N__46599\ : std_logic;
signal \N__46598\ : std_logic;
signal \N__46597\ : std_logic;
signal \N__46596\ : std_logic;
signal \N__46595\ : std_logic;
signal \N__46298\ : std_logic;
signal \N__46295\ : std_logic;
signal \N__46292\ : std_logic;
signal \N__46291\ : std_logic;
signal \N__46288\ : std_logic;
signal \N__46285\ : std_logic;
signal \N__46280\ : std_logic;
signal \N__46277\ : std_logic;
signal \N__46274\ : std_logic;
signal \N__46271\ : std_logic;
signal \N__46270\ : std_logic;
signal \N__46267\ : std_logic;
signal \N__46264\ : std_logic;
signal \N__46259\ : std_logic;
signal \N__46256\ : std_logic;
signal \N__46253\ : std_logic;
signal \N__46250\ : std_logic;
signal \N__46249\ : std_logic;
signal \N__46246\ : std_logic;
signal \N__46243\ : std_logic;
signal \N__46238\ : std_logic;
signal \N__46235\ : std_logic;
signal \N__46232\ : std_logic;
signal \N__46229\ : std_logic;
signal \N__46226\ : std_logic;
signal \N__46225\ : std_logic;
signal \N__46222\ : std_logic;
signal \N__46219\ : std_logic;
signal \N__46214\ : std_logic;
signal \N__46211\ : std_logic;
signal \N__46208\ : std_logic;
signal \N__46205\ : std_logic;
signal \N__46202\ : std_logic;
signal \N__46201\ : std_logic;
signal \N__46198\ : std_logic;
signal \N__46195\ : std_logic;
signal \N__46192\ : std_logic;
signal \N__46187\ : std_logic;
signal \N__46184\ : std_logic;
signal \N__46181\ : std_logic;
signal \N__46178\ : std_logic;
signal \N__46177\ : std_logic;
signal \N__46174\ : std_logic;
signal \N__46171\ : std_logic;
signal \N__46166\ : std_logic;
signal \N__46163\ : std_logic;
signal \N__46160\ : std_logic;
signal \N__46157\ : std_logic;
signal \N__46156\ : std_logic;
signal \N__46153\ : std_logic;
signal \N__46150\ : std_logic;
signal \N__46145\ : std_logic;
signal \N__46142\ : std_logic;
signal \N__46139\ : std_logic;
signal \N__46136\ : std_logic;
signal \N__46135\ : std_logic;
signal \N__46132\ : std_logic;
signal \N__46129\ : std_logic;
signal \N__46124\ : std_logic;
signal \N__46121\ : std_logic;
signal \N__46118\ : std_logic;
signal \N__46115\ : std_logic;
signal \N__46112\ : std_logic;
signal \N__46111\ : std_logic;
signal \N__46108\ : std_logic;
signal \N__46105\ : std_logic;
signal \N__46100\ : std_logic;
signal \N__46097\ : std_logic;
signal \N__46094\ : std_logic;
signal \N__46091\ : std_logic;
signal \N__46090\ : std_logic;
signal \N__46087\ : std_logic;
signal \N__46084\ : std_logic;
signal \N__46079\ : std_logic;
signal \N__46076\ : std_logic;
signal \N__46073\ : std_logic;
signal \N__46070\ : std_logic;
signal \N__46069\ : std_logic;
signal \N__46066\ : std_logic;
signal \N__46063\ : std_logic;
signal \N__46058\ : std_logic;
signal \N__46055\ : std_logic;
signal \N__46052\ : std_logic;
signal \N__46049\ : std_logic;
signal \N__46048\ : std_logic;
signal \N__46045\ : std_logic;
signal \N__46042\ : std_logic;
signal \N__46037\ : std_logic;
signal \N__46034\ : std_logic;
signal \N__46031\ : std_logic;
signal \N__46028\ : std_logic;
signal \N__46027\ : std_logic;
signal \N__46024\ : std_logic;
signal \N__46021\ : std_logic;
signal \N__46016\ : std_logic;
signal \N__46013\ : std_logic;
signal \N__46010\ : std_logic;
signal \N__46007\ : std_logic;
signal \N__46004\ : std_logic;
signal \N__46003\ : std_logic;
signal \N__46000\ : std_logic;
signal \N__45997\ : std_logic;
signal \N__45992\ : std_logic;
signal \N__45989\ : std_logic;
signal \N__45986\ : std_logic;
signal \N__45983\ : std_logic;
signal \N__45982\ : std_logic;
signal \N__45979\ : std_logic;
signal \N__45976\ : std_logic;
signal \N__45971\ : std_logic;
signal \N__45968\ : std_logic;
signal \N__45965\ : std_logic;
signal \N__45962\ : std_logic;
signal \N__45959\ : std_logic;
signal \N__45958\ : std_logic;
signal \N__45955\ : std_logic;
signal \N__45954\ : std_logic;
signal \N__45951\ : std_logic;
signal \N__45948\ : std_logic;
signal \N__45945\ : std_logic;
signal \N__45942\ : std_logic;
signal \N__45935\ : std_logic;
signal \N__45932\ : std_logic;
signal \N__45929\ : std_logic;
signal \N__45926\ : std_logic;
signal \N__45923\ : std_logic;
signal \N__45920\ : std_logic;
signal \N__45917\ : std_logic;
signal \N__45914\ : std_logic;
signal \N__45913\ : std_logic;
signal \N__45910\ : std_logic;
signal \N__45907\ : std_logic;
signal \N__45904\ : std_logic;
signal \N__45899\ : std_logic;
signal \N__45898\ : std_logic;
signal \N__45895\ : std_logic;
signal \N__45892\ : std_logic;
signal \N__45891\ : std_logic;
signal \N__45886\ : std_logic;
signal \N__45883\ : std_logic;
signal \N__45880\ : std_logic;
signal \N__45875\ : std_logic;
signal \N__45872\ : std_logic;
signal \N__45869\ : std_logic;
signal \N__45866\ : std_logic;
signal \N__45863\ : std_logic;
signal \N__45860\ : std_logic;
signal \N__45859\ : std_logic;
signal \N__45856\ : std_logic;
signal \N__45853\ : std_logic;
signal \N__45850\ : std_logic;
signal \N__45845\ : std_logic;
signal \N__45844\ : std_logic;
signal \N__45841\ : std_logic;
signal \N__45838\ : std_logic;
signal \N__45837\ : std_logic;
signal \N__45832\ : std_logic;
signal \N__45829\ : std_logic;
signal \N__45826\ : std_logic;
signal \N__45821\ : std_logic;
signal \N__45818\ : std_logic;
signal \N__45815\ : std_logic;
signal \N__45812\ : std_logic;
signal \N__45809\ : std_logic;
signal \N__45806\ : std_logic;
signal \N__45803\ : std_logic;
signal \N__45802\ : std_logic;
signal \N__45801\ : std_logic;
signal \N__45798\ : std_logic;
signal \N__45797\ : std_logic;
signal \N__45796\ : std_logic;
signal \N__45795\ : std_logic;
signal \N__45794\ : std_logic;
signal \N__45791\ : std_logic;
signal \N__45790\ : std_logic;
signal \N__45787\ : std_logic;
signal \N__45786\ : std_logic;
signal \N__45785\ : std_logic;
signal \N__45782\ : std_logic;
signal \N__45773\ : std_logic;
signal \N__45770\ : std_logic;
signal \N__45765\ : std_logic;
signal \N__45762\ : std_logic;
signal \N__45761\ : std_logic;
signal \N__45760\ : std_logic;
signal \N__45757\ : std_logic;
signal \N__45748\ : std_logic;
signal \N__45741\ : std_logic;
signal \N__45736\ : std_logic;
signal \N__45731\ : std_logic;
signal \N__45728\ : std_logic;
signal \N__45727\ : std_logic;
signal \N__45726\ : std_logic;
signal \N__45725\ : std_logic;
signal \N__45722\ : std_logic;
signal \N__45719\ : std_logic;
signal \N__45718\ : std_logic;
signal \N__45715\ : std_logic;
signal \N__45712\ : std_logic;
signal \N__45707\ : std_logic;
signal \N__45704\ : std_logic;
signal \N__45703\ : std_logic;
signal \N__45698\ : std_logic;
signal \N__45693\ : std_logic;
signal \N__45690\ : std_logic;
signal \N__45687\ : std_logic;
signal \N__45684\ : std_logic;
signal \N__45681\ : std_logic;
signal \N__45674\ : std_logic;
signal \N__45671\ : std_logic;
signal \N__45668\ : std_logic;
signal \N__45665\ : std_logic;
signal \N__45664\ : std_logic;
signal \N__45661\ : std_logic;
signal \N__45660\ : std_logic;
signal \N__45657\ : std_logic;
signal \N__45654\ : std_logic;
signal \N__45651\ : std_logic;
signal \N__45644\ : std_logic;
signal \N__45643\ : std_logic;
signal \N__45640\ : std_logic;
signal \N__45637\ : std_logic;
signal \N__45632\ : std_logic;
signal \N__45629\ : std_logic;
signal \N__45626\ : std_logic;
signal \N__45623\ : std_logic;
signal \N__45620\ : std_logic;
signal \N__45617\ : std_logic;
signal \N__45614\ : std_logic;
signal \N__45611\ : std_logic;
signal \N__45610\ : std_logic;
signal \N__45607\ : std_logic;
signal \N__45604\ : std_logic;
signal \N__45599\ : std_logic;
signal \N__45596\ : std_logic;
signal \N__45593\ : std_logic;
signal \N__45590\ : std_logic;
signal \N__45587\ : std_logic;
signal \N__45584\ : std_logic;
signal \N__45583\ : std_logic;
signal \N__45580\ : std_logic;
signal \N__45579\ : std_logic;
signal \N__45576\ : std_logic;
signal \N__45573\ : std_logic;
signal \N__45570\ : std_logic;
signal \N__45563\ : std_logic;
signal \N__45560\ : std_logic;
signal \N__45557\ : std_logic;
signal \N__45554\ : std_logic;
signal \N__45551\ : std_logic;
signal \N__45548\ : std_logic;
signal \N__45547\ : std_logic;
signal \N__45544\ : std_logic;
signal \N__45541\ : std_logic;
signal \N__45538\ : std_logic;
signal \N__45537\ : std_logic;
signal \N__45534\ : std_logic;
signal \N__45531\ : std_logic;
signal \N__45528\ : std_logic;
signal \N__45525\ : std_logic;
signal \N__45522\ : std_logic;
signal \N__45515\ : std_logic;
signal \N__45512\ : std_logic;
signal \N__45509\ : std_logic;
signal \N__45506\ : std_logic;
signal \N__45505\ : std_logic;
signal \N__45504\ : std_logic;
signal \N__45499\ : std_logic;
signal \N__45496\ : std_logic;
signal \N__45493\ : std_logic;
signal \N__45488\ : std_logic;
signal \N__45485\ : std_logic;
signal \N__45482\ : std_logic;
signal \N__45479\ : std_logic;
signal \N__45478\ : std_logic;
signal \N__45475\ : std_logic;
signal \N__45472\ : std_logic;
signal \N__45471\ : std_logic;
signal \N__45466\ : std_logic;
signal \N__45463\ : std_logic;
signal \N__45460\ : std_logic;
signal \N__45455\ : std_logic;
signal \N__45452\ : std_logic;
signal \N__45449\ : std_logic;
signal \N__45446\ : std_logic;
signal \N__45445\ : std_logic;
signal \N__45442\ : std_logic;
signal \N__45439\ : std_logic;
signal \N__45438\ : std_logic;
signal \N__45433\ : std_logic;
signal \N__45430\ : std_logic;
signal \N__45427\ : std_logic;
signal \N__45422\ : std_logic;
signal \N__45419\ : std_logic;
signal \N__45416\ : std_logic;
signal \N__45413\ : std_logic;
signal \N__45410\ : std_logic;
signal \N__45409\ : std_logic;
signal \N__45408\ : std_logic;
signal \N__45403\ : std_logic;
signal \N__45400\ : std_logic;
signal \N__45397\ : std_logic;
signal \N__45392\ : std_logic;
signal \N__45389\ : std_logic;
signal \N__45386\ : std_logic;
signal \N__45383\ : std_logic;
signal \N__45380\ : std_logic;
signal \N__45377\ : std_logic;
signal \N__45376\ : std_logic;
signal \N__45371\ : std_logic;
signal \N__45370\ : std_logic;
signal \N__45367\ : std_logic;
signal \N__45364\ : std_logic;
signal \N__45361\ : std_logic;
signal \N__45356\ : std_logic;
signal \N__45353\ : std_logic;
signal \N__45350\ : std_logic;
signal \N__45347\ : std_logic;
signal \N__45344\ : std_logic;
signal \N__45341\ : std_logic;
signal \N__45340\ : std_logic;
signal \N__45337\ : std_logic;
signal \N__45336\ : std_logic;
signal \N__45333\ : std_logic;
signal \N__45330\ : std_logic;
signal \N__45327\ : std_logic;
signal \N__45324\ : std_logic;
signal \N__45317\ : std_logic;
signal \N__45314\ : std_logic;
signal \N__45311\ : std_logic;
signal \N__45308\ : std_logic;
signal \N__45305\ : std_logic;
signal \N__45302\ : std_logic;
signal \N__45299\ : std_logic;
signal \N__45298\ : std_logic;
signal \N__45297\ : std_logic;
signal \N__45294\ : std_logic;
signal \N__45291\ : std_logic;
signal \N__45288\ : std_logic;
signal \N__45281\ : std_logic;
signal \N__45278\ : std_logic;
signal \N__45277\ : std_logic;
signal \N__45274\ : std_logic;
signal \N__45271\ : std_logic;
signal \N__45266\ : std_logic;
signal \N__45263\ : std_logic;
signal \N__45260\ : std_logic;
signal \N__45259\ : std_logic;
signal \N__45256\ : std_logic;
signal \N__45253\ : std_logic;
signal \N__45252\ : std_logic;
signal \N__45247\ : std_logic;
signal \N__45244\ : std_logic;
signal \N__45241\ : std_logic;
signal \N__45236\ : std_logic;
signal \N__45235\ : std_logic;
signal \N__45232\ : std_logic;
signal \N__45229\ : std_logic;
signal \N__45226\ : std_logic;
signal \N__45223\ : std_logic;
signal \N__45220\ : std_logic;
signal \N__45217\ : std_logic;
signal \N__45212\ : std_logic;
signal \N__45209\ : std_logic;
signal \N__45208\ : std_logic;
signal \N__45205\ : std_logic;
signal \N__45202\ : std_logic;
signal \N__45201\ : std_logic;
signal \N__45196\ : std_logic;
signal \N__45193\ : std_logic;
signal \N__45190\ : std_logic;
signal \N__45185\ : std_logic;
signal \N__45182\ : std_logic;
signal \N__45181\ : std_logic;
signal \N__45176\ : std_logic;
signal \N__45175\ : std_logic;
signal \N__45172\ : std_logic;
signal \N__45169\ : std_logic;
signal \N__45166\ : std_logic;
signal \N__45161\ : std_logic;
signal \N__45160\ : std_logic;
signal \N__45159\ : std_logic;
signal \N__45156\ : std_logic;
signal \N__45155\ : std_logic;
signal \N__45154\ : std_logic;
signal \N__45153\ : std_logic;
signal \N__45150\ : std_logic;
signal \N__45147\ : std_logic;
signal \N__45144\ : std_logic;
signal \N__45139\ : std_logic;
signal \N__45134\ : std_logic;
signal \N__45131\ : std_logic;
signal \N__45128\ : std_logic;
signal \N__45125\ : std_logic;
signal \N__45122\ : std_logic;
signal \N__45117\ : std_logic;
signal \N__45114\ : std_logic;
signal \N__45111\ : std_logic;
signal \N__45104\ : std_logic;
signal \N__45101\ : std_logic;
signal \N__45100\ : std_logic;
signal \N__45095\ : std_logic;
signal \N__45094\ : std_logic;
signal \N__45091\ : std_logic;
signal \N__45088\ : std_logic;
signal \N__45085\ : std_logic;
signal \N__45080\ : std_logic;
signal \N__45077\ : std_logic;
signal \N__45076\ : std_logic;
signal \N__45075\ : std_logic;
signal \N__45072\ : std_logic;
signal \N__45067\ : std_logic;
signal \N__45062\ : std_logic;
signal \N__45059\ : std_logic;
signal \N__45056\ : std_logic;
signal \N__45055\ : std_logic;
signal \N__45052\ : std_logic;
signal \N__45051\ : std_logic;
signal \N__45048\ : std_logic;
signal \N__45045\ : std_logic;
signal \N__45042\ : std_logic;
signal \N__45039\ : std_logic;
signal \N__45036\ : std_logic;
signal \N__45029\ : std_logic;
signal \N__45026\ : std_logic;
signal \N__45025\ : std_logic;
signal \N__45024\ : std_logic;
signal \N__45021\ : std_logic;
signal \N__45018\ : std_logic;
signal \N__45015\ : std_logic;
signal \N__45008\ : std_logic;
signal \N__45005\ : std_logic;
signal \N__45004\ : std_logic;
signal \N__45001\ : std_logic;
signal \N__44998\ : std_logic;
signal \N__44993\ : std_logic;
signal \N__44992\ : std_logic;
signal \N__44989\ : std_logic;
signal \N__44986\ : std_logic;
signal \N__44983\ : std_logic;
signal \N__44978\ : std_logic;
signal \N__44975\ : std_logic;
signal \N__44974\ : std_logic;
signal \N__44973\ : std_logic;
signal \N__44970\ : std_logic;
signal \N__44965\ : std_logic;
signal \N__44960\ : std_logic;
signal \N__44957\ : std_logic;
signal \N__44954\ : std_logic;
signal \N__44953\ : std_logic;
signal \N__44950\ : std_logic;
signal \N__44949\ : std_logic;
signal \N__44946\ : std_logic;
signal \N__44943\ : std_logic;
signal \N__44940\ : std_logic;
signal \N__44937\ : std_logic;
signal \N__44930\ : std_logic;
signal \N__44927\ : std_logic;
signal \N__44926\ : std_logic;
signal \N__44925\ : std_logic;
signal \N__44922\ : std_logic;
signal \N__44919\ : std_logic;
signal \N__44916\ : std_logic;
signal \N__44913\ : std_logic;
signal \N__44910\ : std_logic;
signal \N__44907\ : std_logic;
signal \N__44900\ : std_logic;
signal \N__44897\ : std_logic;
signal \N__44894\ : std_logic;
signal \N__44893\ : std_logic;
signal \N__44890\ : std_logic;
signal \N__44889\ : std_logic;
signal \N__44886\ : std_logic;
signal \N__44883\ : std_logic;
signal \N__44880\ : std_logic;
signal \N__44877\ : std_logic;
signal \N__44870\ : std_logic;
signal \N__44867\ : std_logic;
signal \N__44866\ : std_logic;
signal \N__44865\ : std_logic;
signal \N__44862\ : std_logic;
signal \N__44859\ : std_logic;
signal \N__44856\ : std_logic;
signal \N__44851\ : std_logic;
signal \N__44846\ : std_logic;
signal \N__44843\ : std_logic;
signal \N__44842\ : std_logic;
signal \N__44839\ : std_logic;
signal \N__44836\ : std_logic;
signal \N__44835\ : std_logic;
signal \N__44830\ : std_logic;
signal \N__44827\ : std_logic;
signal \N__44824\ : std_logic;
signal \N__44819\ : std_logic;
signal \N__44816\ : std_logic;
signal \N__44813\ : std_logic;
signal \N__44812\ : std_logic;
signal \N__44811\ : std_logic;
signal \N__44808\ : std_logic;
signal \N__44803\ : std_logic;
signal \N__44800\ : std_logic;
signal \N__44797\ : std_logic;
signal \N__44792\ : std_logic;
signal \N__44789\ : std_logic;
signal \N__44788\ : std_logic;
signal \N__44785\ : std_logic;
signal \N__44782\ : std_logic;
signal \N__44781\ : std_logic;
signal \N__44776\ : std_logic;
signal \N__44773\ : std_logic;
signal \N__44770\ : std_logic;
signal \N__44765\ : std_logic;
signal \N__44762\ : std_logic;
signal \N__44761\ : std_logic;
signal \N__44760\ : std_logic;
signal \N__44757\ : std_logic;
signal \N__44752\ : std_logic;
signal \N__44749\ : std_logic;
signal \N__44746\ : std_logic;
signal \N__44741\ : std_logic;
signal \N__44738\ : std_logic;
signal \N__44737\ : std_logic;
signal \N__44732\ : std_logic;
signal \N__44731\ : std_logic;
signal \N__44728\ : std_logic;
signal \N__44725\ : std_logic;
signal \N__44722\ : std_logic;
signal \N__44717\ : std_logic;
signal \N__44716\ : std_logic;
signal \N__44715\ : std_logic;
signal \N__44712\ : std_logic;
signal \N__44709\ : std_logic;
signal \N__44706\ : std_logic;
signal \N__44701\ : std_logic;
signal \N__44698\ : std_logic;
signal \N__44695\ : std_logic;
signal \N__44692\ : std_logic;
signal \N__44687\ : std_logic;
signal \N__44684\ : std_logic;
signal \N__44683\ : std_logic;
signal \N__44678\ : std_logic;
signal \N__44677\ : std_logic;
signal \N__44674\ : std_logic;
signal \N__44671\ : std_logic;
signal \N__44668\ : std_logic;
signal \N__44663\ : std_logic;
signal \N__44662\ : std_logic;
signal \N__44659\ : std_logic;
signal \N__44656\ : std_logic;
signal \N__44655\ : std_logic;
signal \N__44652\ : std_logic;
signal \N__44649\ : std_logic;
signal \N__44646\ : std_logic;
signal \N__44639\ : std_logic;
signal \N__44636\ : std_logic;
signal \N__44633\ : std_logic;
signal \N__44630\ : std_logic;
signal \N__44629\ : std_logic;
signal \N__44626\ : std_logic;
signal \N__44625\ : std_logic;
signal \N__44622\ : std_logic;
signal \N__44619\ : std_logic;
signal \N__44616\ : std_logic;
signal \N__44613\ : std_logic;
signal \N__44610\ : std_logic;
signal \N__44603\ : std_logic;
signal \N__44602\ : std_logic;
signal \N__44601\ : std_logic;
signal \N__44598\ : std_logic;
signal \N__44595\ : std_logic;
signal \N__44594\ : std_logic;
signal \N__44591\ : std_logic;
signal \N__44586\ : std_logic;
signal \N__44581\ : std_logic;
signal \N__44576\ : std_logic;
signal \N__44573\ : std_logic;
signal \N__44570\ : std_logic;
signal \N__44569\ : std_logic;
signal \N__44566\ : std_logic;
signal \N__44563\ : std_logic;
signal \N__44558\ : std_logic;
signal \N__44557\ : std_logic;
signal \N__44554\ : std_logic;
signal \N__44551\ : std_logic;
signal \N__44548\ : std_logic;
signal \N__44543\ : std_logic;
signal \N__44542\ : std_logic;
signal \N__44539\ : std_logic;
signal \N__44536\ : std_logic;
signal \N__44533\ : std_logic;
signal \N__44530\ : std_logic;
signal \N__44527\ : std_logic;
signal \N__44524\ : std_logic;
signal \N__44519\ : std_logic;
signal \N__44516\ : std_logic;
signal \N__44515\ : std_logic;
signal \N__44512\ : std_logic;
signal \N__44511\ : std_logic;
signal \N__44508\ : std_logic;
signal \N__44505\ : std_logic;
signal \N__44502\ : std_logic;
signal \N__44499\ : std_logic;
signal \N__44492\ : std_logic;
signal \N__44489\ : std_logic;
signal \N__44488\ : std_logic;
signal \N__44485\ : std_logic;
signal \N__44482\ : std_logic;
signal \N__44477\ : std_logic;
signal \N__44474\ : std_logic;
signal \N__44471\ : std_logic;
signal \N__44468\ : std_logic;
signal \N__44465\ : std_logic;
signal \N__44462\ : std_logic;
signal \N__44459\ : std_logic;
signal \N__44456\ : std_logic;
signal \N__44453\ : std_logic;
signal \N__44450\ : std_logic;
signal \N__44449\ : std_logic;
signal \N__44446\ : std_logic;
signal \N__44445\ : std_logic;
signal \N__44444\ : std_logic;
signal \N__44441\ : std_logic;
signal \N__44438\ : std_logic;
signal \N__44435\ : std_logic;
signal \N__44432\ : std_logic;
signal \N__44429\ : std_logic;
signal \N__44424\ : std_logic;
signal \N__44421\ : std_logic;
signal \N__44418\ : std_logic;
signal \N__44417\ : std_logic;
signal \N__44414\ : std_logic;
signal \N__44411\ : std_logic;
signal \N__44408\ : std_logic;
signal \N__44405\ : std_logic;
signal \N__44402\ : std_logic;
signal \N__44399\ : std_logic;
signal \N__44394\ : std_logic;
signal \N__44387\ : std_logic;
signal \N__44386\ : std_logic;
signal \N__44385\ : std_logic;
signal \N__44384\ : std_logic;
signal \N__44379\ : std_logic;
signal \N__44376\ : std_logic;
signal \N__44373\ : std_logic;
signal \N__44370\ : std_logic;
signal \N__44365\ : std_logic;
signal \N__44362\ : std_logic;
signal \N__44357\ : std_logic;
signal \N__44354\ : std_logic;
signal \N__44351\ : std_logic;
signal \N__44348\ : std_logic;
signal \N__44345\ : std_logic;
signal \N__44342\ : std_logic;
signal \N__44341\ : std_logic;
signal \N__44338\ : std_logic;
signal \N__44335\ : std_logic;
signal \N__44330\ : std_logic;
signal \N__44329\ : std_logic;
signal \N__44326\ : std_logic;
signal \N__44323\ : std_logic;
signal \N__44318\ : std_logic;
signal \N__44317\ : std_logic;
signal \N__44314\ : std_logic;
signal \N__44311\ : std_logic;
signal \N__44308\ : std_logic;
signal \N__44303\ : std_logic;
signal \N__44302\ : std_logic;
signal \N__44299\ : std_logic;
signal \N__44296\ : std_logic;
signal \N__44291\ : std_logic;
signal \N__44288\ : std_logic;
signal \N__44285\ : std_logic;
signal \N__44282\ : std_logic;
signal \N__44281\ : std_logic;
signal \N__44278\ : std_logic;
signal \N__44275\ : std_logic;
signal \N__44274\ : std_logic;
signal \N__44273\ : std_logic;
signal \N__44270\ : std_logic;
signal \N__44267\ : std_logic;
signal \N__44264\ : std_logic;
signal \N__44261\ : std_logic;
signal \N__44260\ : std_logic;
signal \N__44257\ : std_logic;
signal \N__44254\ : std_logic;
signal \N__44251\ : std_logic;
signal \N__44248\ : std_logic;
signal \N__44245\ : std_logic;
signal \N__44236\ : std_logic;
signal \N__44233\ : std_logic;
signal \N__44230\ : std_logic;
signal \N__44225\ : std_logic;
signal \N__44222\ : std_logic;
signal \N__44219\ : std_logic;
signal \N__44216\ : std_logic;
signal \N__44213\ : std_logic;
signal \N__44210\ : std_logic;
signal \N__44207\ : std_logic;
signal \N__44206\ : std_logic;
signal \N__44205\ : std_logic;
signal \N__44204\ : std_logic;
signal \N__44201\ : std_logic;
signal \N__44200\ : std_logic;
signal \N__44199\ : std_logic;
signal \N__44198\ : std_logic;
signal \N__44189\ : std_logic;
signal \N__44188\ : std_logic;
signal \N__44187\ : std_logic;
signal \N__44186\ : std_logic;
signal \N__44185\ : std_logic;
signal \N__44184\ : std_logic;
signal \N__44183\ : std_logic;
signal \N__44182\ : std_logic;
signal \N__44181\ : std_logic;
signal \N__44180\ : std_logic;
signal \N__44179\ : std_logic;
signal \N__44178\ : std_logic;
signal \N__44177\ : std_logic;
signal \N__44174\ : std_logic;
signal \N__44173\ : std_logic;
signal \N__44170\ : std_logic;
signal \N__44169\ : std_logic;
signal \N__44168\ : std_logic;
signal \N__44167\ : std_logic;
signal \N__44166\ : std_logic;
signal \N__44165\ : std_logic;
signal \N__44164\ : std_logic;
signal \N__44161\ : std_logic;
signal \N__44158\ : std_logic;
signal \N__44157\ : std_logic;
signal \N__44156\ : std_logic;
signal \N__44155\ : std_logic;
signal \N__44154\ : std_logic;
signal \N__44151\ : std_logic;
signal \N__44148\ : std_logic;
signal \N__44145\ : std_logic;
signal \N__44144\ : std_logic;
signal \N__44141\ : std_logic;
signal \N__44140\ : std_logic;
signal \N__44139\ : std_logic;
signal \N__44126\ : std_logic;
signal \N__44109\ : std_logic;
signal \N__44100\ : std_logic;
signal \N__44097\ : std_logic;
signal \N__44094\ : std_logic;
signal \N__44091\ : std_logic;
signal \N__44088\ : std_logic;
signal \N__44087\ : std_logic;
signal \N__44086\ : std_logic;
signal \N__44085\ : std_logic;
signal \N__44084\ : std_logic;
signal \N__44081\ : std_logic;
signal \N__44066\ : std_logic;
signal \N__44063\ : std_logic;
signal \N__44062\ : std_logic;
signal \N__44061\ : std_logic;
signal \N__44060\ : std_logic;
signal \N__44055\ : std_logic;
signal \N__44052\ : std_logic;
signal \N__44049\ : std_logic;
signal \N__44046\ : std_logic;
signal \N__44039\ : std_logic;
signal \N__44034\ : std_logic;
signal \N__44031\ : std_logic;
signal \N__44028\ : std_logic;
signal \N__44025\ : std_logic;
signal \N__44018\ : std_logic;
signal \N__44017\ : std_logic;
signal \N__44014\ : std_logic;
signal \N__44009\ : std_logic;
signal \N__44006\ : std_logic;
signal \N__44001\ : std_logic;
signal \N__43998\ : std_logic;
signal \N__43995\ : std_logic;
signal \N__43990\ : std_logic;
signal \N__43987\ : std_logic;
signal \N__43984\ : std_logic;
signal \N__43979\ : std_logic;
signal \N__43976\ : std_logic;
signal \N__43969\ : std_logic;
signal \N__43958\ : std_logic;
signal \N__43957\ : std_logic;
signal \N__43956\ : std_logic;
signal \N__43955\ : std_logic;
signal \N__43954\ : std_logic;
signal \N__43951\ : std_logic;
signal \N__43948\ : std_logic;
signal \N__43945\ : std_logic;
signal \N__43942\ : std_logic;
signal \N__43939\ : std_logic;
signal \N__43936\ : std_logic;
signal \N__43933\ : std_logic;
signal \N__43930\ : std_logic;
signal \N__43927\ : std_logic;
signal \N__43924\ : std_logic;
signal \N__43913\ : std_logic;
signal \N__43912\ : std_logic;
signal \N__43911\ : std_logic;
signal \N__43910\ : std_logic;
signal \N__43901\ : std_logic;
signal \N__43900\ : std_logic;
signal \N__43899\ : std_logic;
signal \N__43898\ : std_logic;
signal \N__43897\ : std_logic;
signal \N__43896\ : std_logic;
signal \N__43895\ : std_logic;
signal \N__43894\ : std_logic;
signal \N__43893\ : std_logic;
signal \N__43892\ : std_logic;
signal \N__43889\ : std_logic;
signal \N__43888\ : std_logic;
signal \N__43887\ : std_logic;
signal \N__43880\ : std_logic;
signal \N__43879\ : std_logic;
signal \N__43878\ : std_logic;
signal \N__43875\ : std_logic;
signal \N__43864\ : std_logic;
signal \N__43863\ : std_logic;
signal \N__43862\ : std_logic;
signal \N__43861\ : std_logic;
signal \N__43860\ : std_logic;
signal \N__43859\ : std_logic;
signal \N__43858\ : std_logic;
signal \N__43857\ : std_logic;
signal \N__43856\ : std_logic;
signal \N__43855\ : std_logic;
signal \N__43854\ : std_logic;
signal \N__43853\ : std_logic;
signal \N__43852\ : std_logic;
signal \N__43851\ : std_logic;
signal \N__43850\ : std_logic;
signal \N__43849\ : std_logic;
signal \N__43848\ : std_logic;
signal \N__43847\ : std_logic;
signal \N__43846\ : std_logic;
signal \N__43845\ : std_logic;
signal \N__43844\ : std_logic;
signal \N__43841\ : std_logic;
signal \N__43836\ : std_logic;
signal \N__43833\ : std_logic;
signal \N__43828\ : std_logic;
signal \N__43827\ : std_logic;
signal \N__43824\ : std_logic;
signal \N__43821\ : std_logic;
signal \N__43804\ : std_logic;
signal \N__43795\ : std_logic;
signal \N__43792\ : std_logic;
signal \N__43777\ : std_logic;
signal \N__43772\ : std_logic;
signal \N__43767\ : std_logic;
signal \N__43764\ : std_logic;
signal \N__43761\ : std_logic;
signal \N__43754\ : std_logic;
signal \N__43749\ : std_logic;
signal \N__43746\ : std_logic;
signal \N__43741\ : std_logic;
signal \N__43730\ : std_logic;
signal \N__43727\ : std_logic;
signal \N__43724\ : std_logic;
signal \N__43721\ : std_logic;
signal \N__43718\ : std_logic;
signal \N__43715\ : std_logic;
signal \N__43712\ : std_logic;
signal \N__43711\ : std_logic;
signal \N__43708\ : std_logic;
signal \N__43707\ : std_logic;
signal \N__43704\ : std_logic;
signal \N__43701\ : std_logic;
signal \N__43700\ : std_logic;
signal \N__43697\ : std_logic;
signal \N__43694\ : std_logic;
signal \N__43691\ : std_logic;
signal \N__43688\ : std_logic;
signal \N__43687\ : std_logic;
signal \N__43684\ : std_logic;
signal \N__43681\ : std_logic;
signal \N__43676\ : std_logic;
signal \N__43673\ : std_logic;
signal \N__43670\ : std_logic;
signal \N__43667\ : std_logic;
signal \N__43662\ : std_logic;
signal \N__43659\ : std_logic;
signal \N__43654\ : std_logic;
signal \N__43649\ : std_logic;
signal \N__43648\ : std_logic;
signal \N__43647\ : std_logic;
signal \N__43646\ : std_logic;
signal \N__43645\ : std_logic;
signal \N__43642\ : std_logic;
signal \N__43639\ : std_logic;
signal \N__43638\ : std_logic;
signal \N__43635\ : std_logic;
signal \N__43632\ : std_logic;
signal \N__43623\ : std_logic;
signal \N__43620\ : std_logic;
signal \N__43619\ : std_logic;
signal \N__43612\ : std_logic;
signal \N__43609\ : std_logic;
signal \N__43604\ : std_logic;
signal \N__43603\ : std_logic;
signal \N__43602\ : std_logic;
signal \N__43601\ : std_logic;
signal \N__43598\ : std_logic;
signal \N__43595\ : std_logic;
signal \N__43594\ : std_logic;
signal \N__43593\ : std_logic;
signal \N__43592\ : std_logic;
signal \N__43591\ : std_logic;
signal \N__43588\ : std_logic;
signal \N__43585\ : std_logic;
signal \N__43582\ : std_logic;
signal \N__43577\ : std_logic;
signal \N__43566\ : std_logic;
signal \N__43563\ : std_logic;
signal \N__43560\ : std_logic;
signal \N__43553\ : std_logic;
signal \N__43550\ : std_logic;
signal \N__43547\ : std_logic;
signal \N__43546\ : std_logic;
signal \N__43545\ : std_logic;
signal \N__43544\ : std_logic;
signal \N__43543\ : std_logic;
signal \N__43542\ : std_logic;
signal \N__43541\ : std_logic;
signal \N__43538\ : std_logic;
signal \N__43527\ : std_logic;
signal \N__43524\ : std_logic;
signal \N__43523\ : std_logic;
signal \N__43520\ : std_logic;
signal \N__43517\ : std_logic;
signal \N__43514\ : std_logic;
signal \N__43511\ : std_logic;
signal \N__43502\ : std_logic;
signal \N__43501\ : std_logic;
signal \N__43498\ : std_logic;
signal \N__43497\ : std_logic;
signal \N__43494\ : std_logic;
signal \N__43491\ : std_logic;
signal \N__43488\ : std_logic;
signal \N__43485\ : std_logic;
signal \N__43480\ : std_logic;
signal \N__43477\ : std_logic;
signal \N__43474\ : std_logic;
signal \N__43471\ : std_logic;
signal \N__43468\ : std_logic;
signal \N__43463\ : std_logic;
signal \N__43462\ : std_logic;
signal \N__43461\ : std_logic;
signal \N__43458\ : std_logic;
signal \N__43455\ : std_logic;
signal \N__43452\ : std_logic;
signal \N__43451\ : std_logic;
signal \N__43448\ : std_logic;
signal \N__43445\ : std_logic;
signal \N__43442\ : std_logic;
signal \N__43439\ : std_logic;
signal \N__43434\ : std_logic;
signal \N__43429\ : std_logic;
signal \N__43424\ : std_logic;
signal \N__43423\ : std_logic;
signal \N__43420\ : std_logic;
signal \N__43419\ : std_logic;
signal \N__43416\ : std_logic;
signal \N__43413\ : std_logic;
signal \N__43410\ : std_logic;
signal \N__43403\ : std_logic;
signal \N__43402\ : std_logic;
signal \N__43401\ : std_logic;
signal \N__43398\ : std_logic;
signal \N__43395\ : std_logic;
signal \N__43392\ : std_logic;
signal \N__43389\ : std_logic;
signal \N__43386\ : std_logic;
signal \N__43383\ : std_logic;
signal \N__43380\ : std_logic;
signal \N__43377\ : std_logic;
signal \N__43370\ : std_logic;
signal \N__43367\ : std_logic;
signal \N__43366\ : std_logic;
signal \N__43363\ : std_logic;
signal \N__43362\ : std_logic;
signal \N__43359\ : std_logic;
signal \N__43356\ : std_logic;
signal \N__43353\ : std_logic;
signal \N__43346\ : std_logic;
signal \N__43345\ : std_logic;
signal \N__43344\ : std_logic;
signal \N__43343\ : std_logic;
signal \N__43338\ : std_logic;
signal \N__43335\ : std_logic;
signal \N__43334\ : std_logic;
signal \N__43333\ : std_logic;
signal \N__43330\ : std_logic;
signal \N__43327\ : std_logic;
signal \N__43320\ : std_logic;
signal \N__43317\ : std_logic;
signal \N__43314\ : std_logic;
signal \N__43311\ : std_logic;
signal \N__43304\ : std_logic;
signal \N__43301\ : std_logic;
signal \N__43298\ : std_logic;
signal \N__43297\ : std_logic;
signal \N__43296\ : std_logic;
signal \N__43293\ : std_logic;
signal \N__43290\ : std_logic;
signal \N__43289\ : std_logic;
signal \N__43286\ : std_logic;
signal \N__43283\ : std_logic;
signal \N__43280\ : std_logic;
signal \N__43275\ : std_logic;
signal \N__43272\ : std_logic;
signal \N__43267\ : std_logic;
signal \N__43264\ : std_logic;
signal \N__43261\ : std_logic;
signal \N__43256\ : std_logic;
signal \N__43255\ : std_logic;
signal \N__43254\ : std_logic;
signal \N__43253\ : std_logic;
signal \N__43246\ : std_logic;
signal \N__43243\ : std_logic;
signal \N__43242\ : std_logic;
signal \N__43241\ : std_logic;
signal \N__43240\ : std_logic;
signal \N__43239\ : std_logic;
signal \N__43236\ : std_logic;
signal \N__43233\ : std_logic;
signal \N__43230\ : std_logic;
signal \N__43225\ : std_logic;
signal \N__43222\ : std_logic;
signal \N__43211\ : std_logic;
signal \N__43210\ : std_logic;
signal \N__43207\ : std_logic;
signal \N__43206\ : std_logic;
signal \N__43205\ : std_logic;
signal \N__43202\ : std_logic;
signal \N__43199\ : std_logic;
signal \N__43194\ : std_logic;
signal \N__43191\ : std_logic;
signal \N__43186\ : std_logic;
signal \N__43183\ : std_logic;
signal \N__43180\ : std_logic;
signal \N__43175\ : std_logic;
signal \N__43172\ : std_logic;
signal \N__43169\ : std_logic;
signal \N__43166\ : std_logic;
signal \N__43163\ : std_logic;
signal \N__43160\ : std_logic;
signal \N__43157\ : std_logic;
signal \N__43154\ : std_logic;
signal \N__43153\ : std_logic;
signal \N__43152\ : std_logic;
signal \N__43151\ : std_logic;
signal \N__43150\ : std_logic;
signal \N__43147\ : std_logic;
signal \N__43144\ : std_logic;
signal \N__43141\ : std_logic;
signal \N__43136\ : std_logic;
signal \N__43127\ : std_logic;
signal \N__43124\ : std_logic;
signal \N__43121\ : std_logic;
signal \N__43118\ : std_logic;
signal \N__43117\ : std_logic;
signal \N__43114\ : std_logic;
signal \N__43111\ : std_logic;
signal \N__43106\ : std_logic;
signal \N__43103\ : std_logic;
signal \N__43100\ : std_logic;
signal \N__43097\ : std_logic;
signal \N__43096\ : std_logic;
signal \N__43093\ : std_logic;
signal \N__43090\ : std_logic;
signal \N__43087\ : std_logic;
signal \N__43084\ : std_logic;
signal \N__43081\ : std_logic;
signal \N__43078\ : std_logic;
signal \N__43077\ : std_logic;
signal \N__43076\ : std_logic;
signal \N__43071\ : std_logic;
signal \N__43068\ : std_logic;
signal \N__43065\ : std_logic;
signal \N__43060\ : std_logic;
signal \N__43055\ : std_logic;
signal \N__43054\ : std_logic;
signal \N__43051\ : std_logic;
signal \N__43050\ : std_logic;
signal \N__43043\ : std_logic;
signal \N__43040\ : std_logic;
signal \N__43037\ : std_logic;
signal \N__43034\ : std_logic;
signal \N__43033\ : std_logic;
signal \N__43030\ : std_logic;
signal \N__43027\ : std_logic;
signal \N__43024\ : std_logic;
signal \N__43023\ : std_logic;
signal \N__43020\ : std_logic;
signal \N__43017\ : std_logic;
signal \N__43014\ : std_logic;
signal \N__43011\ : std_logic;
signal \N__43004\ : std_logic;
signal \N__43003\ : std_logic;
signal \N__42998\ : std_logic;
signal \N__42995\ : std_logic;
signal \N__42992\ : std_logic;
signal \N__42989\ : std_logic;
signal \N__42986\ : std_logic;
signal \N__42983\ : std_logic;
signal \N__42982\ : std_logic;
signal \N__42981\ : std_logic;
signal \N__42980\ : std_logic;
signal \N__42971\ : std_logic;
signal \N__42970\ : std_logic;
signal \N__42969\ : std_logic;
signal \N__42968\ : std_logic;
signal \N__42967\ : std_logic;
signal \N__42966\ : std_logic;
signal \N__42965\ : std_logic;
signal \N__42964\ : std_logic;
signal \N__42963\ : std_logic;
signal \N__42962\ : std_logic;
signal \N__42961\ : std_logic;
signal \N__42960\ : std_logic;
signal \N__42959\ : std_logic;
signal \N__42958\ : std_logic;
signal \N__42957\ : std_logic;
signal \N__42956\ : std_logic;
signal \N__42955\ : std_logic;
signal \N__42954\ : std_logic;
signal \N__42953\ : std_logic;
signal \N__42952\ : std_logic;
signal \N__42951\ : std_logic;
signal \N__42950\ : std_logic;
signal \N__42949\ : std_logic;
signal \N__42948\ : std_logic;
signal \N__42947\ : std_logic;
signal \N__42946\ : std_logic;
signal \N__42945\ : std_logic;
signal \N__42942\ : std_logic;
signal \N__42937\ : std_logic;
signal \N__42928\ : std_logic;
signal \N__42919\ : std_logic;
signal \N__42910\ : std_logic;
signal \N__42901\ : std_logic;
signal \N__42892\ : std_logic;
signal \N__42883\ : std_logic;
signal \N__42878\ : std_logic;
signal \N__42873\ : std_logic;
signal \N__42860\ : std_logic;
signal \N__42857\ : std_logic;
signal \N__42856\ : std_logic;
signal \N__42853\ : std_logic;
signal \N__42850\ : std_logic;
signal \N__42849\ : std_logic;
signal \N__42846\ : std_logic;
signal \N__42843\ : std_logic;
signal \N__42840\ : std_logic;
signal \N__42839\ : std_logic;
signal \N__42832\ : std_logic;
signal \N__42829\ : std_logic;
signal \N__42826\ : std_logic;
signal \N__42823\ : std_logic;
signal \N__42818\ : std_logic;
signal \N__42815\ : std_logic;
signal \N__42812\ : std_logic;
signal \N__42809\ : std_logic;
signal \N__42806\ : std_logic;
signal \N__42803\ : std_logic;
signal \N__42800\ : std_logic;
signal \N__42797\ : std_logic;
signal \N__42796\ : std_logic;
signal \N__42793\ : std_logic;
signal \N__42790\ : std_logic;
signal \N__42789\ : std_logic;
signal \N__42786\ : std_logic;
signal \N__42783\ : std_logic;
signal \N__42780\ : std_logic;
signal \N__42775\ : std_logic;
signal \N__42770\ : std_logic;
signal \N__42769\ : std_logic;
signal \N__42768\ : std_logic;
signal \N__42765\ : std_logic;
signal \N__42764\ : std_logic;
signal \N__42761\ : std_logic;
signal \N__42758\ : std_logic;
signal \N__42755\ : std_logic;
signal \N__42752\ : std_logic;
signal \N__42749\ : std_logic;
signal \N__42744\ : std_logic;
signal \N__42737\ : std_logic;
signal \N__42734\ : std_logic;
signal \N__42731\ : std_logic;
signal \N__42728\ : std_logic;
signal \N__42725\ : std_logic;
signal \N__42722\ : std_logic;
signal \N__42719\ : std_logic;
signal \N__42716\ : std_logic;
signal \N__42713\ : std_logic;
signal \N__42710\ : std_logic;
signal \N__42707\ : std_logic;
signal \N__42704\ : std_logic;
signal \N__42701\ : std_logic;
signal \N__42698\ : std_logic;
signal \N__42695\ : std_logic;
signal \N__42692\ : std_logic;
signal \N__42689\ : std_logic;
signal \N__42686\ : std_logic;
signal \N__42683\ : std_logic;
signal \N__42682\ : std_logic;
signal \N__42679\ : std_logic;
signal \N__42676\ : std_logic;
signal \N__42671\ : std_logic;
signal \N__42668\ : std_logic;
signal \N__42667\ : std_logic;
signal \N__42664\ : std_logic;
signal \N__42661\ : std_logic;
signal \N__42658\ : std_logic;
signal \N__42653\ : std_logic;
signal \N__42652\ : std_logic;
signal \N__42651\ : std_logic;
signal \N__42650\ : std_logic;
signal \N__42649\ : std_logic;
signal \N__42648\ : std_logic;
signal \N__42647\ : std_logic;
signal \N__42646\ : std_logic;
signal \N__42645\ : std_logic;
signal \N__42644\ : std_logic;
signal \N__42641\ : std_logic;
signal \N__42640\ : std_logic;
signal \N__42637\ : std_logic;
signal \N__42636\ : std_logic;
signal \N__42633\ : std_logic;
signal \N__42632\ : std_logic;
signal \N__42631\ : std_logic;
signal \N__42630\ : std_logic;
signal \N__42629\ : std_logic;
signal \N__42628\ : std_logic;
signal \N__42627\ : std_logic;
signal \N__42626\ : std_logic;
signal \N__42625\ : std_logic;
signal \N__42624\ : std_logic;
signal \N__42623\ : std_logic;
signal \N__42622\ : std_logic;
signal \N__42621\ : std_logic;
signal \N__42620\ : std_logic;
signal \N__42615\ : std_logic;
signal \N__42612\ : std_logic;
signal \N__42605\ : std_logic;
signal \N__42594\ : std_logic;
signal \N__42583\ : std_logic;
signal \N__42574\ : std_logic;
signal \N__42571\ : std_logic;
signal \N__42564\ : std_logic;
signal \N__42561\ : std_logic;
signal \N__42560\ : std_logic;
signal \N__42559\ : std_logic;
signal \N__42558\ : std_logic;
signal \N__42555\ : std_logic;
signal \N__42552\ : std_logic;
signal \N__42551\ : std_logic;
signal \N__42544\ : std_logic;
signal \N__42535\ : std_logic;
signal \N__42528\ : std_logic;
signal \N__42527\ : std_logic;
signal \N__42526\ : std_logic;
signal \N__42525\ : std_logic;
signal \N__42522\ : std_logic;
signal \N__42519\ : std_logic;
signal \N__42516\ : std_logic;
signal \N__42509\ : std_logic;
signal \N__42502\ : std_logic;
signal \N__42491\ : std_logic;
signal \N__42488\ : std_logic;
signal \N__42485\ : std_logic;
signal \N__42482\ : std_logic;
signal \N__42481\ : std_logic;
signal \N__42480\ : std_logic;
signal \N__42477\ : std_logic;
signal \N__42472\ : std_logic;
signal \N__42467\ : std_logic;
signal \N__42466\ : std_logic;
signal \N__42465\ : std_logic;
signal \N__42464\ : std_logic;
signal \N__42463\ : std_logic;
signal \N__42462\ : std_logic;
signal \N__42461\ : std_logic;
signal \N__42454\ : std_logic;
signal \N__42447\ : std_logic;
signal \N__42446\ : std_logic;
signal \N__42445\ : std_logic;
signal \N__42444\ : std_logic;
signal \N__42443\ : std_logic;
signal \N__42442\ : std_logic;
signal \N__42441\ : std_logic;
signal \N__42440\ : std_logic;
signal \N__42439\ : std_logic;
signal \N__42438\ : std_logic;
signal \N__42435\ : std_logic;
signal \N__42432\ : std_logic;
signal \N__42429\ : std_logic;
signal \N__42422\ : std_logic;
signal \N__42421\ : std_logic;
signal \N__42420\ : std_logic;
signal \N__42419\ : std_logic;
signal \N__42418\ : std_logic;
signal \N__42417\ : std_logic;
signal \N__42412\ : std_logic;
signal \N__42403\ : std_logic;
signal \N__42400\ : std_logic;
signal \N__42393\ : std_logic;
signal \N__42384\ : std_logic;
signal \N__42381\ : std_logic;
signal \N__42380\ : std_logic;
signal \N__42379\ : std_logic;
signal \N__42378\ : std_logic;
signal \N__42375\ : std_logic;
signal \N__42372\ : std_logic;
signal \N__42363\ : std_logic;
signal \N__42356\ : std_logic;
signal \N__42347\ : std_logic;
signal \N__42346\ : std_logic;
signal \N__42343\ : std_logic;
signal \N__42340\ : std_logic;
signal \N__42339\ : std_logic;
signal \N__42336\ : std_logic;
signal \N__42333\ : std_logic;
signal \N__42330\ : std_logic;
signal \N__42329\ : std_logic;
signal \N__42326\ : std_logic;
signal \N__42323\ : std_logic;
signal \N__42320\ : std_logic;
signal \N__42319\ : std_logic;
signal \N__42316\ : std_logic;
signal \N__42311\ : std_logic;
signal \N__42308\ : std_logic;
signal \N__42305\ : std_logic;
signal \N__42296\ : std_logic;
signal \N__42293\ : std_logic;
signal \N__42290\ : std_logic;
signal \N__42287\ : std_logic;
signal \N__42284\ : std_logic;
signal \N__42281\ : std_logic;
signal \N__42278\ : std_logic;
signal \N__42275\ : std_logic;
signal \N__42274\ : std_logic;
signal \N__42271\ : std_logic;
signal \N__42268\ : std_logic;
signal \N__42265\ : std_logic;
signal \N__42260\ : std_logic;
signal \N__42259\ : std_logic;
signal \N__42256\ : std_logic;
signal \N__42253\ : std_logic;
signal \N__42250\ : std_logic;
signal \N__42247\ : std_logic;
signal \N__42244\ : std_logic;
signal \N__42243\ : std_logic;
signal \N__42240\ : std_logic;
signal \N__42237\ : std_logic;
signal \N__42234\ : std_logic;
signal \N__42233\ : std_logic;
signal \N__42230\ : std_logic;
signal \N__42225\ : std_logic;
signal \N__42222\ : std_logic;
signal \N__42219\ : std_logic;
signal \N__42216\ : std_logic;
signal \N__42209\ : std_logic;
signal \N__42206\ : std_logic;
signal \N__42205\ : std_logic;
signal \N__42204\ : std_logic;
signal \N__42201\ : std_logic;
signal \N__42196\ : std_logic;
signal \N__42191\ : std_logic;
signal \N__42190\ : std_logic;
signal \N__42187\ : std_logic;
signal \N__42184\ : std_logic;
signal \N__42183\ : std_logic;
signal \N__42182\ : std_logic;
signal \N__42181\ : std_logic;
signal \N__42178\ : std_logic;
signal \N__42175\ : std_logic;
signal \N__42172\ : std_logic;
signal \N__42169\ : std_logic;
signal \N__42166\ : std_logic;
signal \N__42163\ : std_logic;
signal \N__42160\ : std_logic;
signal \N__42157\ : std_logic;
signal \N__42154\ : std_logic;
signal \N__42151\ : std_logic;
signal \N__42148\ : std_logic;
signal \N__42141\ : std_logic;
signal \N__42134\ : std_logic;
signal \N__42131\ : std_logic;
signal \N__42130\ : std_logic;
signal \N__42129\ : std_logic;
signal \N__42126\ : std_logic;
signal \N__42123\ : std_logic;
signal \N__42120\ : std_logic;
signal \N__42117\ : std_logic;
signal \N__42114\ : std_logic;
signal \N__42111\ : std_logic;
signal \N__42104\ : std_logic;
signal \N__42103\ : std_logic;
signal \N__42102\ : std_logic;
signal \N__42101\ : std_logic;
signal \N__42100\ : std_logic;
signal \N__42099\ : std_logic;
signal \N__42094\ : std_logic;
signal \N__42093\ : std_logic;
signal \N__42092\ : std_logic;
signal \N__42089\ : std_logic;
signal \N__42082\ : std_logic;
signal \N__42079\ : std_logic;
signal \N__42076\ : std_logic;
signal \N__42073\ : std_logic;
signal \N__42070\ : std_logic;
signal \N__42067\ : std_logic;
signal \N__42062\ : std_logic;
signal \N__42053\ : std_logic;
signal \N__42050\ : std_logic;
signal \N__42049\ : std_logic;
signal \N__42048\ : std_logic;
signal \N__42045\ : std_logic;
signal \N__42042\ : std_logic;
signal \N__42039\ : std_logic;
signal \N__42036\ : std_logic;
signal \N__42033\ : std_logic;
signal \N__42028\ : std_logic;
signal \N__42025\ : std_logic;
signal \N__42020\ : std_logic;
signal \N__42019\ : std_logic;
signal \N__42014\ : std_logic;
signal \N__42013\ : std_logic;
signal \N__42010\ : std_logic;
signal \N__42007\ : std_logic;
signal \N__42004\ : std_logic;
signal \N__41999\ : std_logic;
signal \N__41998\ : std_logic;
signal \N__41995\ : std_logic;
signal \N__41992\ : std_logic;
signal \N__41991\ : std_logic;
signal \N__41988\ : std_logic;
signal \N__41985\ : std_logic;
signal \N__41982\ : std_logic;
signal \N__41979\ : std_logic;
signal \N__41976\ : std_logic;
signal \N__41973\ : std_logic;
signal \N__41966\ : std_logic;
signal \N__41963\ : std_logic;
signal \N__41960\ : std_logic;
signal \N__41957\ : std_logic;
signal \N__41954\ : std_logic;
signal \N__41951\ : std_logic;
signal \N__41948\ : std_logic;
signal \N__41945\ : std_logic;
signal \N__41942\ : std_logic;
signal \N__41939\ : std_logic;
signal \N__41936\ : std_logic;
signal \N__41933\ : std_logic;
signal \N__41932\ : std_logic;
signal \N__41931\ : std_logic;
signal \N__41930\ : std_logic;
signal \N__41927\ : std_logic;
signal \N__41922\ : std_logic;
signal \N__41919\ : std_logic;
signal \N__41916\ : std_logic;
signal \N__41913\ : std_logic;
signal \N__41910\ : std_logic;
signal \N__41907\ : std_logic;
signal \N__41904\ : std_logic;
signal \N__41901\ : std_logic;
signal \N__41894\ : std_logic;
signal \N__41891\ : std_logic;
signal \N__41888\ : std_logic;
signal \N__41887\ : std_logic;
signal \N__41886\ : std_logic;
signal \N__41883\ : std_logic;
signal \N__41880\ : std_logic;
signal \N__41877\ : std_logic;
signal \N__41876\ : std_logic;
signal \N__41873\ : std_logic;
signal \N__41870\ : std_logic;
signal \N__41867\ : std_logic;
signal \N__41864\ : std_logic;
signal \N__41861\ : std_logic;
signal \N__41856\ : std_logic;
signal \N__41853\ : std_logic;
signal \N__41850\ : std_logic;
signal \N__41847\ : std_logic;
signal \N__41844\ : std_logic;
signal \N__41837\ : std_logic;
signal \N__41836\ : std_logic;
signal \N__41833\ : std_logic;
signal \N__41830\ : std_logic;
signal \N__41825\ : std_logic;
signal \N__41824\ : std_logic;
signal \N__41821\ : std_logic;
signal \N__41818\ : std_logic;
signal \N__41813\ : std_logic;
signal \N__41810\ : std_logic;
signal \N__41809\ : std_logic;
signal \N__41804\ : std_logic;
signal \N__41801\ : std_logic;
signal \N__41798\ : std_logic;
signal \N__41797\ : std_logic;
signal \N__41794\ : std_logic;
signal \N__41793\ : std_logic;
signal \N__41792\ : std_logic;
signal \N__41789\ : std_logic;
signal \N__41786\ : std_logic;
signal \N__41783\ : std_logic;
signal \N__41780\ : std_logic;
signal \N__41777\ : std_logic;
signal \N__41768\ : std_logic;
signal \N__41767\ : std_logic;
signal \N__41764\ : std_logic;
signal \N__41763\ : std_logic;
signal \N__41760\ : std_logic;
signal \N__41757\ : std_logic;
signal \N__41756\ : std_logic;
signal \N__41753\ : std_logic;
signal \N__41750\ : std_logic;
signal \N__41747\ : std_logic;
signal \N__41744\ : std_logic;
signal \N__41741\ : std_logic;
signal \N__41740\ : std_logic;
signal \N__41737\ : std_logic;
signal \N__41734\ : std_logic;
signal \N__41731\ : std_logic;
signal \N__41728\ : std_logic;
signal \N__41725\ : std_logic;
signal \N__41722\ : std_logic;
signal \N__41715\ : std_logic;
signal \N__41708\ : std_logic;
signal \N__41705\ : std_logic;
signal \N__41702\ : std_logic;
signal \N__41699\ : std_logic;
signal \N__41698\ : std_logic;
signal \N__41697\ : std_logic;
signal \N__41696\ : std_logic;
signal \N__41693\ : std_logic;
signal \N__41690\ : std_logic;
signal \N__41687\ : std_logic;
signal \N__41684\ : std_logic;
signal \N__41675\ : std_logic;
signal \N__41672\ : std_logic;
signal \N__41671\ : std_logic;
signal \N__41670\ : std_logic;
signal \N__41667\ : std_logic;
signal \N__41664\ : std_logic;
signal \N__41661\ : std_logic;
signal \N__41660\ : std_logic;
signal \N__41655\ : std_logic;
signal \N__41652\ : std_logic;
signal \N__41649\ : std_logic;
signal \N__41648\ : std_logic;
signal \N__41645\ : std_logic;
signal \N__41640\ : std_logic;
signal \N__41637\ : std_logic;
signal \N__41634\ : std_logic;
signal \N__41631\ : std_logic;
signal \N__41624\ : std_logic;
signal \N__41621\ : std_logic;
signal \N__41618\ : std_logic;
signal \N__41615\ : std_logic;
signal \N__41612\ : std_logic;
signal \N__41609\ : std_logic;
signal \N__41606\ : std_logic;
signal \N__41603\ : std_logic;
signal \N__41600\ : std_logic;
signal \N__41597\ : std_logic;
signal \N__41594\ : std_logic;
signal \N__41591\ : std_logic;
signal \N__41588\ : std_logic;
signal \N__41585\ : std_logic;
signal \N__41582\ : std_logic;
signal \N__41579\ : std_logic;
signal \N__41576\ : std_logic;
signal \N__41575\ : std_logic;
signal \N__41572\ : std_logic;
signal \N__41569\ : std_logic;
signal \N__41568\ : std_logic;
signal \N__41567\ : std_logic;
signal \N__41564\ : std_logic;
signal \N__41559\ : std_logic;
signal \N__41556\ : std_logic;
signal \N__41551\ : std_logic;
signal \N__41548\ : std_logic;
signal \N__41545\ : std_logic;
signal \N__41540\ : std_logic;
signal \N__41537\ : std_logic;
signal \N__41534\ : std_logic;
signal \N__41531\ : std_logic;
signal \N__41528\ : std_logic;
signal \N__41527\ : std_logic;
signal \N__41524\ : std_logic;
signal \N__41521\ : std_logic;
signal \N__41520\ : std_logic;
signal \N__41517\ : std_logic;
signal \N__41514\ : std_logic;
signal \N__41511\ : std_logic;
signal \N__41504\ : std_logic;
signal \N__41501\ : std_logic;
signal \N__41498\ : std_logic;
signal \N__41495\ : std_logic;
signal \N__41492\ : std_logic;
signal \N__41491\ : std_logic;
signal \N__41490\ : std_logic;
signal \N__41489\ : std_logic;
signal \N__41486\ : std_logic;
signal \N__41485\ : std_logic;
signal \N__41484\ : std_logic;
signal \N__41483\ : std_logic;
signal \N__41482\ : std_logic;
signal \N__41481\ : std_logic;
signal \N__41480\ : std_logic;
signal \N__41479\ : std_logic;
signal \N__41476\ : std_logic;
signal \N__41473\ : std_logic;
signal \N__41470\ : std_logic;
signal \N__41457\ : std_logic;
signal \N__41454\ : std_logic;
signal \N__41453\ : std_logic;
signal \N__41452\ : std_logic;
signal \N__41451\ : std_logic;
signal \N__41448\ : std_logic;
signal \N__41447\ : std_logic;
signal \N__41444\ : std_logic;
signal \N__41441\ : std_logic;
signal \N__41438\ : std_logic;
signal \N__41437\ : std_logic;
signal \N__41434\ : std_logic;
signal \N__41425\ : std_logic;
signal \N__41420\ : std_logic;
signal \N__41415\ : std_logic;
signal \N__41412\ : std_logic;
signal \N__41409\ : std_logic;
signal \N__41406\ : std_logic;
signal \N__41393\ : std_logic;
signal \N__41390\ : std_logic;
signal \N__41387\ : std_logic;
signal \N__41384\ : std_logic;
signal \N__41381\ : std_logic;
signal \N__41378\ : std_logic;
signal \N__41375\ : std_logic;
signal \N__41372\ : std_logic;
signal \N__41369\ : std_logic;
signal \N__41366\ : std_logic;
signal \N__41363\ : std_logic;
signal \N__41360\ : std_logic;
signal \N__41357\ : std_logic;
signal \N__41354\ : std_logic;
signal \N__41351\ : std_logic;
signal \N__41348\ : std_logic;
signal \N__41345\ : std_logic;
signal \N__41342\ : std_logic;
signal \N__41339\ : std_logic;
signal \N__41336\ : std_logic;
signal \N__41333\ : std_logic;
signal \N__41330\ : std_logic;
signal \N__41327\ : std_logic;
signal \N__41324\ : std_logic;
signal \N__41321\ : std_logic;
signal \N__41318\ : std_logic;
signal \N__41315\ : std_logic;
signal \N__41312\ : std_logic;
signal \N__41309\ : std_logic;
signal \N__41306\ : std_logic;
signal \N__41303\ : std_logic;
signal \N__41300\ : std_logic;
signal \N__41297\ : std_logic;
signal \N__41294\ : std_logic;
signal \N__41291\ : std_logic;
signal \N__41288\ : std_logic;
signal \N__41285\ : std_logic;
signal \N__41282\ : std_logic;
signal \N__41279\ : std_logic;
signal \N__41276\ : std_logic;
signal \N__41275\ : std_logic;
signal \N__41272\ : std_logic;
signal \N__41269\ : std_logic;
signal \N__41266\ : std_logic;
signal \N__41263\ : std_logic;
signal \N__41260\ : std_logic;
signal \N__41257\ : std_logic;
signal \N__41254\ : std_logic;
signal \N__41253\ : std_logic;
signal \N__41252\ : std_logic;
signal \N__41249\ : std_logic;
signal \N__41248\ : std_logic;
signal \N__41245\ : std_logic;
signal \N__41242\ : std_logic;
signal \N__41239\ : std_logic;
signal \N__41236\ : std_logic;
signal \N__41233\ : std_logic;
signal \N__41228\ : std_logic;
signal \N__41225\ : std_logic;
signal \N__41220\ : std_logic;
signal \N__41217\ : std_logic;
signal \N__41210\ : std_logic;
signal \N__41207\ : std_logic;
signal \N__41204\ : std_logic;
signal \N__41201\ : std_logic;
signal \N__41198\ : std_logic;
signal \N__41195\ : std_logic;
signal \N__41192\ : std_logic;
signal \N__41189\ : std_logic;
signal \N__41186\ : std_logic;
signal \N__41183\ : std_logic;
signal \N__41180\ : std_logic;
signal \N__41177\ : std_logic;
signal \N__41174\ : std_logic;
signal \N__41171\ : std_logic;
signal \N__41168\ : std_logic;
signal \N__41165\ : std_logic;
signal \N__41162\ : std_logic;
signal \N__41159\ : std_logic;
signal \N__41156\ : std_logic;
signal \N__41153\ : std_logic;
signal \N__41150\ : std_logic;
signal \N__41147\ : std_logic;
signal \N__41144\ : std_logic;
signal \N__41141\ : std_logic;
signal \N__41138\ : std_logic;
signal \N__41135\ : std_logic;
signal \N__41132\ : std_logic;
signal \N__41129\ : std_logic;
signal \N__41126\ : std_logic;
signal \N__41123\ : std_logic;
signal \N__41120\ : std_logic;
signal \N__41117\ : std_logic;
signal \N__41114\ : std_logic;
signal \N__41111\ : std_logic;
signal \N__41108\ : std_logic;
signal \N__41105\ : std_logic;
signal \N__41102\ : std_logic;
signal \N__41099\ : std_logic;
signal \N__41096\ : std_logic;
signal \N__41093\ : std_logic;
signal \N__41090\ : std_logic;
signal \N__41087\ : std_logic;
signal \N__41084\ : std_logic;
signal \N__41081\ : std_logic;
signal \N__41078\ : std_logic;
signal \N__41075\ : std_logic;
signal \N__41072\ : std_logic;
signal \N__41069\ : std_logic;
signal \N__41068\ : std_logic;
signal \N__41067\ : std_logic;
signal \N__41066\ : std_logic;
signal \N__41065\ : std_logic;
signal \N__41064\ : std_logic;
signal \N__41063\ : std_logic;
signal \N__41062\ : std_logic;
signal \N__41061\ : std_logic;
signal \N__41060\ : std_logic;
signal \N__41059\ : std_logic;
signal \N__41058\ : std_logic;
signal \N__41055\ : std_logic;
signal \N__41054\ : std_logic;
signal \N__41053\ : std_logic;
signal \N__41046\ : std_logic;
signal \N__41037\ : std_logic;
signal \N__41030\ : std_logic;
signal \N__41029\ : std_logic;
signal \N__41028\ : std_logic;
signal \N__41027\ : std_logic;
signal \N__41026\ : std_logic;
signal \N__41023\ : std_logic;
signal \N__41022\ : std_logic;
signal \N__41021\ : std_logic;
signal \N__41018\ : std_logic;
signal \N__41015\ : std_logic;
signal \N__41012\ : std_logic;
signal \N__41009\ : std_logic;
signal \N__41004\ : std_logic;
signal \N__41001\ : std_logic;
signal \N__41000\ : std_logic;
signal \N__40999\ : std_logic;
signal \N__40998\ : std_logic;
signal \N__40991\ : std_logic;
signal \N__40988\ : std_logic;
signal \N__40985\ : std_logic;
signal \N__40982\ : std_logic;
signal \N__40981\ : std_logic;
signal \N__40970\ : std_logic;
signal \N__40961\ : std_logic;
signal \N__40956\ : std_logic;
signal \N__40953\ : std_logic;
signal \N__40950\ : std_logic;
signal \N__40947\ : std_logic;
signal \N__40942\ : std_logic;
signal \N__40937\ : std_logic;
signal \N__40934\ : std_logic;
signal \N__40929\ : std_logic;
signal \N__40926\ : std_logic;
signal \N__40919\ : std_logic;
signal \N__40918\ : std_logic;
signal \N__40917\ : std_logic;
signal \N__40916\ : std_logic;
signal \N__40915\ : std_logic;
signal \N__40914\ : std_logic;
signal \N__40911\ : std_logic;
signal \N__40910\ : std_logic;
signal \N__40909\ : std_logic;
signal \N__40906\ : std_logic;
signal \N__40903\ : std_logic;
signal \N__40902\ : std_logic;
signal \N__40901\ : std_logic;
signal \N__40900\ : std_logic;
signal \N__40899\ : std_logic;
signal \N__40896\ : std_logic;
signal \N__40895\ : std_logic;
signal \N__40894\ : std_logic;
signal \N__40891\ : std_logic;
signal \N__40888\ : std_logic;
signal \N__40885\ : std_logic;
signal \N__40882\ : std_logic;
signal \N__40879\ : std_logic;
signal \N__40876\ : std_logic;
signal \N__40873\ : std_logic;
signal \N__40872\ : std_logic;
signal \N__40869\ : std_logic;
signal \N__40866\ : std_logic;
signal \N__40863\ : std_logic;
signal \N__40862\ : std_logic;
signal \N__40861\ : std_logic;
signal \N__40860\ : std_logic;
signal \N__40859\ : std_logic;
signal \N__40858\ : std_logic;
signal \N__40857\ : std_logic;
signal \N__40854\ : std_logic;
signal \N__40853\ : std_logic;
signal \N__40852\ : std_logic;
signal \N__40849\ : std_logic;
signal \N__40842\ : std_logic;
signal \N__40839\ : std_logic;
signal \N__40836\ : std_logic;
signal \N__40831\ : std_logic;
signal \N__40826\ : std_logic;
signal \N__40821\ : std_logic;
signal \N__40812\ : std_logic;
signal \N__40803\ : std_logic;
signal \N__40802\ : std_logic;
signal \N__40795\ : std_logic;
signal \N__40792\ : std_logic;
signal \N__40789\ : std_logic;
signal \N__40784\ : std_logic;
signal \N__40775\ : std_logic;
signal \N__40772\ : std_logic;
signal \N__40769\ : std_logic;
signal \N__40766\ : std_logic;
signal \N__40763\ : std_logic;
signal \N__40760\ : std_logic;
signal \N__40755\ : std_logic;
signal \N__40752\ : std_logic;
signal \N__40739\ : std_logic;
signal \N__40738\ : std_logic;
signal \N__40735\ : std_logic;
signal \N__40732\ : std_logic;
signal \N__40729\ : std_logic;
signal \N__40728\ : std_logic;
signal \N__40725\ : std_logic;
signal \N__40722\ : std_logic;
signal \N__40719\ : std_logic;
signal \N__40718\ : std_logic;
signal \N__40717\ : std_logic;
signal \N__40716\ : std_logic;
signal \N__40713\ : std_logic;
signal \N__40708\ : std_logic;
signal \N__40705\ : std_logic;
signal \N__40700\ : std_logic;
signal \N__40691\ : std_logic;
signal \N__40690\ : std_logic;
signal \N__40687\ : std_logic;
signal \N__40684\ : std_logic;
signal \N__40683\ : std_logic;
signal \N__40682\ : std_logic;
signal \N__40681\ : std_logic;
signal \N__40680\ : std_logic;
signal \N__40679\ : std_logic;
signal \N__40674\ : std_logic;
signal \N__40671\ : std_logic;
signal \N__40668\ : std_logic;
signal \N__40667\ : std_logic;
signal \N__40666\ : std_logic;
signal \N__40665\ : std_logic;
signal \N__40664\ : std_logic;
signal \N__40663\ : std_logic;
signal \N__40656\ : std_logic;
signal \N__40655\ : std_logic;
signal \N__40650\ : std_logic;
signal \N__40647\ : std_logic;
signal \N__40644\ : std_logic;
signal \N__40641\ : std_logic;
signal \N__40640\ : std_logic;
signal \N__40637\ : std_logic;
signal \N__40636\ : std_logic;
signal \N__40635\ : std_logic;
signal \N__40634\ : std_logic;
signal \N__40633\ : std_logic;
signal \N__40632\ : std_logic;
signal \N__40631\ : std_logic;
signal \N__40630\ : std_logic;
signal \N__40629\ : std_logic;
signal \N__40628\ : std_logic;
signal \N__40625\ : std_logic;
signal \N__40622\ : std_logic;
signal \N__40619\ : std_logic;
signal \N__40616\ : std_logic;
signal \N__40611\ : std_logic;
signal \N__40604\ : std_logic;
signal \N__40595\ : std_logic;
signal \N__40588\ : std_logic;
signal \N__40583\ : std_logic;
signal \N__40580\ : std_logic;
signal \N__40579\ : std_logic;
signal \N__40572\ : std_logic;
signal \N__40569\ : std_logic;
signal \N__40564\ : std_logic;
signal \N__40557\ : std_logic;
signal \N__40554\ : std_logic;
signal \N__40551\ : std_logic;
signal \N__40548\ : std_logic;
signal \N__40543\ : std_logic;
signal \N__40538\ : std_logic;
signal \N__40529\ : std_logic;
signal \N__40526\ : std_logic;
signal \N__40523\ : std_logic;
signal \N__40522\ : std_logic;
signal \N__40519\ : std_logic;
signal \N__40518\ : std_logic;
signal \N__40515\ : std_logic;
signal \N__40514\ : std_logic;
signal \N__40511\ : std_logic;
signal \N__40508\ : std_logic;
signal \N__40505\ : std_logic;
signal \N__40502\ : std_logic;
signal \N__40499\ : std_logic;
signal \N__40496\ : std_logic;
signal \N__40491\ : std_logic;
signal \N__40488\ : std_logic;
signal \N__40485\ : std_logic;
signal \N__40482\ : std_logic;
signal \N__40475\ : std_logic;
signal \N__40472\ : std_logic;
signal \N__40469\ : std_logic;
signal \N__40466\ : std_logic;
signal \N__40463\ : std_logic;
signal \N__40460\ : std_logic;
signal \N__40457\ : std_logic;
signal \N__40454\ : std_logic;
signal \N__40453\ : std_logic;
signal \N__40450\ : std_logic;
signal \N__40447\ : std_logic;
signal \N__40444\ : std_logic;
signal \N__40441\ : std_logic;
signal \N__40440\ : std_logic;
signal \N__40439\ : std_logic;
signal \N__40436\ : std_logic;
signal \N__40433\ : std_logic;
signal \N__40430\ : std_logic;
signal \N__40429\ : std_logic;
signal \N__40426\ : std_logic;
signal \N__40419\ : std_logic;
signal \N__40414\ : std_logic;
signal \N__40409\ : std_logic;
signal \N__40406\ : std_logic;
signal \N__40403\ : std_logic;
signal \N__40400\ : std_logic;
signal \N__40397\ : std_logic;
signal \N__40394\ : std_logic;
signal \N__40393\ : std_logic;
signal \N__40390\ : std_logic;
signal \N__40389\ : std_logic;
signal \N__40386\ : std_logic;
signal \N__40383\ : std_logic;
signal \N__40380\ : std_logic;
signal \N__40377\ : std_logic;
signal \N__40374\ : std_logic;
signal \N__40371\ : std_logic;
signal \N__40368\ : std_logic;
signal \N__40365\ : std_logic;
signal \N__40360\ : std_logic;
signal \N__40355\ : std_logic;
signal \N__40352\ : std_logic;
signal \N__40349\ : std_logic;
signal \N__40346\ : std_logic;
signal \N__40345\ : std_logic;
signal \N__40344\ : std_logic;
signal \N__40343\ : std_logic;
signal \N__40342\ : std_logic;
signal \N__40337\ : std_logic;
signal \N__40336\ : std_logic;
signal \N__40335\ : std_logic;
signal \N__40332\ : std_logic;
signal \N__40329\ : std_logic;
signal \N__40328\ : std_logic;
signal \N__40327\ : std_logic;
signal \N__40326\ : std_logic;
signal \N__40323\ : std_logic;
signal \N__40320\ : std_logic;
signal \N__40319\ : std_logic;
signal \N__40318\ : std_logic;
signal \N__40317\ : std_logic;
signal \N__40316\ : std_logic;
signal \N__40311\ : std_logic;
signal \N__40308\ : std_logic;
signal \N__40299\ : std_logic;
signal \N__40296\ : std_logic;
signal \N__40293\ : std_logic;
signal \N__40284\ : std_logic;
signal \N__40281\ : std_logic;
signal \N__40278\ : std_logic;
signal \N__40275\ : std_logic;
signal \N__40272\ : std_logic;
signal \N__40269\ : std_logic;
signal \N__40262\ : std_logic;
signal \N__40259\ : std_logic;
signal \N__40250\ : std_logic;
signal \N__40249\ : std_logic;
signal \N__40248\ : std_logic;
signal \N__40245\ : std_logic;
signal \N__40242\ : std_logic;
signal \N__40239\ : std_logic;
signal \N__40236\ : std_logic;
signal \N__40233\ : std_logic;
signal \N__40230\ : std_logic;
signal \N__40225\ : std_logic;
signal \N__40222\ : std_logic;
signal \N__40217\ : std_logic;
signal \N__40216\ : std_logic;
signal \N__40215\ : std_logic;
signal \N__40210\ : std_logic;
signal \N__40207\ : std_logic;
signal \N__40206\ : std_logic;
signal \N__40205\ : std_logic;
signal \N__40202\ : std_logic;
signal \N__40195\ : std_logic;
signal \N__40192\ : std_logic;
signal \N__40189\ : std_logic;
signal \N__40186\ : std_logic;
signal \N__40183\ : std_logic;
signal \N__40178\ : std_logic;
signal \N__40177\ : std_logic;
signal \N__40174\ : std_logic;
signal \N__40171\ : std_logic;
signal \N__40168\ : std_logic;
signal \N__40165\ : std_logic;
signal \N__40164\ : std_logic;
signal \N__40161\ : std_logic;
signal \N__40158\ : std_logic;
signal \N__40155\ : std_logic;
signal \N__40150\ : std_logic;
signal \N__40147\ : std_logic;
signal \N__40142\ : std_logic;
signal \N__40139\ : std_logic;
signal \N__40138\ : std_logic;
signal \N__40135\ : std_logic;
signal \N__40132\ : std_logic;
signal \N__40129\ : std_logic;
signal \N__40126\ : std_logic;
signal \N__40121\ : std_logic;
signal \N__40118\ : std_logic;
signal \N__40117\ : std_logic;
signal \N__40114\ : std_logic;
signal \N__40111\ : std_logic;
signal \N__40108\ : std_logic;
signal \N__40105\ : std_logic;
signal \N__40102\ : std_logic;
signal \N__40099\ : std_logic;
signal \N__40094\ : std_logic;
signal \N__40093\ : std_logic;
signal \N__40092\ : std_logic;
signal \N__40089\ : std_logic;
signal \N__40084\ : std_logic;
signal \N__40081\ : std_logic;
signal \N__40078\ : std_logic;
signal \N__40075\ : std_logic;
signal \N__40072\ : std_logic;
signal \N__40067\ : std_logic;
signal \N__40066\ : std_logic;
signal \N__40065\ : std_logic;
signal \N__40064\ : std_logic;
signal \N__40061\ : std_logic;
signal \N__40056\ : std_logic;
signal \N__40053\ : std_logic;
signal \N__40050\ : std_logic;
signal \N__40047\ : std_logic;
signal \N__40044\ : std_logic;
signal \N__40041\ : std_logic;
signal \N__40040\ : std_logic;
signal \N__40039\ : std_logic;
signal \N__40036\ : std_logic;
signal \N__40031\ : std_logic;
signal \N__40026\ : std_logic;
signal \N__40019\ : std_logic;
signal \N__40018\ : std_logic;
signal \N__40017\ : std_logic;
signal \N__40016\ : std_logic;
signal \N__40015\ : std_logic;
signal \N__40014\ : std_logic;
signal \N__40013\ : std_logic;
signal \N__40012\ : std_logic;
signal \N__40011\ : std_logic;
signal \N__40008\ : std_logic;
signal \N__40007\ : std_logic;
signal \N__40006\ : std_logic;
signal \N__40003\ : std_logic;
signal \N__40002\ : std_logic;
signal \N__40001\ : std_logic;
signal \N__39998\ : std_logic;
signal \N__39995\ : std_logic;
signal \N__39994\ : std_logic;
signal \N__39991\ : std_logic;
signal \N__39990\ : std_logic;
signal \N__39989\ : std_logic;
signal \N__39988\ : std_logic;
signal \N__39985\ : std_logic;
signal \N__39982\ : std_logic;
signal \N__39979\ : std_logic;
signal \N__39978\ : std_logic;
signal \N__39977\ : std_logic;
signal \N__39972\ : std_logic;
signal \N__39969\ : std_logic;
signal \N__39966\ : std_logic;
signal \N__39963\ : std_logic;
signal \N__39962\ : std_logic;
signal \N__39961\ : std_logic;
signal \N__39946\ : std_logic;
signal \N__39933\ : std_logic;
signal \N__39932\ : std_logic;
signal \N__39929\ : std_logic;
signal \N__39928\ : std_logic;
signal \N__39925\ : std_logic;
signal \N__39920\ : std_logic;
signal \N__39917\ : std_logic;
signal \N__39914\ : std_logic;
signal \N__39911\ : std_logic;
signal \N__39910\ : std_logic;
signal \N__39907\ : std_logic;
signal \N__39904\ : std_logic;
signal \N__39899\ : std_logic;
signal \N__39896\ : std_logic;
signal \N__39893\ : std_logic;
signal \N__39890\ : std_logic;
signal \N__39883\ : std_logic;
signal \N__39880\ : std_logic;
signal \N__39873\ : std_logic;
signal \N__39870\ : std_logic;
signal \N__39863\ : std_logic;
signal \N__39854\ : std_logic;
signal \N__39853\ : std_logic;
signal \N__39852\ : std_logic;
signal \N__39851\ : std_logic;
signal \N__39850\ : std_logic;
signal \N__39849\ : std_logic;
signal \N__39848\ : std_logic;
signal \N__39847\ : std_logic;
signal \N__39846\ : std_logic;
signal \N__39845\ : std_logic;
signal \N__39842\ : std_logic;
signal \N__39839\ : std_logic;
signal \N__39836\ : std_logic;
signal \N__39833\ : std_logic;
signal \N__39830\ : std_logic;
signal \N__39827\ : std_logic;
signal \N__39824\ : std_logic;
signal \N__39823\ : std_logic;
signal \N__39822\ : std_logic;
signal \N__39821\ : std_logic;
signal \N__39820\ : std_logic;
signal \N__39819\ : std_logic;
signal \N__39818\ : std_logic;
signal \N__39813\ : std_logic;
signal \N__39812\ : std_logic;
signal \N__39811\ : std_logic;
signal \N__39808\ : std_logic;
signal \N__39799\ : std_logic;
signal \N__39792\ : std_logic;
signal \N__39785\ : std_logic;
signal \N__39778\ : std_logic;
signal \N__39775\ : std_logic;
signal \N__39770\ : std_logic;
signal \N__39769\ : std_logic;
signal \N__39768\ : std_logic;
signal \N__39767\ : std_logic;
signal \N__39766\ : std_logic;
signal \N__39755\ : std_logic;
signal \N__39750\ : std_logic;
signal \N__39747\ : std_logic;
signal \N__39744\ : std_logic;
signal \N__39739\ : std_logic;
signal \N__39738\ : std_logic;
signal \N__39735\ : std_logic;
signal \N__39732\ : std_logic;
signal \N__39729\ : std_logic;
signal \N__39726\ : std_logic;
signal \N__39723\ : std_logic;
signal \N__39720\ : std_logic;
signal \N__39719\ : std_logic;
signal \N__39716\ : std_logic;
signal \N__39713\ : std_logic;
signal \N__39710\ : std_logic;
signal \N__39705\ : std_logic;
signal \N__39700\ : std_logic;
signal \N__39697\ : std_logic;
signal \N__39694\ : std_logic;
signal \N__39689\ : std_logic;
signal \N__39680\ : std_logic;
signal \N__39679\ : std_logic;
signal \N__39678\ : std_logic;
signal \N__39675\ : std_logic;
signal \N__39670\ : std_logic;
signal \N__39669\ : std_logic;
signal \N__39668\ : std_logic;
signal \N__39667\ : std_logic;
signal \N__39666\ : std_logic;
signal \N__39665\ : std_logic;
signal \N__39664\ : std_logic;
signal \N__39663\ : std_logic;
signal \N__39662\ : std_logic;
signal \N__39661\ : std_logic;
signal \N__39660\ : std_logic;
signal \N__39659\ : std_logic;
signal \N__39658\ : std_logic;
signal \N__39657\ : std_logic;
signal \N__39656\ : std_logic;
signal \N__39655\ : std_logic;
signal \N__39654\ : std_logic;
signal \N__39651\ : std_logic;
signal \N__39648\ : std_logic;
signal \N__39645\ : std_logic;
signal \N__39642\ : std_logic;
signal \N__39629\ : std_logic;
signal \N__39614\ : std_logic;
signal \N__39611\ : std_logic;
signal \N__39610\ : std_logic;
signal \N__39609\ : std_logic;
signal \N__39608\ : std_logic;
signal \N__39601\ : std_logic;
signal \N__39594\ : std_logic;
signal \N__39591\ : std_logic;
signal \N__39588\ : std_logic;
signal \N__39583\ : std_logic;
signal \N__39580\ : std_logic;
signal \N__39577\ : std_logic;
signal \N__39570\ : std_logic;
signal \N__39569\ : std_logic;
signal \N__39568\ : std_logic;
signal \N__39565\ : std_logic;
signal \N__39562\ : std_logic;
signal \N__39559\ : std_logic;
signal \N__39554\ : std_logic;
signal \N__39551\ : std_logic;
signal \N__39548\ : std_logic;
signal \N__39545\ : std_logic;
signal \N__39536\ : std_logic;
signal \N__39535\ : std_logic;
signal \N__39532\ : std_logic;
signal \N__39529\ : std_logic;
signal \N__39524\ : std_logic;
signal \N__39521\ : std_logic;
signal \N__39518\ : std_logic;
signal \N__39515\ : std_logic;
signal \N__39514\ : std_logic;
signal \N__39513\ : std_logic;
signal \N__39512\ : std_logic;
signal \N__39503\ : std_logic;
signal \N__39500\ : std_logic;
signal \N__39497\ : std_logic;
signal \N__39496\ : std_logic;
signal \N__39493\ : std_logic;
signal \N__39490\ : std_logic;
signal \N__39489\ : std_logic;
signal \N__39486\ : std_logic;
signal \N__39483\ : std_logic;
signal \N__39480\ : std_logic;
signal \N__39473\ : std_logic;
signal \N__39470\ : std_logic;
signal \N__39469\ : std_logic;
signal \N__39466\ : std_logic;
signal \N__39463\ : std_logic;
signal \N__39462\ : std_logic;
signal \N__39459\ : std_logic;
signal \N__39456\ : std_logic;
signal \N__39453\ : std_logic;
signal \N__39446\ : std_logic;
signal \N__39443\ : std_logic;
signal \N__39440\ : std_logic;
signal \N__39437\ : std_logic;
signal \N__39434\ : std_logic;
signal \N__39431\ : std_logic;
signal \N__39428\ : std_logic;
signal \N__39425\ : std_logic;
signal \N__39422\ : std_logic;
signal \N__39419\ : std_logic;
signal \N__39416\ : std_logic;
signal \N__39413\ : std_logic;
signal \N__39410\ : std_logic;
signal \N__39407\ : std_logic;
signal \N__39406\ : std_logic;
signal \N__39405\ : std_logic;
signal \N__39402\ : std_logic;
signal \N__39401\ : std_logic;
signal \N__39398\ : std_logic;
signal \N__39395\ : std_logic;
signal \N__39392\ : std_logic;
signal \N__39389\ : std_logic;
signal \N__39386\ : std_logic;
signal \N__39383\ : std_logic;
signal \N__39380\ : std_logic;
signal \N__39379\ : std_logic;
signal \N__39376\ : std_logic;
signal \N__39373\ : std_logic;
signal \N__39368\ : std_logic;
signal \N__39365\ : std_logic;
signal \N__39362\ : std_logic;
signal \N__39353\ : std_logic;
signal \N__39352\ : std_logic;
signal \N__39351\ : std_logic;
signal \N__39350\ : std_logic;
signal \N__39347\ : std_logic;
signal \N__39344\ : std_logic;
signal \N__39341\ : std_logic;
signal \N__39338\ : std_logic;
signal \N__39335\ : std_logic;
signal \N__39332\ : std_logic;
signal \N__39331\ : std_logic;
signal \N__39328\ : std_logic;
signal \N__39325\ : std_logic;
signal \N__39322\ : std_logic;
signal \N__39319\ : std_logic;
signal \N__39316\ : std_logic;
signal \N__39313\ : std_logic;
signal \N__39302\ : std_logic;
signal \N__39299\ : std_logic;
signal \N__39296\ : std_logic;
signal \N__39293\ : std_logic;
signal \N__39290\ : std_logic;
signal \N__39287\ : std_logic;
signal \N__39284\ : std_logic;
signal \N__39281\ : std_logic;
signal \N__39278\ : std_logic;
signal \N__39275\ : std_logic;
signal \N__39272\ : std_logic;
signal \N__39269\ : std_logic;
signal \N__39266\ : std_logic;
signal \N__39263\ : std_logic;
signal \N__39260\ : std_logic;
signal \N__39259\ : std_logic;
signal \N__39256\ : std_logic;
signal \N__39255\ : std_logic;
signal \N__39254\ : std_logic;
signal \N__39251\ : std_logic;
signal \N__39248\ : std_logic;
signal \N__39243\ : std_logic;
signal \N__39240\ : std_logic;
signal \N__39233\ : std_logic;
signal \N__39232\ : std_logic;
signal \N__39231\ : std_logic;
signal \N__39228\ : std_logic;
signal \N__39225\ : std_logic;
signal \N__39222\ : std_logic;
signal \N__39217\ : std_logic;
signal \N__39212\ : std_logic;
signal \N__39209\ : std_logic;
signal \N__39208\ : std_logic;
signal \N__39207\ : std_logic;
signal \N__39204\ : std_logic;
signal \N__39201\ : std_logic;
signal \N__39198\ : std_logic;
signal \N__39193\ : std_logic;
signal \N__39188\ : std_logic;
signal \N__39185\ : std_logic;
signal \N__39184\ : std_logic;
signal \N__39183\ : std_logic;
signal \N__39180\ : std_logic;
signal \N__39177\ : std_logic;
signal \N__39174\ : std_logic;
signal \N__39171\ : std_logic;
signal \N__39164\ : std_logic;
signal \N__39161\ : std_logic;
signal \N__39160\ : std_logic;
signal \N__39159\ : std_logic;
signal \N__39156\ : std_logic;
signal \N__39153\ : std_logic;
signal \N__39150\ : std_logic;
signal \N__39147\ : std_logic;
signal \N__39140\ : std_logic;
signal \N__39137\ : std_logic;
signal \N__39136\ : std_logic;
signal \N__39135\ : std_logic;
signal \N__39132\ : std_logic;
signal \N__39129\ : std_logic;
signal \N__39126\ : std_logic;
signal \N__39121\ : std_logic;
signal \N__39116\ : std_logic;
signal \N__39113\ : std_logic;
signal \N__39112\ : std_logic;
signal \N__39111\ : std_logic;
signal \N__39108\ : std_logic;
signal \N__39105\ : std_logic;
signal \N__39102\ : std_logic;
signal \N__39097\ : std_logic;
signal \N__39092\ : std_logic;
signal \N__39089\ : std_logic;
signal \N__39088\ : std_logic;
signal \N__39085\ : std_logic;
signal \N__39082\ : std_logic;
signal \N__39077\ : std_logic;
signal \N__39074\ : std_logic;
signal \N__39073\ : std_logic;
signal \N__39072\ : std_logic;
signal \N__39071\ : std_logic;
signal \N__39070\ : std_logic;
signal \N__39069\ : std_logic;
signal \N__39068\ : std_logic;
signal \N__39067\ : std_logic;
signal \N__39066\ : std_logic;
signal \N__39065\ : std_logic;
signal \N__39064\ : std_logic;
signal \N__39063\ : std_logic;
signal \N__39062\ : std_logic;
signal \N__39061\ : std_logic;
signal \N__39060\ : std_logic;
signal \N__39059\ : std_logic;
signal \N__39058\ : std_logic;
signal \N__39057\ : std_logic;
signal \N__39056\ : std_logic;
signal \N__39055\ : std_logic;
signal \N__39054\ : std_logic;
signal \N__39053\ : std_logic;
signal \N__39052\ : std_logic;
signal \N__39051\ : std_logic;
signal \N__39050\ : std_logic;
signal \N__39049\ : std_logic;
signal \N__39044\ : std_logic;
signal \N__39035\ : std_logic;
signal \N__39034\ : std_logic;
signal \N__39033\ : std_logic;
signal \N__39032\ : std_logic;
signal \N__39031\ : std_logic;
signal \N__39022\ : std_logic;
signal \N__39013\ : std_logic;
signal \N__39004\ : std_logic;
signal \N__38995\ : std_logic;
signal \N__38986\ : std_logic;
signal \N__38983\ : std_logic;
signal \N__38980\ : std_logic;
signal \N__38971\ : std_logic;
signal \N__38962\ : std_logic;
signal \N__38959\ : std_logic;
signal \N__38956\ : std_logic;
signal \N__38953\ : std_logic;
signal \N__38948\ : std_logic;
signal \N__38939\ : std_logic;
signal \N__38936\ : std_logic;
signal \N__38935\ : std_logic;
signal \N__38932\ : std_logic;
signal \N__38929\ : std_logic;
signal \N__38924\ : std_logic;
signal \N__38921\ : std_logic;
signal \N__38918\ : std_logic;
signal \N__38917\ : std_logic;
signal \N__38916\ : std_logic;
signal \N__38913\ : std_logic;
signal \N__38910\ : std_logic;
signal \N__38909\ : std_logic;
signal \N__38906\ : std_logic;
signal \N__38901\ : std_logic;
signal \N__38898\ : std_logic;
signal \N__38895\ : std_logic;
signal \N__38890\ : std_logic;
signal \N__38887\ : std_logic;
signal \N__38884\ : std_logic;
signal \N__38879\ : std_logic;
signal \N__38878\ : std_logic;
signal \N__38877\ : std_logic;
signal \N__38874\ : std_logic;
signal \N__38871\ : std_logic;
signal \N__38868\ : std_logic;
signal \N__38863\ : std_logic;
signal \N__38858\ : std_logic;
signal \N__38855\ : std_logic;
signal \N__38854\ : std_logic;
signal \N__38853\ : std_logic;
signal \N__38850\ : std_logic;
signal \N__38847\ : std_logic;
signal \N__38844\ : std_logic;
signal \N__38839\ : std_logic;
signal \N__38834\ : std_logic;
signal \N__38831\ : std_logic;
signal \N__38830\ : std_logic;
signal \N__38829\ : std_logic;
signal \N__38826\ : std_logic;
signal \N__38823\ : std_logic;
signal \N__38820\ : std_logic;
signal \N__38817\ : std_logic;
signal \N__38810\ : std_logic;
signal \N__38807\ : std_logic;
signal \N__38806\ : std_logic;
signal \N__38805\ : std_logic;
signal \N__38802\ : std_logic;
signal \N__38799\ : std_logic;
signal \N__38796\ : std_logic;
signal \N__38793\ : std_logic;
signal \N__38786\ : std_logic;
signal \N__38783\ : std_logic;
signal \N__38782\ : std_logic;
signal \N__38781\ : std_logic;
signal \N__38778\ : std_logic;
signal \N__38775\ : std_logic;
signal \N__38772\ : std_logic;
signal \N__38767\ : std_logic;
signal \N__38762\ : std_logic;
signal \N__38759\ : std_logic;
signal \N__38758\ : std_logic;
signal \N__38757\ : std_logic;
signal \N__38754\ : std_logic;
signal \N__38751\ : std_logic;
signal \N__38748\ : std_logic;
signal \N__38743\ : std_logic;
signal \N__38738\ : std_logic;
signal \N__38735\ : std_logic;
signal \N__38734\ : std_logic;
signal \N__38733\ : std_logic;
signal \N__38730\ : std_logic;
signal \N__38725\ : std_logic;
signal \N__38720\ : std_logic;
signal \N__38717\ : std_logic;
signal \N__38716\ : std_logic;
signal \N__38715\ : std_logic;
signal \N__38712\ : std_logic;
signal \N__38707\ : std_logic;
signal \N__38702\ : std_logic;
signal \N__38699\ : std_logic;
signal \N__38698\ : std_logic;
signal \N__38697\ : std_logic;
signal \N__38694\ : std_logic;
signal \N__38691\ : std_logic;
signal \N__38688\ : std_logic;
signal \N__38683\ : std_logic;
signal \N__38678\ : std_logic;
signal \N__38675\ : std_logic;
signal \N__38674\ : std_logic;
signal \N__38673\ : std_logic;
signal \N__38670\ : std_logic;
signal \N__38667\ : std_logic;
signal \N__38664\ : std_logic;
signal \N__38659\ : std_logic;
signal \N__38654\ : std_logic;
signal \N__38651\ : std_logic;
signal \N__38650\ : std_logic;
signal \N__38649\ : std_logic;
signal \N__38646\ : std_logic;
signal \N__38643\ : std_logic;
signal \N__38640\ : std_logic;
signal \N__38637\ : std_logic;
signal \N__38630\ : std_logic;
signal \N__38627\ : std_logic;
signal \N__38626\ : std_logic;
signal \N__38625\ : std_logic;
signal \N__38622\ : std_logic;
signal \N__38619\ : std_logic;
signal \N__38616\ : std_logic;
signal \N__38613\ : std_logic;
signal \N__38606\ : std_logic;
signal \N__38603\ : std_logic;
signal \N__38602\ : std_logic;
signal \N__38601\ : std_logic;
signal \N__38598\ : std_logic;
signal \N__38595\ : std_logic;
signal \N__38592\ : std_logic;
signal \N__38587\ : std_logic;
signal \N__38582\ : std_logic;
signal \N__38579\ : std_logic;
signal \N__38578\ : std_logic;
signal \N__38577\ : std_logic;
signal \N__38574\ : std_logic;
signal \N__38571\ : std_logic;
signal \N__38568\ : std_logic;
signal \N__38563\ : std_logic;
signal \N__38558\ : std_logic;
signal \N__38555\ : std_logic;
signal \N__38554\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38550\ : std_logic;
signal \N__38545\ : std_logic;
signal \N__38540\ : std_logic;
signal \N__38537\ : std_logic;
signal \N__38536\ : std_logic;
signal \N__38535\ : std_logic;
signal \N__38532\ : std_logic;
signal \N__38527\ : std_logic;
signal \N__38522\ : std_logic;
signal \N__38519\ : std_logic;
signal \N__38516\ : std_logic;
signal \N__38513\ : std_logic;
signal \N__38510\ : std_logic;
signal \N__38509\ : std_logic;
signal \N__38506\ : std_logic;
signal \N__38503\ : std_logic;
signal \N__38500\ : std_logic;
signal \N__38497\ : std_logic;
signal \N__38494\ : std_logic;
signal \N__38489\ : std_logic;
signal \N__38486\ : std_logic;
signal \N__38483\ : std_logic;
signal \N__38480\ : std_logic;
signal \N__38477\ : std_logic;
signal \N__38476\ : std_logic;
signal \N__38473\ : std_logic;
signal \N__38470\ : std_logic;
signal \N__38467\ : std_logic;
signal \N__38464\ : std_logic;
signal \N__38461\ : std_logic;
signal \N__38456\ : std_logic;
signal \N__38455\ : std_logic;
signal \N__38454\ : std_logic;
signal \N__38451\ : std_logic;
signal \N__38448\ : std_logic;
signal \N__38445\ : std_logic;
signal \N__38438\ : std_logic;
signal \N__38435\ : std_logic;
signal \N__38434\ : std_logic;
signal \N__38433\ : std_logic;
signal \N__38430\ : std_logic;
signal \N__38427\ : std_logic;
signal \N__38424\ : std_logic;
signal \N__38417\ : std_logic;
signal \N__38414\ : std_logic;
signal \N__38413\ : std_logic;
signal \N__38412\ : std_logic;
signal \N__38409\ : std_logic;
signal \N__38406\ : std_logic;
signal \N__38403\ : std_logic;
signal \N__38398\ : std_logic;
signal \N__38393\ : std_logic;
signal \N__38390\ : std_logic;
signal \N__38389\ : std_logic;
signal \N__38388\ : std_logic;
signal \N__38385\ : std_logic;
signal \N__38382\ : std_logic;
signal \N__38379\ : std_logic;
signal \N__38374\ : std_logic;
signal \N__38369\ : std_logic;
signal \N__38366\ : std_logic;
signal \N__38365\ : std_logic;
signal \N__38364\ : std_logic;
signal \N__38361\ : std_logic;
signal \N__38356\ : std_logic;
signal \N__38351\ : std_logic;
signal \N__38348\ : std_logic;
signal \N__38347\ : std_logic;
signal \N__38346\ : std_logic;
signal \N__38343\ : std_logic;
signal \N__38338\ : std_logic;
signal \N__38333\ : std_logic;
signal \N__38330\ : std_logic;
signal \N__38327\ : std_logic;
signal \N__38324\ : std_logic;
signal \N__38321\ : std_logic;
signal \N__38320\ : std_logic;
signal \N__38317\ : std_logic;
signal \N__38314\ : std_logic;
signal \N__38311\ : std_logic;
signal \N__38306\ : std_logic;
signal \N__38303\ : std_logic;
signal \N__38300\ : std_logic;
signal \N__38297\ : std_logic;
signal \N__38294\ : std_logic;
signal \N__38291\ : std_logic;
signal \N__38288\ : std_logic;
signal \N__38287\ : std_logic;
signal \N__38286\ : std_logic;
signal \N__38283\ : std_logic;
signal \N__38280\ : std_logic;
signal \N__38277\ : std_logic;
signal \N__38274\ : std_logic;
signal \N__38269\ : std_logic;
signal \N__38264\ : std_logic;
signal \N__38261\ : std_logic;
signal \N__38258\ : std_logic;
signal \N__38255\ : std_logic;
signal \N__38252\ : std_logic;
signal \N__38251\ : std_logic;
signal \N__38248\ : std_logic;
signal \N__38245\ : std_logic;
signal \N__38242\ : std_logic;
signal \N__38239\ : std_logic;
signal \N__38234\ : std_logic;
signal \N__38231\ : std_logic;
signal \N__38228\ : std_logic;
signal \N__38225\ : std_logic;
signal \N__38222\ : std_logic;
signal \N__38219\ : std_logic;
signal \N__38218\ : std_logic;
signal \N__38215\ : std_logic;
signal \N__38212\ : std_logic;
signal \N__38209\ : std_logic;
signal \N__38204\ : std_logic;
signal \N__38201\ : std_logic;
signal \N__38198\ : std_logic;
signal \N__38195\ : std_logic;
signal \N__38194\ : std_logic;
signal \N__38191\ : std_logic;
signal \N__38188\ : std_logic;
signal \N__38185\ : std_logic;
signal \N__38180\ : std_logic;
signal \N__38179\ : std_logic;
signal \N__38178\ : std_logic;
signal \N__38177\ : std_logic;
signal \N__38176\ : std_logic;
signal \N__38175\ : std_logic;
signal \N__38174\ : std_logic;
signal \N__38173\ : std_logic;
signal \N__38170\ : std_logic;
signal \N__38167\ : std_logic;
signal \N__38166\ : std_logic;
signal \N__38165\ : std_logic;
signal \N__38164\ : std_logic;
signal \N__38163\ : std_logic;
signal \N__38162\ : std_logic;
signal \N__38161\ : std_logic;
signal \N__38160\ : std_logic;
signal \N__38159\ : std_logic;
signal \N__38148\ : std_logic;
signal \N__38147\ : std_logic;
signal \N__38146\ : std_logic;
signal \N__38145\ : std_logic;
signal \N__38144\ : std_logic;
signal \N__38143\ : std_logic;
signal \N__38142\ : std_logic;
signal \N__38127\ : std_logic;
signal \N__38118\ : std_logic;
signal \N__38117\ : std_logic;
signal \N__38114\ : std_logic;
signal \N__38107\ : std_logic;
signal \N__38104\ : std_logic;
signal \N__38103\ : std_logic;
signal \N__38098\ : std_logic;
signal \N__38093\ : std_logic;
signal \N__38090\ : std_logic;
signal \N__38085\ : std_logic;
signal \N__38080\ : std_logic;
signal \N__38075\ : std_logic;
signal \N__38072\ : std_logic;
signal \N__38069\ : std_logic;
signal \N__38064\ : std_logic;
signal \N__38061\ : std_logic;
signal \N__38058\ : std_logic;
signal \N__38051\ : std_logic;
signal \N__38050\ : std_logic;
signal \N__38049\ : std_logic;
signal \N__38048\ : std_logic;
signal \N__38047\ : std_logic;
signal \N__38046\ : std_logic;
signal \N__38045\ : std_logic;
signal \N__38044\ : std_logic;
signal \N__38043\ : std_logic;
signal \N__38040\ : std_logic;
signal \N__38039\ : std_logic;
signal \N__38038\ : std_logic;
signal \N__38037\ : std_logic;
signal \N__38034\ : std_logic;
signal \N__38031\ : std_logic;
signal \N__38028\ : std_logic;
signal \N__38025\ : std_logic;
signal \N__38024\ : std_logic;
signal \N__38023\ : std_logic;
signal \N__38022\ : std_logic;
signal \N__38019\ : std_logic;
signal \N__38018\ : std_logic;
signal \N__38017\ : std_logic;
signal \N__38016\ : std_logic;
signal \N__38015\ : std_logic;
signal \N__38012\ : std_logic;
signal \N__38009\ : std_logic;
signal \N__38006\ : std_logic;
signal \N__38005\ : std_logic;
signal \N__38004\ : std_logic;
signal \N__37999\ : std_logic;
signal \N__37998\ : std_logic;
signal \N__37987\ : std_logic;
signal \N__37982\ : std_logic;
signal \N__37967\ : std_logic;
signal \N__37964\ : std_logic;
signal \N__37955\ : std_logic;
signal \N__37952\ : std_logic;
signal \N__37951\ : std_logic;
signal \N__37948\ : std_logic;
signal \N__37947\ : std_logic;
signal \N__37944\ : std_logic;
signal \N__37937\ : std_logic;
signal \N__37934\ : std_logic;
signal \N__37931\ : std_logic;
signal \N__37924\ : std_logic;
signal \N__37919\ : std_logic;
signal \N__37910\ : std_logic;
signal \N__37907\ : std_logic;
signal \N__37904\ : std_logic;
signal \N__37901\ : std_logic;
signal \N__37900\ : std_logic;
signal \N__37899\ : std_logic;
signal \N__37898\ : std_logic;
signal \N__37897\ : std_logic;
signal \N__37896\ : std_logic;
signal \N__37895\ : std_logic;
signal \N__37894\ : std_logic;
signal \N__37893\ : std_logic;
signal \N__37892\ : std_logic;
signal \N__37889\ : std_logic;
signal \N__37886\ : std_logic;
signal \N__37885\ : std_logic;
signal \N__37884\ : std_logic;
signal \N__37881\ : std_logic;
signal \N__37878\ : std_logic;
signal \N__37877\ : std_logic;
signal \N__37876\ : std_logic;
signal \N__37875\ : std_logic;
signal \N__37874\ : std_logic;
signal \N__37873\ : std_logic;
signal \N__37862\ : std_logic;
signal \N__37861\ : std_logic;
signal \N__37860\ : std_logic;
signal \N__37859\ : std_logic;
signal \N__37858\ : std_logic;
signal \N__37855\ : std_logic;
signal \N__37850\ : std_logic;
signal \N__37845\ : std_logic;
signal \N__37830\ : std_logic;
signal \N__37827\ : std_logic;
signal \N__37826\ : std_logic;
signal \N__37823\ : std_logic;
signal \N__37818\ : std_logic;
signal \N__37815\ : std_logic;
signal \N__37812\ : std_logic;
signal \N__37803\ : std_logic;
signal \N__37800\ : std_logic;
signal \N__37795\ : std_logic;
signal \N__37794\ : std_logic;
signal \N__37793\ : std_logic;
signal \N__37786\ : std_logic;
signal \N__37783\ : std_logic;
signal \N__37780\ : std_logic;
signal \N__37775\ : std_logic;
signal \N__37770\ : std_logic;
signal \N__37767\ : std_logic;
signal \N__37760\ : std_logic;
signal \N__37757\ : std_logic;
signal \N__37756\ : std_logic;
signal \N__37753\ : std_logic;
signal \N__37750\ : std_logic;
signal \N__37747\ : std_logic;
signal \N__37742\ : std_logic;
signal \N__37739\ : std_logic;
signal \N__37736\ : std_logic;
signal \N__37733\ : std_logic;
signal \N__37732\ : std_logic;
signal \N__37729\ : std_logic;
signal \N__37726\ : std_logic;
signal \N__37723\ : std_logic;
signal \N__37720\ : std_logic;
signal \N__37715\ : std_logic;
signal \N__37712\ : std_logic;
signal \N__37709\ : std_logic;
signal \N__37706\ : std_logic;
signal \N__37705\ : std_logic;
signal \N__37702\ : std_logic;
signal \N__37699\ : std_logic;
signal \N__37696\ : std_logic;
signal \N__37693\ : std_logic;
signal \N__37690\ : std_logic;
signal \N__37685\ : std_logic;
signal \N__37682\ : std_logic;
signal \N__37679\ : std_logic;
signal \N__37676\ : std_logic;
signal \N__37675\ : std_logic;
signal \N__37672\ : std_logic;
signal \N__37669\ : std_logic;
signal \N__37666\ : std_logic;
signal \N__37661\ : std_logic;
signal \N__37658\ : std_logic;
signal \N__37655\ : std_logic;
signal \N__37652\ : std_logic;
signal \N__37651\ : std_logic;
signal \N__37648\ : std_logic;
signal \N__37645\ : std_logic;
signal \N__37642\ : std_logic;
signal \N__37637\ : std_logic;
signal \N__37634\ : std_logic;
signal \N__37631\ : std_logic;
signal \N__37628\ : std_logic;
signal \N__37627\ : std_logic;
signal \N__37624\ : std_logic;
signal \N__37621\ : std_logic;
signal \N__37618\ : std_logic;
signal \N__37613\ : std_logic;
signal \N__37610\ : std_logic;
signal \N__37607\ : std_logic;
signal \N__37604\ : std_logic;
signal \N__37601\ : std_logic;
signal \N__37598\ : std_logic;
signal \N__37597\ : std_logic;
signal \N__37594\ : std_logic;
signal \N__37591\ : std_logic;
signal \N__37588\ : std_logic;
signal \N__37585\ : std_logic;
signal \N__37580\ : std_logic;
signal \N__37577\ : std_logic;
signal \N__37574\ : std_logic;
signal \N__37571\ : std_logic;
signal \N__37568\ : std_logic;
signal \N__37565\ : std_logic;
signal \N__37564\ : std_logic;
signal \N__37561\ : std_logic;
signal \N__37558\ : std_logic;
signal \N__37555\ : std_logic;
signal \N__37552\ : std_logic;
signal \N__37547\ : std_logic;
signal \N__37544\ : std_logic;
signal \N__37541\ : std_logic;
signal \N__37538\ : std_logic;
signal \N__37537\ : std_logic;
signal \N__37534\ : std_logic;
signal \N__37531\ : std_logic;
signal \N__37528\ : std_logic;
signal \N__37523\ : std_logic;
signal \N__37520\ : std_logic;
signal \N__37517\ : std_logic;
signal \N__37514\ : std_logic;
signal \N__37513\ : std_logic;
signal \N__37510\ : std_logic;
signal \N__37507\ : std_logic;
signal \N__37504\ : std_logic;
signal \N__37499\ : std_logic;
signal \N__37496\ : std_logic;
signal \N__37493\ : std_logic;
signal \N__37490\ : std_logic;
signal \N__37487\ : std_logic;
signal \N__37486\ : std_logic;
signal \N__37483\ : std_logic;
signal \N__37480\ : std_logic;
signal \N__37477\ : std_logic;
signal \N__37474\ : std_logic;
signal \N__37469\ : std_logic;
signal \N__37466\ : std_logic;
signal \N__37465\ : std_logic;
signal \N__37464\ : std_logic;
signal \N__37457\ : std_logic;
signal \N__37456\ : std_logic;
signal \N__37455\ : std_logic;
signal \N__37454\ : std_logic;
signal \N__37451\ : std_logic;
signal \N__37444\ : std_logic;
signal \N__37439\ : std_logic;
signal \N__37438\ : std_logic;
signal \N__37437\ : std_logic;
signal \N__37434\ : std_logic;
signal \N__37429\ : std_logic;
signal \N__37424\ : std_logic;
signal \N__37423\ : std_logic;
signal \N__37422\ : std_logic;
signal \N__37419\ : std_logic;
signal \N__37414\ : std_logic;
signal \N__37409\ : std_logic;
signal \N__37406\ : std_logic;
signal \N__37405\ : std_logic;
signal \N__37402\ : std_logic;
signal \N__37399\ : std_logic;
signal \N__37398\ : std_logic;
signal \N__37395\ : std_logic;
signal \N__37390\ : std_logic;
signal \N__37385\ : std_logic;
signal \N__37382\ : std_logic;
signal \N__37379\ : std_logic;
signal \N__37378\ : std_logic;
signal \N__37375\ : std_logic;
signal \N__37372\ : std_logic;
signal \N__37369\ : std_logic;
signal \N__37364\ : std_logic;
signal \N__37363\ : std_logic;
signal \N__37362\ : std_logic;
signal \N__37361\ : std_logic;
signal \N__37354\ : std_logic;
signal \N__37351\ : std_logic;
signal \N__37350\ : std_logic;
signal \N__37349\ : std_logic;
signal \N__37346\ : std_logic;
signal \N__37343\ : std_logic;
signal \N__37338\ : std_logic;
signal \N__37333\ : std_logic;
signal \N__37328\ : std_logic;
signal \N__37327\ : std_logic;
signal \N__37326\ : std_logic;
signal \N__37323\ : std_logic;
signal \N__37320\ : std_logic;
signal \N__37317\ : std_logic;
signal \N__37314\ : std_logic;
signal \N__37313\ : std_logic;
signal \N__37310\ : std_logic;
signal \N__37307\ : std_logic;
signal \N__37304\ : std_logic;
signal \N__37301\ : std_logic;
signal \N__37296\ : std_logic;
signal \N__37293\ : std_logic;
signal \N__37290\ : std_logic;
signal \N__37287\ : std_logic;
signal \N__37280\ : std_logic;
signal \N__37279\ : std_logic;
signal \N__37278\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37276\ : std_logic;
signal \N__37275\ : std_logic;
signal \N__37264\ : std_logic;
signal \N__37261\ : std_logic;
signal \N__37260\ : std_logic;
signal \N__37257\ : std_logic;
signal \N__37256\ : std_logic;
signal \N__37255\ : std_logic;
signal \N__37254\ : std_logic;
signal \N__37251\ : std_logic;
signal \N__37248\ : std_logic;
signal \N__37245\ : std_logic;
signal \N__37238\ : std_logic;
signal \N__37235\ : std_logic;
signal \N__37226\ : std_logic;
signal \N__37225\ : std_logic;
signal \N__37224\ : std_logic;
signal \N__37221\ : std_logic;
signal \N__37218\ : std_logic;
signal \N__37215\ : std_logic;
signal \N__37212\ : std_logic;
signal \N__37209\ : std_logic;
signal \N__37206\ : std_logic;
signal \N__37203\ : std_logic;
signal \N__37202\ : std_logic;
signal \N__37197\ : std_logic;
signal \N__37194\ : std_logic;
signal \N__37191\ : std_logic;
signal \N__37188\ : std_logic;
signal \N__37181\ : std_logic;
signal \N__37178\ : std_logic;
signal \N__37175\ : std_logic;
signal \N__37174\ : std_logic;
signal \N__37171\ : std_logic;
signal \N__37168\ : std_logic;
signal \N__37165\ : std_logic;
signal \N__37160\ : std_logic;
signal \N__37157\ : std_logic;
signal \N__37154\ : std_logic;
signal \N__37151\ : std_logic;
signal \N__37150\ : std_logic;
signal \N__37147\ : std_logic;
signal \N__37144\ : std_logic;
signal \N__37141\ : std_logic;
signal \N__37136\ : std_logic;
signal \N__37133\ : std_logic;
signal \N__37130\ : std_logic;
signal \N__37127\ : std_logic;
signal \N__37126\ : std_logic;
signal \N__37123\ : std_logic;
signal \N__37120\ : std_logic;
signal \N__37117\ : std_logic;
signal \N__37112\ : std_logic;
signal \N__37109\ : std_logic;
signal \N__37106\ : std_logic;
signal \N__37103\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37099\ : std_logic;
signal \N__37096\ : std_logic;
signal \N__37093\ : std_logic;
signal \N__37090\ : std_logic;
signal \N__37085\ : std_logic;
signal \N__37082\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37076\ : std_logic;
signal \N__37075\ : std_logic;
signal \N__37072\ : std_logic;
signal \N__37069\ : std_logic;
signal \N__37066\ : std_logic;
signal \N__37063\ : std_logic;
signal \N__37062\ : std_logic;
signal \N__37059\ : std_logic;
signal \N__37056\ : std_logic;
signal \N__37053\ : std_logic;
signal \N__37046\ : std_logic;
signal \N__37043\ : std_logic;
signal \N__37040\ : std_logic;
signal \N__37037\ : std_logic;
signal \N__37034\ : std_logic;
signal \N__37031\ : std_logic;
signal \N__37028\ : std_logic;
signal \N__37025\ : std_logic;
signal \N__37022\ : std_logic;
signal \N__37019\ : std_logic;
signal \N__37016\ : std_logic;
signal \N__37013\ : std_logic;
signal \N__37010\ : std_logic;
signal \N__37007\ : std_logic;
signal \N__37004\ : std_logic;
signal \N__37001\ : std_logic;
signal \N__36998\ : std_logic;
signal \N__36995\ : std_logic;
signal \N__36992\ : std_logic;
signal \N__36989\ : std_logic;
signal \N__36986\ : std_logic;
signal \N__36983\ : std_logic;
signal \N__36980\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36974\ : std_logic;
signal \N__36971\ : std_logic;
signal \N__36968\ : std_logic;
signal \N__36965\ : std_logic;
signal \N__36962\ : std_logic;
signal \N__36961\ : std_logic;
signal \N__36958\ : std_logic;
signal \N__36955\ : std_logic;
signal \N__36952\ : std_logic;
signal \N__36947\ : std_logic;
signal \N__36944\ : std_logic;
signal \N__36941\ : std_logic;
signal \N__36938\ : std_logic;
signal \N__36935\ : std_logic;
signal \N__36934\ : std_logic;
signal \N__36931\ : std_logic;
signal \N__36928\ : std_logic;
signal \N__36925\ : std_logic;
signal \N__36920\ : std_logic;
signal \N__36917\ : std_logic;
signal \N__36914\ : std_logic;
signal \N__36911\ : std_logic;
signal \N__36908\ : std_logic;
signal \N__36905\ : std_logic;
signal \N__36902\ : std_logic;
signal \N__36899\ : std_logic;
signal \N__36896\ : std_logic;
signal \N__36895\ : std_logic;
signal \N__36892\ : std_logic;
signal \N__36889\ : std_logic;
signal \N__36886\ : std_logic;
signal \N__36881\ : std_logic;
signal \N__36878\ : std_logic;
signal \N__36875\ : std_logic;
signal \N__36872\ : std_logic;
signal \N__36869\ : std_logic;
signal \N__36866\ : std_logic;
signal \N__36863\ : std_logic;
signal \N__36860\ : std_logic;
signal \N__36857\ : std_logic;
signal \N__36854\ : std_logic;
signal \N__36851\ : std_logic;
signal \N__36848\ : std_logic;
signal \N__36845\ : std_logic;
signal \N__36842\ : std_logic;
signal \N__36839\ : std_logic;
signal \N__36836\ : std_logic;
signal \N__36833\ : std_logic;
signal \N__36830\ : std_logic;
signal \N__36827\ : std_logic;
signal \N__36826\ : std_logic;
signal \N__36823\ : std_logic;
signal \N__36820\ : std_logic;
signal \N__36817\ : std_logic;
signal \N__36814\ : std_logic;
signal \N__36809\ : std_logic;
signal \N__36806\ : std_logic;
signal \N__36803\ : std_logic;
signal \N__36800\ : std_logic;
signal \N__36797\ : std_logic;
signal \N__36794\ : std_logic;
signal \N__36791\ : std_logic;
signal \N__36788\ : std_logic;
signal \N__36785\ : std_logic;
signal \N__36782\ : std_logic;
signal \N__36779\ : std_logic;
signal \N__36776\ : std_logic;
signal \N__36773\ : std_logic;
signal \N__36770\ : std_logic;
signal \N__36767\ : std_logic;
signal \N__36764\ : std_logic;
signal \N__36761\ : std_logic;
signal \N__36758\ : std_logic;
signal \N__36755\ : std_logic;
signal \N__36752\ : std_logic;
signal \N__36749\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36743\ : std_logic;
signal \N__36742\ : std_logic;
signal \N__36739\ : std_logic;
signal \N__36736\ : std_logic;
signal \N__36731\ : std_logic;
signal \N__36728\ : std_logic;
signal \N__36725\ : std_logic;
signal \N__36722\ : std_logic;
signal \N__36719\ : std_logic;
signal \N__36718\ : std_logic;
signal \N__36715\ : std_logic;
signal \N__36712\ : std_logic;
signal \N__36707\ : std_logic;
signal \N__36704\ : std_logic;
signal \N__36701\ : std_logic;
signal \N__36700\ : std_logic;
signal \N__36697\ : std_logic;
signal \N__36694\ : std_logic;
signal \N__36693\ : std_logic;
signal \N__36688\ : std_logic;
signal \N__36685\ : std_logic;
signal \N__36682\ : std_logic;
signal \N__36677\ : std_logic;
signal \N__36674\ : std_logic;
signal \N__36673\ : std_logic;
signal \N__36670\ : std_logic;
signal \N__36669\ : std_logic;
signal \N__36666\ : std_logic;
signal \N__36663\ : std_logic;
signal \N__36660\ : std_logic;
signal \N__36655\ : std_logic;
signal \N__36650\ : std_logic;
signal \N__36647\ : std_logic;
signal \N__36646\ : std_logic;
signal \N__36643\ : std_logic;
signal \N__36642\ : std_logic;
signal \N__36639\ : std_logic;
signal \N__36636\ : std_logic;
signal \N__36633\ : std_logic;
signal \N__36628\ : std_logic;
signal \N__36623\ : std_logic;
signal \N__36620\ : std_logic;
signal \N__36619\ : std_logic;
signal \N__36616\ : std_logic;
signal \N__36613\ : std_logic;
signal \N__36612\ : std_logic;
signal \N__36607\ : std_logic;
signal \N__36604\ : std_logic;
signal \N__36601\ : std_logic;
signal \N__36596\ : std_logic;
signal \N__36593\ : std_logic;
signal \N__36592\ : std_logic;
signal \N__36589\ : std_logic;
signal \N__36586\ : std_logic;
signal \N__36585\ : std_logic;
signal \N__36580\ : std_logic;
signal \N__36577\ : std_logic;
signal \N__36574\ : std_logic;
signal \N__36569\ : std_logic;
signal \N__36566\ : std_logic;
signal \N__36565\ : std_logic;
signal \N__36562\ : std_logic;
signal \N__36559\ : std_logic;
signal \N__36556\ : std_logic;
signal \N__36551\ : std_logic;
signal \N__36548\ : std_logic;
signal \N__36547\ : std_logic;
signal \N__36546\ : std_logic;
signal \N__36545\ : std_logic;
signal \N__36544\ : std_logic;
signal \N__36543\ : std_logic;
signal \N__36542\ : std_logic;
signal \N__36541\ : std_logic;
signal \N__36540\ : std_logic;
signal \N__36539\ : std_logic;
signal \N__36538\ : std_logic;
signal \N__36537\ : std_logic;
signal \N__36536\ : std_logic;
signal \N__36535\ : std_logic;
signal \N__36534\ : std_logic;
signal \N__36533\ : std_logic;
signal \N__36532\ : std_logic;
signal \N__36531\ : std_logic;
signal \N__36530\ : std_logic;
signal \N__36529\ : std_logic;
signal \N__36528\ : std_logic;
signal \N__36527\ : std_logic;
signal \N__36526\ : std_logic;
signal \N__36525\ : std_logic;
signal \N__36524\ : std_logic;
signal \N__36523\ : std_logic;
signal \N__36522\ : std_logic;
signal \N__36521\ : std_logic;
signal \N__36520\ : std_logic;
signal \N__36519\ : std_logic;
signal \N__36510\ : std_logic;
signal \N__36501\ : std_logic;
signal \N__36492\ : std_logic;
signal \N__36483\ : std_logic;
signal \N__36478\ : std_logic;
signal \N__36469\ : std_logic;
signal \N__36460\ : std_logic;
signal \N__36451\ : std_logic;
signal \N__36448\ : std_logic;
signal \N__36433\ : std_logic;
signal \N__36428\ : std_logic;
signal \N__36425\ : std_logic;
signal \N__36424\ : std_logic;
signal \N__36421\ : std_logic;
signal \N__36418\ : std_logic;
signal \N__36415\ : std_logic;
signal \N__36410\ : std_logic;
signal \N__36409\ : std_logic;
signal \N__36408\ : std_logic;
signal \N__36407\ : std_logic;
signal \N__36404\ : std_logic;
signal \N__36401\ : std_logic;
signal \N__36398\ : std_logic;
signal \N__36395\ : std_logic;
signal \N__36390\ : std_logic;
signal \N__36385\ : std_logic;
signal \N__36382\ : std_logic;
signal \N__36377\ : std_logic;
signal \N__36374\ : std_logic;
signal \N__36371\ : std_logic;
signal \N__36368\ : std_logic;
signal \N__36365\ : std_logic;
signal \N__36364\ : std_logic;
signal \N__36361\ : std_logic;
signal \N__36358\ : std_logic;
signal \N__36357\ : std_logic;
signal \N__36352\ : std_logic;
signal \N__36349\ : std_logic;
signal \N__36346\ : std_logic;
signal \N__36341\ : std_logic;
signal \N__36338\ : std_logic;
signal \N__36337\ : std_logic;
signal \N__36334\ : std_logic;
signal \N__36331\ : std_logic;
signal \N__36330\ : std_logic;
signal \N__36325\ : std_logic;
signal \N__36322\ : std_logic;
signal \N__36319\ : std_logic;
signal \N__36314\ : std_logic;
signal \N__36311\ : std_logic;
signal \N__36310\ : std_logic;
signal \N__36307\ : std_logic;
signal \N__36304\ : std_logic;
signal \N__36303\ : std_logic;
signal \N__36300\ : std_logic;
signal \N__36297\ : std_logic;
signal \N__36294\ : std_logic;
signal \N__36289\ : std_logic;
signal \N__36284\ : std_logic;
signal \N__36281\ : std_logic;
signal \N__36280\ : std_logic;
signal \N__36277\ : std_logic;
signal \N__36276\ : std_logic;
signal \N__36273\ : std_logic;
signal \N__36270\ : std_logic;
signal \N__36267\ : std_logic;
signal \N__36262\ : std_logic;
signal \N__36257\ : std_logic;
signal \N__36254\ : std_logic;
signal \N__36253\ : std_logic;
signal \N__36250\ : std_logic;
signal \N__36247\ : std_logic;
signal \N__36246\ : std_logic;
signal \N__36241\ : std_logic;
signal \N__36238\ : std_logic;
signal \N__36235\ : std_logic;
signal \N__36230\ : std_logic;
signal \N__36227\ : std_logic;
signal \N__36226\ : std_logic;
signal \N__36223\ : std_logic;
signal \N__36220\ : std_logic;
signal \N__36219\ : std_logic;
signal \N__36214\ : std_logic;
signal \N__36211\ : std_logic;
signal \N__36208\ : std_logic;
signal \N__36203\ : std_logic;
signal \N__36200\ : std_logic;
signal \N__36199\ : std_logic;
signal \N__36198\ : std_logic;
signal \N__36193\ : std_logic;
signal \N__36190\ : std_logic;
signal \N__36187\ : std_logic;
signal \N__36182\ : std_logic;
signal \N__36179\ : std_logic;
signal \N__36178\ : std_logic;
signal \N__36177\ : std_logic;
signal \N__36172\ : std_logic;
signal \N__36169\ : std_logic;
signal \N__36166\ : std_logic;
signal \N__36161\ : std_logic;
signal \N__36158\ : std_logic;
signal \N__36157\ : std_logic;
signal \N__36154\ : std_logic;
signal \N__36151\ : std_logic;
signal \N__36150\ : std_logic;
signal \N__36145\ : std_logic;
signal \N__36142\ : std_logic;
signal \N__36139\ : std_logic;
signal \N__36134\ : std_logic;
signal \N__36131\ : std_logic;
signal \N__36130\ : std_logic;
signal \N__36129\ : std_logic;
signal \N__36124\ : std_logic;
signal \N__36121\ : std_logic;
signal \N__36118\ : std_logic;
signal \N__36113\ : std_logic;
signal \N__36110\ : std_logic;
signal \N__36109\ : std_logic;
signal \N__36108\ : std_logic;
signal \N__36103\ : std_logic;
signal \N__36100\ : std_logic;
signal \N__36097\ : std_logic;
signal \N__36092\ : std_logic;
signal \N__36089\ : std_logic;
signal \N__36086\ : std_logic;
signal \N__36083\ : std_logic;
signal \N__36082\ : std_logic;
signal \N__36079\ : std_logic;
signal \N__36078\ : std_logic;
signal \N__36075\ : std_logic;
signal \N__36072\ : std_logic;
signal \N__36069\ : std_logic;
signal \N__36064\ : std_logic;
signal \N__36059\ : std_logic;
signal \N__36056\ : std_logic;
signal \N__36055\ : std_logic;
signal \N__36052\ : std_logic;
signal \N__36049\ : std_logic;
signal \N__36046\ : std_logic;
signal \N__36045\ : std_logic;
signal \N__36040\ : std_logic;
signal \N__36037\ : std_logic;
signal \N__36034\ : std_logic;
signal \N__36029\ : std_logic;
signal \N__36026\ : std_logic;
signal \N__36025\ : std_logic;
signal \N__36022\ : std_logic;
signal \N__36019\ : std_logic;
signal \N__36018\ : std_logic;
signal \N__36013\ : std_logic;
signal \N__36010\ : std_logic;
signal \N__36007\ : std_logic;
signal \N__36002\ : std_logic;
signal \N__35999\ : std_logic;
signal \N__35998\ : std_logic;
signal \N__35995\ : std_logic;
signal \N__35992\ : std_logic;
signal \N__35991\ : std_logic;
signal \N__35986\ : std_logic;
signal \N__35983\ : std_logic;
signal \N__35980\ : std_logic;
signal \N__35975\ : std_logic;
signal \N__35972\ : std_logic;
signal \N__35971\ : std_logic;
signal \N__35970\ : std_logic;
signal \N__35965\ : std_logic;
signal \N__35962\ : std_logic;
signal \N__35959\ : std_logic;
signal \N__35954\ : std_logic;
signal \N__35951\ : std_logic;
signal \N__35950\ : std_logic;
signal \N__35949\ : std_logic;
signal \N__35944\ : std_logic;
signal \N__35941\ : std_logic;
signal \N__35938\ : std_logic;
signal \N__35933\ : std_logic;
signal \N__35930\ : std_logic;
signal \N__35929\ : std_logic;
signal \N__35926\ : std_logic;
signal \N__35923\ : std_logic;
signal \N__35920\ : std_logic;
signal \N__35917\ : std_logic;
signal \N__35916\ : std_logic;
signal \N__35911\ : std_logic;
signal \N__35908\ : std_logic;
signal \N__35903\ : std_logic;
signal \N__35900\ : std_logic;
signal \N__35899\ : std_logic;
signal \N__35896\ : std_logic;
signal \N__35893\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35885\ : std_logic;
signal \N__35882\ : std_logic;
signal \N__35881\ : std_logic;
signal \N__35878\ : std_logic;
signal \N__35875\ : std_logic;
signal \N__35872\ : std_logic;
signal \N__35869\ : std_logic;
signal \N__35868\ : std_logic;
signal \N__35863\ : std_logic;
signal \N__35860\ : std_logic;
signal \N__35855\ : std_logic;
signal \N__35854\ : std_logic;
signal \N__35851\ : std_logic;
signal \N__35850\ : std_logic;
signal \N__35847\ : std_logic;
signal \N__35844\ : std_logic;
signal \N__35841\ : std_logic;
signal \N__35836\ : std_logic;
signal \N__35831\ : std_logic;
signal \N__35828\ : std_logic;
signal \N__35827\ : std_logic;
signal \N__35824\ : std_logic;
signal \N__35821\ : std_logic;
signal \N__35820\ : std_logic;
signal \N__35817\ : std_logic;
signal \N__35814\ : std_logic;
signal \N__35811\ : std_logic;
signal \N__35808\ : std_logic;
signal \N__35801\ : std_logic;
signal \N__35798\ : std_logic;
signal \N__35797\ : std_logic;
signal \N__35796\ : std_logic;
signal \N__35791\ : std_logic;
signal \N__35788\ : std_logic;
signal \N__35785\ : std_logic;
signal \N__35780\ : std_logic;
signal \N__35777\ : std_logic;
signal \N__35776\ : std_logic;
signal \N__35775\ : std_logic;
signal \N__35770\ : std_logic;
signal \N__35767\ : std_logic;
signal \N__35764\ : std_logic;
signal \N__35759\ : std_logic;
signal \N__35756\ : std_logic;
signal \N__35755\ : std_logic;
signal \N__35752\ : std_logic;
signal \N__35749\ : std_logic;
signal \N__35744\ : std_logic;
signal \N__35743\ : std_logic;
signal \N__35740\ : std_logic;
signal \N__35737\ : std_logic;
signal \N__35734\ : std_logic;
signal \N__35729\ : std_logic;
signal \N__35726\ : std_logic;
signal \N__35725\ : std_logic;
signal \N__35722\ : std_logic;
signal \N__35719\ : std_logic;
signal \N__35718\ : std_logic;
signal \N__35713\ : std_logic;
signal \N__35710\ : std_logic;
signal \N__35707\ : std_logic;
signal \N__35702\ : std_logic;
signal \N__35699\ : std_logic;
signal \N__35698\ : std_logic;
signal \N__35697\ : std_logic;
signal \N__35696\ : std_logic;
signal \N__35695\ : std_logic;
signal \N__35684\ : std_logic;
signal \N__35681\ : std_logic;
signal \N__35678\ : std_logic;
signal \N__35677\ : std_logic;
signal \N__35674\ : std_logic;
signal \N__35671\ : std_logic;
signal \N__35670\ : std_logic;
signal \N__35667\ : std_logic;
signal \N__35664\ : std_logic;
signal \N__35661\ : std_logic;
signal \N__35658\ : std_logic;
signal \N__35657\ : std_logic;
signal \N__35656\ : std_logic;
signal \N__35651\ : std_logic;
signal \N__35648\ : std_logic;
signal \N__35645\ : std_logic;
signal \N__35642\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35630\ : std_logic;
signal \N__35627\ : std_logic;
signal \N__35624\ : std_logic;
signal \N__35621\ : std_logic;
signal \N__35618\ : std_logic;
signal \N__35615\ : std_logic;
signal \N__35612\ : std_logic;
signal \N__35609\ : std_logic;
signal \N__35606\ : std_logic;
signal \N__35603\ : std_logic;
signal \N__35600\ : std_logic;
signal \N__35597\ : std_logic;
signal \N__35594\ : std_logic;
signal \N__35593\ : std_logic;
signal \N__35592\ : std_logic;
signal \N__35589\ : std_logic;
signal \N__35584\ : std_logic;
signal \N__35579\ : std_logic;
signal \N__35576\ : std_logic;
signal \N__35573\ : std_logic;
signal \N__35570\ : std_logic;
signal \N__35569\ : std_logic;
signal \N__35566\ : std_logic;
signal \N__35563\ : std_logic;
signal \N__35560\ : std_logic;
signal \N__35559\ : std_logic;
signal \N__35558\ : std_logic;
signal \N__35553\ : std_logic;
signal \N__35548\ : std_logic;
signal \N__35543\ : std_logic;
signal \N__35540\ : std_logic;
signal \N__35539\ : std_logic;
signal \N__35538\ : std_logic;
signal \N__35535\ : std_logic;
signal \N__35532\ : std_logic;
signal \N__35529\ : std_logic;
signal \N__35522\ : std_logic;
signal \N__35519\ : std_logic;
signal \N__35518\ : std_logic;
signal \N__35517\ : std_logic;
signal \N__35514\ : std_logic;
signal \N__35513\ : std_logic;
signal \N__35510\ : std_logic;
signal \N__35507\ : std_logic;
signal \N__35504\ : std_logic;
signal \N__35501\ : std_logic;
signal \N__35500\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35494\ : std_logic;
signal \N__35491\ : std_logic;
signal \N__35488\ : std_logic;
signal \N__35485\ : std_logic;
signal \N__35482\ : std_logic;
signal \N__35479\ : std_logic;
signal \N__35474\ : std_logic;
signal \N__35471\ : std_logic;
signal \N__35468\ : std_logic;
signal \N__35465\ : std_logic;
signal \N__35462\ : std_logic;
signal \N__35453\ : std_logic;
signal \N__35450\ : std_logic;
signal \N__35449\ : std_logic;
signal \N__35448\ : std_logic;
signal \N__35445\ : std_logic;
signal \N__35442\ : std_logic;
signal \N__35439\ : std_logic;
signal \N__35432\ : std_logic;
signal \N__35431\ : std_logic;
signal \N__35428\ : std_logic;
signal \N__35427\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35422\ : std_logic;
signal \N__35419\ : std_logic;
signal \N__35416\ : std_logic;
signal \N__35413\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35407\ : std_logic;
signal \N__35404\ : std_logic;
signal \N__35401\ : std_logic;
signal \N__35398\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35389\ : std_logic;
signal \N__35386\ : std_logic;
signal \N__35383\ : std_logic;
signal \N__35380\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35363\ : std_logic;
signal \N__35360\ : std_logic;
signal \N__35357\ : std_logic;
signal \N__35354\ : std_logic;
signal \N__35351\ : std_logic;
signal \N__35348\ : std_logic;
signal \N__35345\ : std_logic;
signal \N__35342\ : std_logic;
signal \N__35339\ : std_logic;
signal \N__35336\ : std_logic;
signal \N__35333\ : std_logic;
signal \N__35330\ : std_logic;
signal \N__35327\ : std_logic;
signal \N__35324\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35318\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35314\ : std_logic;
signal \N__35313\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35302\ : std_logic;
signal \N__35299\ : std_logic;
signal \N__35298\ : std_logic;
signal \N__35295\ : std_logic;
signal \N__35292\ : std_logic;
signal \N__35289\ : std_logic;
signal \N__35288\ : std_logic;
signal \N__35285\ : std_logic;
signal \N__35280\ : std_logic;
signal \N__35277\ : std_logic;
signal \N__35270\ : std_logic;
signal \N__35267\ : std_logic;
signal \N__35264\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35260\ : std_logic;
signal \N__35259\ : std_logic;
signal \N__35258\ : std_logic;
signal \N__35257\ : std_logic;
signal \N__35256\ : std_logic;
signal \N__35253\ : std_logic;
signal \N__35250\ : std_logic;
signal \N__35249\ : std_logic;
signal \N__35246\ : std_logic;
signal \N__35243\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35232\ : std_logic;
signal \N__35229\ : std_logic;
signal \N__35224\ : std_logic;
signal \N__35213\ : std_logic;
signal \N__35210\ : std_logic;
signal \N__35207\ : std_logic;
signal \N__35206\ : std_logic;
signal \N__35203\ : std_logic;
signal \N__35200\ : std_logic;
signal \N__35195\ : std_logic;
signal \N__35194\ : std_logic;
signal \N__35191\ : std_logic;
signal \N__35188\ : std_logic;
signal \N__35183\ : std_logic;
signal \N__35180\ : std_logic;
signal \N__35177\ : std_logic;
signal \N__35174\ : std_logic;
signal \N__35171\ : std_logic;
signal \N__35170\ : std_logic;
signal \N__35167\ : std_logic;
signal \N__35162\ : std_logic;
signal \N__35159\ : std_logic;
signal \N__35156\ : std_logic;
signal \N__35155\ : std_logic;
signal \N__35150\ : std_logic;
signal \N__35147\ : std_logic;
signal \N__35144\ : std_logic;
signal \N__35143\ : std_logic;
signal \N__35140\ : std_logic;
signal \N__35137\ : std_logic;
signal \N__35132\ : std_logic;
signal \N__35129\ : std_logic;
signal \N__35128\ : std_logic;
signal \N__35125\ : std_logic;
signal \N__35124\ : std_logic;
signal \N__35121\ : std_logic;
signal \N__35118\ : std_logic;
signal \N__35117\ : std_logic;
signal \N__35114\ : std_logic;
signal \N__35111\ : std_logic;
signal \N__35108\ : std_logic;
signal \N__35105\ : std_logic;
signal \N__35102\ : std_logic;
signal \N__35099\ : std_logic;
signal \N__35090\ : std_logic;
signal \N__35087\ : std_logic;
signal \N__35084\ : std_logic;
signal \N__35081\ : std_logic;
signal \N__35080\ : std_logic;
signal \N__35077\ : std_logic;
signal \N__35076\ : std_logic;
signal \N__35075\ : std_logic;
signal \N__35072\ : std_logic;
signal \N__35069\ : std_logic;
signal \N__35066\ : std_logic;
signal \N__35063\ : std_logic;
signal \N__35060\ : std_logic;
signal \N__35057\ : std_logic;
signal \N__35054\ : std_logic;
signal \N__35049\ : std_logic;
signal \N__35042\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35035\ : std_logic;
signal \N__35032\ : std_logic;
signal \N__35031\ : std_logic;
signal \N__35028\ : std_logic;
signal \N__35025\ : std_logic;
signal \N__35022\ : std_logic;
signal \N__35015\ : std_logic;
signal \N__35012\ : std_logic;
signal \N__35011\ : std_logic;
signal \N__35008\ : std_logic;
signal \N__35003\ : std_logic;
signal \N__35002\ : std_logic;
signal \N__34999\ : std_logic;
signal \N__34996\ : std_logic;
signal \N__34991\ : std_logic;
signal \N__34988\ : std_logic;
signal \N__34985\ : std_logic;
signal \N__34984\ : std_logic;
signal \N__34983\ : std_logic;
signal \N__34978\ : std_logic;
signal \N__34975\ : std_logic;
signal \N__34972\ : std_logic;
signal \N__34969\ : std_logic;
signal \N__34964\ : std_logic;
signal \N__34961\ : std_logic;
signal \N__34960\ : std_logic;
signal \N__34957\ : std_logic;
signal \N__34954\ : std_logic;
signal \N__34951\ : std_logic;
signal \N__34948\ : std_logic;
signal \N__34947\ : std_logic;
signal \N__34944\ : std_logic;
signal \N__34941\ : std_logic;
signal \N__34938\ : std_logic;
signal \N__34935\ : std_logic;
signal \N__34928\ : std_logic;
signal \N__34925\ : std_logic;
signal \N__34922\ : std_logic;
signal \N__34919\ : std_logic;
signal \N__34916\ : std_logic;
signal \N__34913\ : std_logic;
signal \N__34910\ : std_logic;
signal \N__34907\ : std_logic;
signal \N__34906\ : std_logic;
signal \N__34905\ : std_logic;
signal \N__34904\ : std_logic;
signal \N__34901\ : std_logic;
signal \N__34894\ : std_logic;
signal \N__34891\ : std_logic;
signal \N__34888\ : std_logic;
signal \N__34885\ : std_logic;
signal \N__34882\ : std_logic;
signal \N__34879\ : std_logic;
signal \N__34876\ : std_logic;
signal \N__34871\ : std_logic;
signal \N__34868\ : std_logic;
signal \N__34865\ : std_logic;
signal \N__34862\ : std_logic;
signal \N__34859\ : std_logic;
signal \N__34858\ : std_logic;
signal \N__34855\ : std_logic;
signal \N__34852\ : std_logic;
signal \N__34847\ : std_logic;
signal \N__34844\ : std_logic;
signal \N__34841\ : std_logic;
signal \N__34840\ : std_logic;
signal \N__34839\ : std_logic;
signal \N__34836\ : std_logic;
signal \N__34833\ : std_logic;
signal \N__34830\ : std_logic;
signal \N__34823\ : std_logic;
signal \N__34820\ : std_logic;
signal \N__34817\ : std_logic;
signal \N__34814\ : std_logic;
signal \N__34813\ : std_logic;
signal \N__34810\ : std_logic;
signal \N__34807\ : std_logic;
signal \N__34804\ : std_logic;
signal \N__34803\ : std_logic;
signal \N__34800\ : std_logic;
signal \N__34797\ : std_logic;
signal \N__34794\ : std_logic;
signal \N__34791\ : std_logic;
signal \N__34784\ : std_logic;
signal \N__34781\ : std_logic;
signal \N__34778\ : std_logic;
signal \N__34775\ : std_logic;
signal \N__34772\ : std_logic;
signal \N__34769\ : std_logic;
signal \N__34766\ : std_logic;
signal \N__34763\ : std_logic;
signal \N__34760\ : std_logic;
signal \N__34757\ : std_logic;
signal \N__34754\ : std_logic;
signal \N__34751\ : std_logic;
signal \N__34748\ : std_logic;
signal \N__34745\ : std_logic;
signal \N__34742\ : std_logic;
signal \N__34739\ : std_logic;
signal \N__34736\ : std_logic;
signal \N__34733\ : std_logic;
signal \N__34730\ : std_logic;
signal \N__34727\ : std_logic;
signal \N__34726\ : std_logic;
signal \N__34723\ : std_logic;
signal \N__34720\ : std_logic;
signal \N__34715\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34709\ : std_logic;
signal \N__34706\ : std_logic;
signal \N__34703\ : std_logic;
signal \N__34700\ : std_logic;
signal \N__34699\ : std_logic;
signal \N__34696\ : std_logic;
signal \N__34693\ : std_logic;
signal \N__34688\ : std_logic;
signal \N__34685\ : std_logic;
signal \N__34682\ : std_logic;
signal \N__34679\ : std_logic;
signal \N__34676\ : std_logic;
signal \N__34673\ : std_logic;
signal \N__34670\ : std_logic;
signal \N__34667\ : std_logic;
signal \N__34666\ : std_logic;
signal \N__34663\ : std_logic;
signal \N__34660\ : std_logic;
signal \N__34655\ : std_logic;
signal \N__34652\ : std_logic;
signal \N__34649\ : std_logic;
signal \N__34646\ : std_logic;
signal \N__34643\ : std_logic;
signal \N__34640\ : std_logic;
signal \N__34637\ : std_logic;
signal \N__34636\ : std_logic;
signal \N__34633\ : std_logic;
signal \N__34630\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34624\ : std_logic;
signal \N__34619\ : std_logic;
signal \N__34616\ : std_logic;
signal \N__34613\ : std_logic;
signal \N__34610\ : std_logic;
signal \N__34607\ : std_logic;
signal \N__34606\ : std_logic;
signal \N__34603\ : std_logic;
signal \N__34600\ : std_logic;
signal \N__34597\ : std_logic;
signal \N__34592\ : std_logic;
signal \N__34589\ : std_logic;
signal \N__34586\ : std_logic;
signal \N__34583\ : std_logic;
signal \N__34580\ : std_logic;
signal \N__34577\ : std_logic;
signal \N__34574\ : std_logic;
signal \N__34571\ : std_logic;
signal \N__34568\ : std_logic;
signal \N__34565\ : std_logic;
signal \N__34564\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34557\ : std_logic;
signal \N__34552\ : std_logic;
signal \N__34549\ : std_logic;
signal \N__34546\ : std_logic;
signal \N__34545\ : std_logic;
signal \N__34544\ : std_logic;
signal \N__34541\ : std_logic;
signal \N__34538\ : std_logic;
signal \N__34537\ : std_logic;
signal \N__34536\ : std_logic;
signal \N__34531\ : std_logic;
signal \N__34528\ : std_logic;
signal \N__34525\ : std_logic;
signal \N__34522\ : std_logic;
signal \N__34519\ : std_logic;
signal \N__34516\ : std_logic;
signal \N__34513\ : std_logic;
signal \N__34510\ : std_logic;
signal \N__34507\ : std_logic;
signal \N__34504\ : std_logic;
signal \N__34501\ : std_logic;
signal \N__34498\ : std_logic;
signal \N__34491\ : std_logic;
signal \N__34488\ : std_logic;
signal \N__34483\ : std_logic;
signal \N__34480\ : std_logic;
signal \N__34475\ : std_logic;
signal \N__34474\ : std_logic;
signal \N__34471\ : std_logic;
signal \N__34468\ : std_logic;
signal \N__34465\ : std_logic;
signal \N__34462\ : std_logic;
signal \N__34459\ : std_logic;
signal \N__34454\ : std_logic;
signal \N__34453\ : std_logic;
signal \N__34448\ : std_logic;
signal \N__34445\ : std_logic;
signal \N__34442\ : std_logic;
signal \N__34439\ : std_logic;
signal \N__34436\ : std_logic;
signal \N__34433\ : std_logic;
signal \N__34432\ : std_logic;
signal \N__34431\ : std_logic;
signal \N__34428\ : std_logic;
signal \N__34423\ : std_logic;
signal \N__34418\ : std_logic;
signal \N__34417\ : std_logic;
signal \N__34412\ : std_logic;
signal \N__34411\ : std_logic;
signal \N__34410\ : std_logic;
signal \N__34407\ : std_logic;
signal \N__34404\ : std_logic;
signal \N__34403\ : std_logic;
signal \N__34402\ : std_logic;
signal \N__34399\ : std_logic;
signal \N__34396\ : std_logic;
signal \N__34393\ : std_logic;
signal \N__34388\ : std_logic;
signal \N__34379\ : std_logic;
signal \N__34376\ : std_logic;
signal \N__34373\ : std_logic;
signal \N__34370\ : std_logic;
signal \N__34369\ : std_logic;
signal \N__34366\ : std_logic;
signal \N__34365\ : std_logic;
signal \N__34362\ : std_logic;
signal \N__34359\ : std_logic;
signal \N__34356\ : std_logic;
signal \N__34349\ : std_logic;
signal \N__34346\ : std_logic;
signal \N__34345\ : std_logic;
signal \N__34342\ : std_logic;
signal \N__34339\ : std_logic;
signal \N__34334\ : std_logic;
signal \N__34331\ : std_logic;
signal \N__34328\ : std_logic;
signal \N__34325\ : std_logic;
signal \N__34322\ : std_logic;
signal \N__34319\ : std_logic;
signal \N__34316\ : std_logic;
signal \N__34313\ : std_logic;
signal \N__34310\ : std_logic;
signal \N__34309\ : std_logic;
signal \N__34306\ : std_logic;
signal \N__34303\ : std_logic;
signal \N__34298\ : std_logic;
signal \N__34295\ : std_logic;
signal \N__34292\ : std_logic;
signal \N__34289\ : std_logic;
signal \N__34286\ : std_logic;
signal \N__34283\ : std_logic;
signal \N__34280\ : std_logic;
signal \N__34279\ : std_logic;
signal \N__34276\ : std_logic;
signal \N__34273\ : std_logic;
signal \N__34268\ : std_logic;
signal \N__34265\ : std_logic;
signal \N__34262\ : std_logic;
signal \N__34259\ : std_logic;
signal \N__34256\ : std_logic;
signal \N__34253\ : std_logic;
signal \N__34250\ : std_logic;
signal \N__34249\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34243\ : std_logic;
signal \N__34238\ : std_logic;
signal \N__34235\ : std_logic;
signal \N__34232\ : std_logic;
signal \N__34229\ : std_logic;
signal \N__34226\ : std_logic;
signal \N__34223\ : std_logic;
signal \N__34220\ : std_logic;
signal \N__34217\ : std_logic;
signal \N__34214\ : std_logic;
signal \N__34211\ : std_logic;
signal \N__34208\ : std_logic;
signal \N__34205\ : std_logic;
signal \N__34202\ : std_logic;
signal \N__34199\ : std_logic;
signal \N__34196\ : std_logic;
signal \N__34193\ : std_logic;
signal \N__34190\ : std_logic;
signal \N__34187\ : std_logic;
signal \N__34184\ : std_logic;
signal \N__34181\ : std_logic;
signal \N__34178\ : std_logic;
signal \N__34175\ : std_logic;
signal \N__34172\ : std_logic;
signal \N__34169\ : std_logic;
signal \N__34166\ : std_logic;
signal \N__34165\ : std_logic;
signal \N__34162\ : std_logic;
signal \N__34159\ : std_logic;
signal \N__34158\ : std_logic;
signal \N__34155\ : std_logic;
signal \N__34152\ : std_logic;
signal \N__34151\ : std_logic;
signal \N__34150\ : std_logic;
signal \N__34147\ : std_logic;
signal \N__34144\ : std_logic;
signal \N__34141\ : std_logic;
signal \N__34138\ : std_logic;
signal \N__34135\ : std_logic;
signal \N__34132\ : std_logic;
signal \N__34125\ : std_logic;
signal \N__34122\ : std_logic;
signal \N__34115\ : std_logic;
signal \N__34114\ : std_logic;
signal \N__34111\ : std_logic;
signal \N__34108\ : std_logic;
signal \N__34107\ : std_logic;
signal \N__34106\ : std_logic;
signal \N__34103\ : std_logic;
signal \N__34100\ : std_logic;
signal \N__34099\ : std_logic;
signal \N__34096\ : std_logic;
signal \N__34093\ : std_logic;
signal \N__34090\ : std_logic;
signal \N__34087\ : std_logic;
signal \N__34084\ : std_logic;
signal \N__34081\ : std_logic;
signal \N__34078\ : std_logic;
signal \N__34075\ : std_logic;
signal \N__34072\ : std_logic;
signal \N__34069\ : std_logic;
signal \N__34066\ : std_logic;
signal \N__34055\ : std_logic;
signal \N__34052\ : std_logic;
signal \N__34049\ : std_logic;
signal \N__34048\ : std_logic;
signal \N__34047\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34043\ : std_logic;
signal \N__34040\ : std_logic;
signal \N__34037\ : std_logic;
signal \N__34034\ : std_logic;
signal \N__34031\ : std_logic;
signal \N__34030\ : std_logic;
signal \N__34029\ : std_logic;
signal \N__34024\ : std_logic;
signal \N__34021\ : std_logic;
signal \N__34018\ : std_logic;
signal \N__34015\ : std_logic;
signal \N__34012\ : std_logic;
signal \N__34009\ : std_logic;
signal \N__33998\ : std_logic;
signal \N__33995\ : std_logic;
signal \N__33992\ : std_logic;
signal \N__33989\ : std_logic;
signal \N__33986\ : std_logic;
signal \N__33983\ : std_logic;
signal \N__33980\ : std_logic;
signal \N__33977\ : std_logic;
signal \N__33974\ : std_logic;
signal \N__33971\ : std_logic;
signal \N__33968\ : std_logic;
signal \N__33965\ : std_logic;
signal \N__33962\ : std_logic;
signal \N__33959\ : std_logic;
signal \N__33956\ : std_logic;
signal \N__33953\ : std_logic;
signal \N__33950\ : std_logic;
signal \N__33947\ : std_logic;
signal \N__33944\ : std_logic;
signal \N__33941\ : std_logic;
signal \N__33938\ : std_logic;
signal \N__33935\ : std_logic;
signal \N__33932\ : std_logic;
signal \N__33929\ : std_logic;
signal \N__33926\ : std_logic;
signal \N__33923\ : std_logic;
signal \N__33920\ : std_logic;
signal \N__33917\ : std_logic;
signal \N__33916\ : std_logic;
signal \N__33913\ : std_logic;
signal \N__33910\ : std_logic;
signal \N__33907\ : std_logic;
signal \N__33904\ : std_logic;
signal \N__33903\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33901\ : std_logic;
signal \N__33898\ : std_logic;
signal \N__33895\ : std_logic;
signal \N__33892\ : std_logic;
signal \N__33887\ : std_logic;
signal \N__33878\ : std_logic;
signal \N__33877\ : std_logic;
signal \N__33876\ : std_logic;
signal \N__33873\ : std_logic;
signal \N__33870\ : std_logic;
signal \N__33867\ : std_logic;
signal \N__33866\ : std_logic;
signal \N__33863\ : std_logic;
signal \N__33860\ : std_logic;
signal \N__33857\ : std_logic;
signal \N__33854\ : std_logic;
signal \N__33853\ : std_logic;
signal \N__33850\ : std_logic;
signal \N__33845\ : std_logic;
signal \N__33840\ : std_logic;
signal \N__33833\ : std_logic;
signal \N__33832\ : std_logic;
signal \N__33827\ : std_logic;
signal \N__33826\ : std_logic;
signal \N__33823\ : std_logic;
signal \N__33820\ : std_logic;
signal \N__33817\ : std_logic;
signal \N__33812\ : std_logic;
signal \N__33809\ : std_logic;
signal \N__33806\ : std_logic;
signal \N__33805\ : std_logic;
signal \N__33804\ : std_logic;
signal \N__33801\ : std_logic;
signal \N__33796\ : std_logic;
signal \N__33791\ : std_logic;
signal \N__33788\ : std_logic;
signal \N__33787\ : std_logic;
signal \N__33784\ : std_logic;
signal \N__33783\ : std_logic;
signal \N__33780\ : std_logic;
signal \N__33777\ : std_logic;
signal \N__33774\ : std_logic;
signal \N__33773\ : std_logic;
signal \N__33770\ : std_logic;
signal \N__33767\ : std_logic;
signal \N__33762\ : std_logic;
signal \N__33755\ : std_logic;
signal \N__33752\ : std_logic;
signal \N__33749\ : std_logic;
signal \N__33746\ : std_logic;
signal \N__33743\ : std_logic;
signal \N__33740\ : std_logic;
signal \N__33737\ : std_logic;
signal \N__33734\ : std_logic;
signal \N__33731\ : std_logic;
signal \N__33728\ : std_logic;
signal \N__33725\ : std_logic;
signal \N__33722\ : std_logic;
signal \N__33719\ : std_logic;
signal \N__33716\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33712\ : std_logic;
signal \N__33711\ : std_logic;
signal \N__33704\ : std_logic;
signal \N__33701\ : std_logic;
signal \N__33698\ : std_logic;
signal \N__33695\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33691\ : std_logic;
signal \N__33688\ : std_logic;
signal \N__33685\ : std_logic;
signal \N__33680\ : std_logic;
signal \N__33677\ : std_logic;
signal \N__33674\ : std_logic;
signal \N__33671\ : std_logic;
signal \N__33668\ : std_logic;
signal \N__33665\ : std_logic;
signal \N__33662\ : std_logic;
signal \N__33659\ : std_logic;
signal \N__33656\ : std_logic;
signal \N__33653\ : std_logic;
signal \N__33650\ : std_logic;
signal \N__33647\ : std_logic;
signal \N__33646\ : std_logic;
signal \N__33641\ : std_logic;
signal \N__33638\ : std_logic;
signal \N__33635\ : std_logic;
signal \N__33632\ : std_logic;
signal \N__33629\ : std_logic;
signal \N__33628\ : std_logic;
signal \N__33623\ : std_logic;
signal \N__33620\ : std_logic;
signal \N__33617\ : std_logic;
signal \N__33614\ : std_logic;
signal \N__33611\ : std_logic;
signal \N__33608\ : std_logic;
signal \N__33605\ : std_logic;
signal \N__33602\ : std_logic;
signal \N__33599\ : std_logic;
signal \N__33596\ : std_logic;
signal \N__33593\ : std_logic;
signal \N__33592\ : std_logic;
signal \N__33591\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33585\ : std_logic;
signal \N__33582\ : std_logic;
signal \N__33579\ : std_logic;
signal \N__33576\ : std_logic;
signal \N__33569\ : std_logic;
signal \N__33566\ : std_logic;
signal \N__33563\ : std_logic;
signal \N__33560\ : std_logic;
signal \N__33557\ : std_logic;
signal \N__33554\ : std_logic;
signal \N__33553\ : std_logic;
signal \N__33550\ : std_logic;
signal \N__33547\ : std_logic;
signal \N__33542\ : std_logic;
signal \N__33541\ : std_logic;
signal \N__33538\ : std_logic;
signal \N__33535\ : std_logic;
signal \N__33530\ : std_logic;
signal \N__33529\ : std_logic;
signal \N__33526\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33520\ : std_logic;
signal \N__33515\ : std_logic;
signal \N__33514\ : std_logic;
signal \N__33513\ : std_logic;
signal \N__33512\ : std_logic;
signal \N__33509\ : std_logic;
signal \N__33506\ : std_logic;
signal \N__33503\ : std_logic;
signal \N__33500\ : std_logic;
signal \N__33491\ : std_logic;
signal \N__33490\ : std_logic;
signal \N__33489\ : std_logic;
signal \N__33486\ : std_logic;
signal \N__33483\ : std_logic;
signal \N__33482\ : std_logic;
signal \N__33479\ : std_logic;
signal \N__33476\ : std_logic;
signal \N__33473\ : std_logic;
signal \N__33470\ : std_logic;
signal \N__33463\ : std_logic;
signal \N__33460\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33452\ : std_logic;
signal \N__33449\ : std_logic;
signal \N__33446\ : std_logic;
signal \N__33443\ : std_logic;
signal \N__33440\ : std_logic;
signal \N__33437\ : std_logic;
signal \N__33434\ : std_logic;
signal \N__33431\ : std_logic;
signal \N__33428\ : std_logic;
signal \N__33427\ : std_logic;
signal \N__33426\ : std_logic;
signal \N__33423\ : std_logic;
signal \N__33420\ : std_logic;
signal \N__33417\ : std_logic;
signal \N__33412\ : std_logic;
signal \N__33409\ : std_logic;
signal \N__33404\ : std_logic;
signal \N__33401\ : std_logic;
signal \N__33398\ : std_logic;
signal \N__33395\ : std_logic;
signal \N__33392\ : std_logic;
signal \N__33389\ : std_logic;
signal \N__33386\ : std_logic;
signal \N__33383\ : std_logic;
signal \N__33380\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33374\ : std_logic;
signal \N__33371\ : std_logic;
signal \N__33368\ : std_logic;
signal \N__33365\ : std_logic;
signal \N__33362\ : std_logic;
signal \N__33359\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33353\ : std_logic;
signal \N__33350\ : std_logic;
signal \N__33347\ : std_logic;
signal \N__33344\ : std_logic;
signal \N__33341\ : std_logic;
signal \N__33338\ : std_logic;
signal \N__33335\ : std_logic;
signal \N__33332\ : std_logic;
signal \N__33329\ : std_logic;
signal \N__33326\ : std_logic;
signal \N__33323\ : std_logic;
signal \N__33320\ : std_logic;
signal \N__33317\ : std_logic;
signal \N__33314\ : std_logic;
signal \N__33311\ : std_logic;
signal \N__33308\ : std_logic;
signal \N__33305\ : std_logic;
signal \N__33304\ : std_logic;
signal \N__33303\ : std_logic;
signal \N__33298\ : std_logic;
signal \N__33295\ : std_logic;
signal \N__33290\ : std_logic;
signal \N__33289\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33287\ : std_logic;
signal \N__33284\ : std_logic;
signal \N__33281\ : std_logic;
signal \N__33278\ : std_logic;
signal \N__33273\ : std_logic;
signal \N__33266\ : std_logic;
signal \N__33263\ : std_logic;
signal \N__33260\ : std_logic;
signal \N__33257\ : std_logic;
signal \N__33254\ : std_logic;
signal \N__33251\ : std_logic;
signal \N__33248\ : std_logic;
signal \N__33247\ : std_logic;
signal \N__33244\ : std_logic;
signal \N__33243\ : std_logic;
signal \N__33242\ : std_logic;
signal \N__33239\ : std_logic;
signal \N__33236\ : std_logic;
signal \N__33231\ : std_logic;
signal \N__33224\ : std_logic;
signal \N__33221\ : std_logic;
signal \N__33218\ : std_logic;
signal \N__33215\ : std_logic;
signal \N__33212\ : std_logic;
signal \N__33209\ : std_logic;
signal \N__33206\ : std_logic;
signal \N__33203\ : std_logic;
signal \N__33200\ : std_logic;
signal \N__33197\ : std_logic;
signal \N__33194\ : std_logic;
signal \N__33191\ : std_logic;
signal \N__33188\ : std_logic;
signal \N__33185\ : std_logic;
signal \N__33182\ : std_logic;
signal \N__33179\ : std_logic;
signal \N__33176\ : std_logic;
signal \N__33173\ : std_logic;
signal \N__33170\ : std_logic;
signal \N__33167\ : std_logic;
signal \N__33164\ : std_logic;
signal \N__33161\ : std_logic;
signal \N__33158\ : std_logic;
signal \N__33155\ : std_logic;
signal \N__33152\ : std_logic;
signal \N__33149\ : std_logic;
signal \N__33146\ : std_logic;
signal \N__33143\ : std_logic;
signal \N__33140\ : std_logic;
signal \N__33137\ : std_logic;
signal \N__33134\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33128\ : std_logic;
signal \N__33125\ : std_logic;
signal \N__33122\ : std_logic;
signal \N__33119\ : std_logic;
signal \N__33116\ : std_logic;
signal \N__33113\ : std_logic;
signal \N__33110\ : std_logic;
signal \N__33107\ : std_logic;
signal \N__33104\ : std_logic;
signal \N__33101\ : std_logic;
signal \N__33098\ : std_logic;
signal \N__33095\ : std_logic;
signal \N__33092\ : std_logic;
signal \N__33089\ : std_logic;
signal \N__33086\ : std_logic;
signal \N__33083\ : std_logic;
signal \N__33080\ : std_logic;
signal \N__33077\ : std_logic;
signal \N__33074\ : std_logic;
signal \N__33071\ : std_logic;
signal \N__33068\ : std_logic;
signal \N__33065\ : std_logic;
signal \N__33062\ : std_logic;
signal \N__33059\ : std_logic;
signal \N__33056\ : std_logic;
signal \N__33053\ : std_logic;
signal \N__33050\ : std_logic;
signal \N__33047\ : std_logic;
signal \N__33044\ : std_logic;
signal \N__33041\ : std_logic;
signal \N__33038\ : std_logic;
signal \N__33035\ : std_logic;
signal \N__33032\ : std_logic;
signal \N__33029\ : std_logic;
signal \N__33026\ : std_logic;
signal \N__33023\ : std_logic;
signal \N__33020\ : std_logic;
signal \N__33017\ : std_logic;
signal \N__33014\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33008\ : std_logic;
signal \N__33005\ : std_logic;
signal \N__33002\ : std_logic;
signal \N__32999\ : std_logic;
signal \N__32996\ : std_logic;
signal \N__32993\ : std_logic;
signal \N__32990\ : std_logic;
signal \N__32987\ : std_logic;
signal \N__32984\ : std_logic;
signal \N__32981\ : std_logic;
signal \N__32978\ : std_logic;
signal \N__32975\ : std_logic;
signal \N__32972\ : std_logic;
signal \N__32969\ : std_logic;
signal \N__32966\ : std_logic;
signal \N__32963\ : std_logic;
signal \N__32960\ : std_logic;
signal \N__32957\ : std_logic;
signal \N__32954\ : std_logic;
signal \N__32951\ : std_logic;
signal \N__32948\ : std_logic;
signal \N__32945\ : std_logic;
signal \N__32942\ : std_logic;
signal \N__32939\ : std_logic;
signal \N__32936\ : std_logic;
signal \N__32933\ : std_logic;
signal \N__32930\ : std_logic;
signal \N__32927\ : std_logic;
signal \N__32924\ : std_logic;
signal \N__32921\ : std_logic;
signal \N__32918\ : std_logic;
signal \N__32915\ : std_logic;
signal \N__32912\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32906\ : std_logic;
signal \N__32903\ : std_logic;
signal \N__32900\ : std_logic;
signal \N__32897\ : std_logic;
signal \N__32894\ : std_logic;
signal \N__32891\ : std_logic;
signal \N__32888\ : std_logic;
signal \N__32885\ : std_logic;
signal \N__32882\ : std_logic;
signal \N__32879\ : std_logic;
signal \N__32876\ : std_logic;
signal \N__32875\ : std_logic;
signal \N__32872\ : std_logic;
signal \N__32869\ : std_logic;
signal \N__32866\ : std_logic;
signal \N__32863\ : std_logic;
signal \N__32858\ : std_logic;
signal \N__32855\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32846\ : std_logic;
signal \N__32843\ : std_logic;
signal \N__32842\ : std_logic;
signal \N__32839\ : std_logic;
signal \N__32838\ : std_logic;
signal \N__32835\ : std_logic;
signal \N__32832\ : std_logic;
signal \N__32827\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32819\ : std_logic;
signal \N__32816\ : std_logic;
signal \N__32815\ : std_logic;
signal \N__32810\ : std_logic;
signal \N__32807\ : std_logic;
signal \N__32804\ : std_logic;
signal \N__32801\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32795\ : std_logic;
signal \N__32794\ : std_logic;
signal \N__32789\ : std_logic;
signal \N__32786\ : std_logic;
signal \N__32783\ : std_logic;
signal \N__32780\ : std_logic;
signal \N__32777\ : std_logic;
signal \N__32774\ : std_logic;
signal \N__32771\ : std_logic;
signal \N__32768\ : std_logic;
signal \N__32765\ : std_logic;
signal \N__32762\ : std_logic;
signal \N__32759\ : std_logic;
signal \N__32756\ : std_logic;
signal \N__32753\ : std_logic;
signal \N__32750\ : std_logic;
signal \N__32747\ : std_logic;
signal \N__32744\ : std_logic;
signal \N__32741\ : std_logic;
signal \N__32740\ : std_logic;
signal \N__32739\ : std_logic;
signal \N__32738\ : std_logic;
signal \N__32737\ : std_logic;
signal \N__32726\ : std_logic;
signal \N__32723\ : std_logic;
signal \N__32720\ : std_logic;
signal \N__32717\ : std_logic;
signal \N__32716\ : std_logic;
signal \N__32711\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32705\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32701\ : std_logic;
signal \N__32700\ : std_logic;
signal \N__32699\ : std_logic;
signal \N__32698\ : std_logic;
signal \N__32697\ : std_logic;
signal \N__32696\ : std_logic;
signal \N__32691\ : std_logic;
signal \N__32680\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32672\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32663\ : std_logic;
signal \N__32660\ : std_logic;
signal \N__32657\ : std_logic;
signal \N__32654\ : std_logic;
signal \N__32651\ : std_logic;
signal \N__32648\ : std_logic;
signal \N__32645\ : std_logic;
signal \N__32642\ : std_logic;
signal \N__32639\ : std_logic;
signal \N__32636\ : std_logic;
signal \N__32633\ : std_logic;
signal \N__32630\ : std_logic;
signal \N__32627\ : std_logic;
signal \N__32624\ : std_logic;
signal \N__32621\ : std_logic;
signal \N__32618\ : std_logic;
signal \N__32615\ : std_logic;
signal \N__32612\ : std_logic;
signal \N__32609\ : std_logic;
signal \N__32606\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32600\ : std_logic;
signal \N__32597\ : std_logic;
signal \N__32594\ : std_logic;
signal \N__32591\ : std_logic;
signal \N__32588\ : std_logic;
signal \N__32585\ : std_logic;
signal \N__32582\ : std_logic;
signal \N__32579\ : std_logic;
signal \N__32576\ : std_logic;
signal \N__32573\ : std_logic;
signal \N__32570\ : std_logic;
signal \N__32567\ : std_logic;
signal \N__32564\ : std_logic;
signal \N__32561\ : std_logic;
signal \N__32558\ : std_logic;
signal \N__32555\ : std_logic;
signal \N__32552\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32546\ : std_logic;
signal \N__32543\ : std_logic;
signal \N__32540\ : std_logic;
signal \N__32539\ : std_logic;
signal \N__32538\ : std_logic;
signal \N__32535\ : std_logic;
signal \N__32532\ : std_logic;
signal \N__32529\ : std_logic;
signal \N__32526\ : std_logic;
signal \N__32521\ : std_logic;
signal \N__32518\ : std_logic;
signal \N__32515\ : std_logic;
signal \N__32510\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32506\ : std_logic;
signal \N__32505\ : std_logic;
signal \N__32504\ : std_logic;
signal \N__32499\ : std_logic;
signal \N__32496\ : std_logic;
signal \N__32493\ : std_logic;
signal \N__32486\ : std_logic;
signal \N__32483\ : std_logic;
signal \N__32480\ : std_logic;
signal \N__32477\ : std_logic;
signal \N__32474\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32468\ : std_logic;
signal \N__32465\ : std_logic;
signal \N__32462\ : std_logic;
signal \N__32459\ : std_logic;
signal \N__32456\ : std_logic;
signal \N__32453\ : std_logic;
signal \N__32450\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32444\ : std_logic;
signal \N__32441\ : std_logic;
signal \N__32438\ : std_logic;
signal \N__32435\ : std_logic;
signal \N__32432\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32426\ : std_logic;
signal \N__32423\ : std_logic;
signal \N__32420\ : std_logic;
signal \N__32417\ : std_logic;
signal \N__32414\ : std_logic;
signal \N__32411\ : std_logic;
signal \N__32408\ : std_logic;
signal \N__32405\ : std_logic;
signal \N__32402\ : std_logic;
signal \N__32399\ : std_logic;
signal \N__32396\ : std_logic;
signal \N__32393\ : std_logic;
signal \N__32392\ : std_logic;
signal \N__32389\ : std_logic;
signal \N__32386\ : std_logic;
signal \N__32385\ : std_logic;
signal \N__32382\ : std_logic;
signal \N__32381\ : std_logic;
signal \N__32380\ : std_logic;
signal \N__32375\ : std_logic;
signal \N__32372\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32362\ : std_logic;
signal \N__32357\ : std_logic;
signal \N__32356\ : std_logic;
signal \N__32353\ : std_logic;
signal \N__32352\ : std_logic;
signal \N__32351\ : std_logic;
signal \N__32350\ : std_logic;
signal \N__32347\ : std_logic;
signal \N__32342\ : std_logic;
signal \N__32335\ : std_logic;
signal \N__32330\ : std_logic;
signal \N__32329\ : std_logic;
signal \N__32328\ : std_logic;
signal \N__32327\ : std_logic;
signal \N__32324\ : std_logic;
signal \N__32321\ : std_logic;
signal \N__32316\ : std_logic;
signal \N__32309\ : std_logic;
signal \N__32308\ : std_logic;
signal \N__32307\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32305\ : std_logic;
signal \N__32304\ : std_logic;
signal \N__32301\ : std_logic;
signal \N__32300\ : std_logic;
signal \N__32293\ : std_logic;
signal \N__32288\ : std_logic;
signal \N__32283\ : std_logic;
signal \N__32276\ : std_logic;
signal \N__32273\ : std_logic;
signal \N__32270\ : std_logic;
signal \N__32267\ : std_logic;
signal \N__32264\ : std_logic;
signal \N__32261\ : std_logic;
signal \N__32258\ : std_logic;
signal \N__32255\ : std_logic;
signal \N__32252\ : std_logic;
signal \N__32251\ : std_logic;
signal \N__32250\ : std_logic;
signal \N__32247\ : std_logic;
signal \N__32246\ : std_logic;
signal \N__32243\ : std_logic;
signal \N__32240\ : std_logic;
signal \N__32237\ : std_logic;
signal \N__32234\ : std_logic;
signal \N__32231\ : std_logic;
signal \N__32228\ : std_logic;
signal \N__32219\ : std_logic;
signal \N__32218\ : std_logic;
signal \N__32217\ : std_logic;
signal \N__32214\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32203\ : std_logic;
signal \N__32200\ : std_logic;
signal \N__32197\ : std_logic;
signal \N__32194\ : std_logic;
signal \N__32191\ : std_logic;
signal \N__32188\ : std_logic;
signal \N__32185\ : std_logic;
signal \N__32182\ : std_logic;
signal \N__32179\ : std_logic;
signal \N__32176\ : std_logic;
signal \N__32171\ : std_logic;
signal \N__32168\ : std_logic;
signal \N__32167\ : std_logic;
signal \N__32166\ : std_logic;
signal \N__32163\ : std_logic;
signal \N__32158\ : std_logic;
signal \N__32153\ : std_logic;
signal \N__32152\ : std_logic;
signal \N__32151\ : std_logic;
signal \N__32150\ : std_logic;
signal \N__32145\ : std_logic;
signal \N__32140\ : std_logic;
signal \N__32135\ : std_logic;
signal \N__32134\ : std_logic;
signal \N__32133\ : std_logic;
signal \N__32130\ : std_logic;
signal \N__32127\ : std_logic;
signal \N__32126\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32114\ : std_logic;
signal \N__32111\ : std_logic;
signal \N__32106\ : std_logic;
signal \N__32103\ : std_logic;
signal \N__32098\ : std_logic;
signal \N__32095\ : std_logic;
signal \N__32090\ : std_logic;
signal \N__32089\ : std_logic;
signal \N__32088\ : std_logic;
signal \N__32087\ : std_logic;
signal \N__32086\ : std_logic;
signal \N__32085\ : std_logic;
signal \N__32084\ : std_logic;
signal \N__32083\ : std_logic;
signal \N__32082\ : std_logic;
signal \N__32081\ : std_logic;
signal \N__32080\ : std_logic;
signal \N__32079\ : std_logic;
signal \N__32078\ : std_logic;
signal \N__32077\ : std_logic;
signal \N__32076\ : std_logic;
signal \N__32075\ : std_logic;
signal \N__32074\ : std_logic;
signal \N__32073\ : std_logic;
signal \N__32072\ : std_logic;
signal \N__32071\ : std_logic;
signal \N__32070\ : std_logic;
signal \N__32069\ : std_logic;
signal \N__32068\ : std_logic;
signal \N__32067\ : std_logic;
signal \N__32066\ : std_logic;
signal \N__32065\ : std_logic;
signal \N__32064\ : std_logic;
signal \N__32063\ : std_logic;
signal \N__32062\ : std_logic;
signal \N__32061\ : std_logic;
signal \N__32056\ : std_logic;
signal \N__32047\ : std_logic;
signal \N__32038\ : std_logic;
signal \N__32029\ : std_logic;
signal \N__32020\ : std_logic;
signal \N__32011\ : std_logic;
signal \N__32002\ : std_logic;
signal \N__31993\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31983\ : std_logic;
signal \N__31978\ : std_logic;
signal \N__31973\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31955\ : std_logic;
signal \N__31952\ : std_logic;
signal \N__31949\ : std_logic;
signal \N__31946\ : std_logic;
signal \N__31943\ : std_logic;
signal \N__31940\ : std_logic;
signal \N__31937\ : std_logic;
signal \N__31934\ : std_logic;
signal \N__31931\ : std_logic;
signal \N__31928\ : std_logic;
signal \N__31925\ : std_logic;
signal \N__31922\ : std_logic;
signal \N__31919\ : std_logic;
signal \N__31916\ : std_logic;
signal \N__31913\ : std_logic;
signal \N__31910\ : std_logic;
signal \N__31907\ : std_logic;
signal \N__31904\ : std_logic;
signal \N__31903\ : std_logic;
signal \N__31900\ : std_logic;
signal \N__31897\ : std_logic;
signal \N__31894\ : std_logic;
signal \N__31891\ : std_logic;
signal \N__31886\ : std_logic;
signal \N__31883\ : std_logic;
signal \N__31880\ : std_logic;
signal \N__31877\ : std_logic;
signal \N__31874\ : std_logic;
signal \N__31871\ : std_logic;
signal \N__31868\ : std_logic;
signal \N__31867\ : std_logic;
signal \N__31866\ : std_logic;
signal \N__31863\ : std_logic;
signal \N__31860\ : std_logic;
signal \N__31859\ : std_logic;
signal \N__31856\ : std_logic;
signal \N__31853\ : std_logic;
signal \N__31850\ : std_logic;
signal \N__31847\ : std_logic;
signal \N__31842\ : std_logic;
signal \N__31837\ : std_logic;
signal \N__31832\ : std_logic;
signal \N__31829\ : std_logic;
signal \N__31826\ : std_logic;
signal \N__31825\ : std_logic;
signal \N__31824\ : std_logic;
signal \N__31823\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31817\ : std_logic;
signal \N__31814\ : std_logic;
signal \N__31811\ : std_logic;
signal \N__31806\ : std_logic;
signal \N__31803\ : std_logic;
signal \N__31796\ : std_logic;
signal \N__31793\ : std_logic;
signal \N__31790\ : std_logic;
signal \N__31787\ : std_logic;
signal \N__31784\ : std_logic;
signal \N__31783\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31779\ : std_logic;
signal \N__31774\ : std_logic;
signal \N__31769\ : std_logic;
signal \N__31768\ : std_logic;
signal \N__31765\ : std_logic;
signal \N__31762\ : std_logic;
signal \N__31759\ : std_logic;
signal \N__31756\ : std_logic;
signal \N__31751\ : std_logic;
signal \N__31750\ : std_logic;
signal \N__31749\ : std_logic;
signal \N__31748\ : std_logic;
signal \N__31743\ : std_logic;
signal \N__31740\ : std_logic;
signal \N__31737\ : std_logic;
signal \N__31730\ : std_logic;
signal \N__31727\ : std_logic;
signal \N__31724\ : std_logic;
signal \N__31721\ : std_logic;
signal \N__31718\ : std_logic;
signal \N__31715\ : std_logic;
signal \N__31712\ : std_logic;
signal \N__31709\ : std_logic;
signal \N__31706\ : std_logic;
signal \N__31705\ : std_logic;
signal \N__31704\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31698\ : std_logic;
signal \N__31695\ : std_logic;
signal \N__31692\ : std_logic;
signal \N__31689\ : std_logic;
signal \N__31686\ : std_logic;
signal \N__31679\ : std_logic;
signal \N__31676\ : std_logic;
signal \N__31675\ : std_logic;
signal \N__31672\ : std_logic;
signal \N__31671\ : std_logic;
signal \N__31668\ : std_logic;
signal \N__31665\ : std_logic;
signal \N__31662\ : std_logic;
signal \N__31655\ : std_logic;
signal \N__31654\ : std_logic;
signal \N__31651\ : std_logic;
signal \N__31648\ : std_logic;
signal \N__31645\ : std_logic;
signal \N__31642\ : std_logic;
signal \N__31639\ : std_logic;
signal \N__31636\ : std_logic;
signal \N__31631\ : std_logic;
signal \N__31628\ : std_logic;
signal \N__31627\ : std_logic;
signal \N__31626\ : std_logic;
signal \N__31623\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31617\ : std_logic;
signal \N__31614\ : std_logic;
signal \N__31611\ : std_logic;
signal \N__31608\ : std_logic;
signal \N__31603\ : std_logic;
signal \N__31600\ : std_logic;
signal \N__31597\ : std_logic;
signal \N__31592\ : std_logic;
signal \N__31589\ : std_logic;
signal \N__31588\ : std_logic;
signal \N__31587\ : std_logic;
signal \N__31584\ : std_logic;
signal \N__31581\ : std_logic;
signal \N__31578\ : std_logic;
signal \N__31573\ : std_logic;
signal \N__31572\ : std_logic;
signal \N__31569\ : std_logic;
signal \N__31566\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31556\ : std_logic;
signal \N__31553\ : std_logic;
signal \N__31550\ : std_logic;
signal \N__31549\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31545\ : std_logic;
signal \N__31544\ : std_logic;
signal \N__31541\ : std_logic;
signal \N__31538\ : std_logic;
signal \N__31535\ : std_logic;
signal \N__31532\ : std_logic;
signal \N__31529\ : std_logic;
signal \N__31526\ : std_logic;
signal \N__31521\ : std_logic;
signal \N__31518\ : std_logic;
signal \N__31515\ : std_logic;
signal \N__31508\ : std_logic;
signal \N__31507\ : std_logic;
signal \N__31504\ : std_logic;
signal \N__31503\ : std_logic;
signal \N__31502\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31496\ : std_logic;
signal \N__31491\ : std_logic;
signal \N__31488\ : std_logic;
signal \N__31481\ : std_logic;
signal \N__31478\ : std_logic;
signal \N__31475\ : std_logic;
signal \N__31472\ : std_logic;
signal \N__31469\ : std_logic;
signal \N__31466\ : std_logic;
signal \N__31463\ : std_logic;
signal \N__31460\ : std_logic;
signal \N__31457\ : std_logic;
signal \N__31454\ : std_logic;
signal \N__31451\ : std_logic;
signal \N__31448\ : std_logic;
signal \N__31445\ : std_logic;
signal \N__31442\ : std_logic;
signal \N__31439\ : std_logic;
signal \N__31436\ : std_logic;
signal \N__31435\ : std_logic;
signal \N__31432\ : std_logic;
signal \N__31429\ : std_logic;
signal \N__31426\ : std_logic;
signal \N__31423\ : std_logic;
signal \N__31418\ : std_logic;
signal \N__31417\ : std_logic;
signal \N__31414\ : std_logic;
signal \N__31411\ : std_logic;
signal \N__31408\ : std_logic;
signal \N__31405\ : std_logic;
signal \N__31400\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31394\ : std_logic;
signal \N__31391\ : std_logic;
signal \N__31388\ : std_logic;
signal \N__31385\ : std_logic;
signal \N__31382\ : std_logic;
signal \N__31379\ : std_logic;
signal \N__31376\ : std_logic;
signal \N__31373\ : std_logic;
signal \N__31370\ : std_logic;
signal \N__31367\ : std_logic;
signal \N__31364\ : std_logic;
signal \N__31361\ : std_logic;
signal \N__31358\ : std_logic;
signal \N__31355\ : std_logic;
signal \N__31352\ : std_logic;
signal \N__31349\ : std_logic;
signal \N__31346\ : std_logic;
signal \N__31343\ : std_logic;
signal \N__31340\ : std_logic;
signal \N__31337\ : std_logic;
signal \N__31334\ : std_logic;
signal \N__31331\ : std_logic;
signal \N__31328\ : std_logic;
signal \N__31325\ : std_logic;
signal \N__31322\ : std_logic;
signal \N__31319\ : std_logic;
signal \N__31316\ : std_logic;
signal \N__31313\ : std_logic;
signal \N__31310\ : std_logic;
signal \N__31307\ : std_logic;
signal \N__31304\ : std_logic;
signal \N__31301\ : std_logic;
signal \N__31298\ : std_logic;
signal \N__31295\ : std_logic;
signal \N__31292\ : std_logic;
signal \N__31289\ : std_logic;
signal \N__31286\ : std_logic;
signal \N__31283\ : std_logic;
signal \N__31280\ : std_logic;
signal \N__31277\ : std_logic;
signal \N__31274\ : std_logic;
signal \N__31271\ : std_logic;
signal \N__31268\ : std_logic;
signal \N__31265\ : std_logic;
signal \N__31262\ : std_logic;
signal \N__31259\ : std_logic;
signal \N__31256\ : std_logic;
signal \N__31253\ : std_logic;
signal \N__31250\ : std_logic;
signal \N__31247\ : std_logic;
signal \N__31244\ : std_logic;
signal \N__31241\ : std_logic;
signal \N__31238\ : std_logic;
signal \N__31235\ : std_logic;
signal \N__31232\ : std_logic;
signal \N__31229\ : std_logic;
signal \N__31228\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31226\ : std_logic;
signal \N__31225\ : std_logic;
signal \N__31224\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31215\ : std_logic;
signal \N__31212\ : std_logic;
signal \N__31209\ : std_logic;
signal \N__31206\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31200\ : std_logic;
signal \N__31197\ : std_logic;
signal \N__31194\ : std_logic;
signal \N__31191\ : std_logic;
signal \N__31188\ : std_logic;
signal \N__31185\ : std_logic;
signal \N__31180\ : std_logic;
signal \N__31177\ : std_logic;
signal \N__31174\ : std_logic;
signal \N__31163\ : std_logic;
signal \N__31160\ : std_logic;
signal \N__31157\ : std_logic;
signal \N__31154\ : std_logic;
signal \N__31151\ : std_logic;
signal \N__31148\ : std_logic;
signal \N__31145\ : std_logic;
signal \N__31142\ : std_logic;
signal \N__31139\ : std_logic;
signal \N__31138\ : std_logic;
signal \N__31135\ : std_logic;
signal \N__31132\ : std_logic;
signal \N__31129\ : std_logic;
signal \N__31124\ : std_logic;
signal \N__31121\ : std_logic;
signal \N__31118\ : std_logic;
signal \N__31115\ : std_logic;
signal \N__31112\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31110\ : std_logic;
signal \N__31107\ : std_logic;
signal \N__31106\ : std_logic;
signal \N__31101\ : std_logic;
signal \N__31098\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31092\ : std_logic;
signal \N__31085\ : std_logic;
signal \N__31082\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31072\ : std_logic;
signal \N__31071\ : std_logic;
signal \N__31070\ : std_logic;
signal \N__31067\ : std_logic;
signal \N__31062\ : std_logic;
signal \N__31059\ : std_logic;
signal \N__31054\ : std_logic;
signal \N__31051\ : std_logic;
signal \N__31046\ : std_logic;
signal \N__31045\ : std_logic;
signal \N__31042\ : std_logic;
signal \N__31041\ : std_logic;
signal \N__31034\ : std_logic;
signal \N__31033\ : std_logic;
signal \N__31030\ : std_logic;
signal \N__31027\ : std_logic;
signal \N__31022\ : std_logic;
signal \N__31019\ : std_logic;
signal \N__31016\ : std_logic;
signal \N__31013\ : std_logic;
signal \N__31010\ : std_logic;
signal \N__31007\ : std_logic;
signal \N__31004\ : std_logic;
signal \N__31003\ : std_logic;
signal \N__31002\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30993\ : std_logic;
signal \N__30992\ : std_logic;
signal \N__30989\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30981\ : std_logic;
signal \N__30978\ : std_logic;
signal \N__30973\ : std_logic;
signal \N__30968\ : std_logic;
signal \N__30965\ : std_logic;
signal \N__30964\ : std_logic;
signal \N__30963\ : std_logic;
signal \N__30960\ : std_logic;
signal \N__30955\ : std_logic;
signal \N__30954\ : std_logic;
signal \N__30951\ : std_logic;
signal \N__30948\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30938\ : std_logic;
signal \N__30935\ : std_logic;
signal \N__30932\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30926\ : std_logic;
signal \N__30923\ : std_logic;
signal \N__30920\ : std_logic;
signal \N__30917\ : std_logic;
signal \N__30914\ : std_logic;
signal \N__30911\ : std_logic;
signal \N__30908\ : std_logic;
signal \N__30905\ : std_logic;
signal \N__30902\ : std_logic;
signal \N__30899\ : std_logic;
signal \N__30896\ : std_logic;
signal \N__30893\ : std_logic;
signal \N__30890\ : std_logic;
signal \N__30887\ : std_logic;
signal \N__30884\ : std_logic;
signal \N__30883\ : std_logic;
signal \N__30880\ : std_logic;
signal \N__30879\ : std_logic;
signal \N__30876\ : std_logic;
signal \N__30873\ : std_logic;
signal \N__30870\ : std_logic;
signal \N__30869\ : std_logic;
signal \N__30864\ : std_logic;
signal \N__30861\ : std_logic;
signal \N__30858\ : std_logic;
signal \N__30855\ : std_logic;
signal \N__30852\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30842\ : std_logic;
signal \N__30839\ : std_logic;
signal \N__30838\ : std_logic;
signal \N__30835\ : std_logic;
signal \N__30832\ : std_logic;
signal \N__30831\ : std_logic;
signal \N__30828\ : std_logic;
signal \N__30827\ : std_logic;
signal \N__30824\ : std_logic;
signal \N__30821\ : std_logic;
signal \N__30818\ : std_logic;
signal \N__30815\ : std_logic;
signal \N__30812\ : std_logic;
signal \N__30809\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30797\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30788\ : std_logic;
signal \N__30785\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30776\ : std_logic;
signal \N__30773\ : std_logic;
signal \N__30772\ : std_logic;
signal \N__30771\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30763\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30759\ : std_logic;
signal \N__30756\ : std_logic;
signal \N__30753\ : std_logic;
signal \N__30750\ : std_logic;
signal \N__30745\ : std_logic;
signal \N__30740\ : std_logic;
signal \N__30739\ : std_logic;
signal \N__30738\ : std_logic;
signal \N__30737\ : std_logic;
signal \N__30730\ : std_logic;
signal \N__30727\ : std_logic;
signal \N__30724\ : std_logic;
signal \N__30721\ : std_logic;
signal \N__30716\ : std_logic;
signal \N__30715\ : std_logic;
signal \N__30712\ : std_logic;
signal \N__30709\ : std_logic;
signal \N__30708\ : std_logic;
signal \N__30707\ : std_logic;
signal \N__30704\ : std_logic;
signal \N__30701\ : std_logic;
signal \N__30698\ : std_logic;
signal \N__30695\ : std_logic;
signal \N__30688\ : std_logic;
signal \N__30685\ : std_logic;
signal \N__30680\ : std_logic;
signal \N__30679\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30673\ : std_logic;
signal \N__30672\ : std_logic;
signal \N__30669\ : std_logic;
signal \N__30664\ : std_logic;
signal \N__30663\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30650\ : std_logic;
signal \N__30647\ : std_logic;
signal \N__30644\ : std_logic;
signal \N__30641\ : std_logic;
signal \N__30638\ : std_logic;
signal \N__30635\ : std_logic;
signal \N__30632\ : std_logic;
signal \N__30631\ : std_logic;
signal \N__30630\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30624\ : std_logic;
signal \N__30621\ : std_logic;
signal \N__30618\ : std_logic;
signal \N__30615\ : std_logic;
signal \N__30612\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30604\ : std_logic;
signal \N__30603\ : std_logic;
signal \N__30600\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30598\ : std_logic;
signal \N__30595\ : std_logic;
signal \N__30594\ : std_logic;
signal \N__30591\ : std_logic;
signal \N__30590\ : std_logic;
signal \N__30587\ : std_logic;
signal \N__30584\ : std_logic;
signal \N__30575\ : std_logic;
signal \N__30574\ : std_logic;
signal \N__30571\ : std_logic;
signal \N__30564\ : std_logic;
signal \N__30561\ : std_logic;
signal \N__30560\ : std_logic;
signal \N__30557\ : std_logic;
signal \N__30554\ : std_logic;
signal \N__30551\ : std_logic;
signal \N__30548\ : std_logic;
signal \N__30539\ : std_logic;
signal \N__30536\ : std_logic;
signal \N__30533\ : std_logic;
signal \N__30530\ : std_logic;
signal \N__30529\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30523\ : std_logic;
signal \N__30520\ : std_logic;
signal \N__30517\ : std_logic;
signal \N__30514\ : std_logic;
signal \N__30511\ : std_logic;
signal \N__30508\ : std_logic;
signal \N__30505\ : std_logic;
signal \N__30500\ : std_logic;
signal \N__30499\ : std_logic;
signal \N__30496\ : std_logic;
signal \N__30493\ : std_logic;
signal \N__30490\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30484\ : std_logic;
signal \N__30481\ : std_logic;
signal \N__30476\ : std_logic;
signal \N__30473\ : std_logic;
signal \N__30470\ : std_logic;
signal \N__30467\ : std_logic;
signal \N__30464\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30462\ : std_logic;
signal \N__30459\ : std_logic;
signal \N__30456\ : std_logic;
signal \N__30453\ : std_logic;
signal \N__30452\ : std_logic;
signal \N__30449\ : std_logic;
signal \N__30446\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30440\ : std_logic;
signal \N__30435\ : std_logic;
signal \N__30430\ : std_logic;
signal \N__30425\ : std_logic;
signal \N__30424\ : std_logic;
signal \N__30421\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30417\ : std_logic;
signal \N__30416\ : std_logic;
signal \N__30413\ : std_logic;
signal \N__30410\ : std_logic;
signal \N__30407\ : std_logic;
signal \N__30404\ : std_logic;
signal \N__30401\ : std_logic;
signal \N__30398\ : std_logic;
signal \N__30395\ : std_logic;
signal \N__30392\ : std_logic;
signal \N__30383\ : std_logic;
signal \N__30380\ : std_logic;
signal \N__30377\ : std_logic;
signal \N__30374\ : std_logic;
signal \N__30371\ : std_logic;
signal \N__30368\ : std_logic;
signal \N__30365\ : std_logic;
signal \N__30362\ : std_logic;
signal \N__30359\ : std_logic;
signal \N__30358\ : std_logic;
signal \N__30357\ : std_logic;
signal \N__30354\ : std_logic;
signal \N__30351\ : std_logic;
signal \N__30350\ : std_logic;
signal \N__30347\ : std_logic;
signal \N__30344\ : std_logic;
signal \N__30341\ : std_logic;
signal \N__30338\ : std_logic;
signal \N__30335\ : std_logic;
signal \N__30332\ : std_logic;
signal \N__30325\ : std_logic;
signal \N__30320\ : std_logic;
signal \N__30319\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30313\ : std_logic;
signal \N__30312\ : std_logic;
signal \N__30307\ : std_logic;
signal \N__30304\ : std_logic;
signal \N__30303\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30297\ : std_logic;
signal \N__30294\ : std_logic;
signal \N__30287\ : std_logic;
signal \N__30284\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30272\ : std_logic;
signal \N__30271\ : std_logic;
signal \N__30270\ : std_logic;
signal \N__30269\ : std_logic;
signal \N__30266\ : std_logic;
signal \N__30263\ : std_logic;
signal \N__30260\ : std_logic;
signal \N__30257\ : std_logic;
signal \N__30254\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30246\ : std_logic;
signal \N__30239\ : std_logic;
signal \N__30236\ : std_logic;
signal \N__30235\ : std_logic;
signal \N__30234\ : std_logic;
signal \N__30233\ : std_logic;
signal \N__30226\ : std_logic;
signal \N__30223\ : std_logic;
signal \N__30220\ : std_logic;
signal \N__30217\ : std_logic;
signal \N__30212\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30208\ : std_logic;
signal \N__30207\ : std_logic;
signal \N__30204\ : std_logic;
signal \N__30201\ : std_logic;
signal \N__30198\ : std_logic;
signal \N__30197\ : std_logic;
signal \N__30194\ : std_logic;
signal \N__30191\ : std_logic;
signal \N__30188\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30182\ : std_logic;
signal \N__30177\ : std_logic;
signal \N__30174\ : std_logic;
signal \N__30167\ : std_logic;
signal \N__30166\ : std_logic;
signal \N__30165\ : std_logic;
signal \N__30164\ : std_logic;
signal \N__30157\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30151\ : std_logic;
signal \N__30148\ : std_logic;
signal \N__30145\ : std_logic;
signal \N__30142\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30134\ : std_logic;
signal \N__30131\ : std_logic;
signal \N__30128\ : std_logic;
signal \N__30125\ : std_logic;
signal \N__30122\ : std_logic;
signal \N__30121\ : std_logic;
signal \N__30120\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30112\ : std_logic;
signal \N__30111\ : std_logic;
signal \N__30108\ : std_logic;
signal \N__30105\ : std_logic;
signal \N__30102\ : std_logic;
signal \N__30099\ : std_logic;
signal \N__30096\ : std_logic;
signal \N__30093\ : std_logic;
signal \N__30086\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30080\ : std_logic;
signal \N__30077\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30070\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30065\ : std_logic;
signal \N__30062\ : std_logic;
signal \N__30059\ : std_logic;
signal \N__30056\ : std_logic;
signal \N__30053\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30041\ : std_logic;
signal \N__30038\ : std_logic;
signal \N__30037\ : std_logic;
signal \N__30034\ : std_logic;
signal \N__30031\ : std_logic;
signal \N__30030\ : std_logic;
signal \N__30029\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30015\ : std_logic;
signal \N__30012\ : std_logic;
signal \N__30009\ : std_logic;
signal \N__30002\ : std_logic;
signal \N__29999\ : std_logic;
signal \N__29996\ : std_logic;
signal \N__29993\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29987\ : std_logic;
signal \N__29984\ : std_logic;
signal \N__29981\ : std_logic;
signal \N__29978\ : std_logic;
signal \N__29975\ : std_logic;
signal \N__29972\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29968\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29964\ : std_logic;
signal \N__29961\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29957\ : std_logic;
signal \N__29952\ : std_logic;
signal \N__29949\ : std_logic;
signal \N__29946\ : std_logic;
signal \N__29943\ : std_logic;
signal \N__29938\ : std_logic;
signal \N__29933\ : std_logic;
signal \N__29930\ : std_logic;
signal \N__29929\ : std_logic;
signal \N__29926\ : std_logic;
signal \N__29925\ : std_logic;
signal \N__29922\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29918\ : std_logic;
signal \N__29915\ : std_logic;
signal \N__29912\ : std_logic;
signal \N__29909\ : std_logic;
signal \N__29904\ : std_logic;
signal \N__29901\ : std_logic;
signal \N__29898\ : std_logic;
signal \N__29891\ : std_logic;
signal \N__29888\ : std_logic;
signal \N__29885\ : std_logic;
signal \N__29882\ : std_logic;
signal \N__29881\ : std_logic;
signal \N__29880\ : std_logic;
signal \N__29877\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29873\ : std_logic;
signal \N__29870\ : std_logic;
signal \N__29865\ : std_logic;
signal \N__29862\ : std_logic;
signal \N__29859\ : std_logic;
signal \N__29856\ : std_logic;
signal \N__29853\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29845\ : std_logic;
signal \N__29842\ : std_logic;
signal \N__29839\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29837\ : std_logic;
signal \N__29834\ : std_logic;
signal \N__29831\ : std_logic;
signal \N__29828\ : std_logic;
signal \N__29825\ : std_logic;
signal \N__29822\ : std_logic;
signal \N__29817\ : std_logic;
signal \N__29814\ : std_logic;
signal \N__29807\ : std_logic;
signal \N__29804\ : std_logic;
signal \N__29801\ : std_logic;
signal \N__29798\ : std_logic;
signal \N__29795\ : std_logic;
signal \N__29792\ : std_logic;
signal \N__29789\ : std_logic;
signal \N__29786\ : std_logic;
signal \N__29783\ : std_logic;
signal \N__29780\ : std_logic;
signal \N__29779\ : std_logic;
signal \N__29778\ : std_logic;
signal \N__29771\ : std_logic;
signal \N__29770\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29764\ : std_logic;
signal \N__29761\ : std_logic;
signal \N__29758\ : std_logic;
signal \N__29753\ : std_logic;
signal \N__29750\ : std_logic;
signal \N__29747\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29741\ : std_logic;
signal \N__29738\ : std_logic;
signal \N__29737\ : std_logic;
signal \N__29736\ : std_logic;
signal \N__29733\ : std_logic;
signal \N__29728\ : std_logic;
signal \N__29725\ : std_logic;
signal \N__29722\ : std_logic;
signal \N__29721\ : std_logic;
signal \N__29718\ : std_logic;
signal \N__29715\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29702\ : std_logic;
signal \N__29699\ : std_logic;
signal \N__29696\ : std_logic;
signal \N__29693\ : std_logic;
signal \N__29690\ : std_logic;
signal \N__29687\ : std_logic;
signal \N__29684\ : std_logic;
signal \N__29681\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29679\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29671\ : std_logic;
signal \N__29670\ : std_logic;
signal \N__29667\ : std_logic;
signal \N__29664\ : std_logic;
signal \N__29661\ : std_logic;
signal \N__29656\ : std_logic;
signal \N__29653\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29645\ : std_logic;
signal \N__29642\ : std_logic;
signal \N__29641\ : std_logic;
signal \N__29640\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29632\ : std_logic;
signal \N__29631\ : std_logic;
signal \N__29628\ : std_logic;
signal \N__29625\ : std_logic;
signal \N__29622\ : std_logic;
signal \N__29615\ : std_logic;
signal \N__29614\ : std_logic;
signal \N__29611\ : std_logic;
signal \N__29608\ : std_logic;
signal \N__29605\ : std_logic;
signal \N__29604\ : std_logic;
signal \N__29599\ : std_logic;
signal \N__29596\ : std_logic;
signal \N__29593\ : std_logic;
signal \N__29590\ : std_logic;
signal \N__29585\ : std_logic;
signal \N__29582\ : std_logic;
signal \N__29581\ : std_logic;
signal \N__29578\ : std_logic;
signal \N__29575\ : std_logic;
signal \N__29570\ : std_logic;
signal \N__29569\ : std_logic;
signal \N__29566\ : std_logic;
signal \N__29563\ : std_logic;
signal \N__29558\ : std_logic;
signal \N__29555\ : std_logic;
signal \N__29552\ : std_logic;
signal \N__29549\ : std_logic;
signal \N__29548\ : std_logic;
signal \N__29545\ : std_logic;
signal \N__29542\ : std_logic;
signal \N__29537\ : std_logic;
signal \N__29534\ : std_logic;
signal \N__29531\ : std_logic;
signal \N__29530\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29526\ : std_logic;
signal \N__29523\ : std_logic;
signal \N__29520\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29514\ : std_logic;
signal \N__29511\ : std_logic;
signal \N__29508\ : std_logic;
signal \N__29505\ : std_logic;
signal \N__29502\ : std_logic;
signal \N__29499\ : std_logic;
signal \N__29492\ : std_logic;
signal \N__29489\ : std_logic;
signal \N__29488\ : std_logic;
signal \N__29487\ : std_logic;
signal \N__29484\ : std_logic;
signal \N__29479\ : std_logic;
signal \N__29476\ : std_logic;
signal \N__29473\ : std_logic;
signal \N__29472\ : std_logic;
signal \N__29469\ : std_logic;
signal \N__29466\ : std_logic;
signal \N__29463\ : std_logic;
signal \N__29456\ : std_logic;
signal \N__29453\ : std_logic;
signal \N__29452\ : std_logic;
signal \N__29451\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29443\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29433\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29427\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29414\ : std_logic;
signal \N__29411\ : std_logic;
signal \N__29408\ : std_logic;
signal \N__29407\ : std_logic;
signal \N__29404\ : std_logic;
signal \N__29403\ : std_logic;
signal \N__29400\ : std_logic;
signal \N__29397\ : std_logic;
signal \N__29392\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29388\ : std_logic;
signal \N__29385\ : std_logic;
signal \N__29382\ : std_logic;
signal \N__29379\ : std_logic;
signal \N__29376\ : std_logic;
signal \N__29373\ : std_logic;
signal \N__29366\ : std_logic;
signal \N__29363\ : std_logic;
signal \N__29360\ : std_logic;
signal \N__29357\ : std_logic;
signal \N__29354\ : std_logic;
signal \N__29351\ : std_logic;
signal \N__29348\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29342\ : std_logic;
signal \N__29339\ : std_logic;
signal \N__29336\ : std_logic;
signal \N__29333\ : std_logic;
signal \N__29330\ : std_logic;
signal \N__29327\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29322\ : std_logic;
signal \N__29319\ : std_logic;
signal \N__29316\ : std_logic;
signal \N__29313\ : std_logic;
signal \N__29306\ : std_logic;
signal \N__29303\ : std_logic;
signal \N__29300\ : std_logic;
signal \N__29297\ : std_logic;
signal \N__29294\ : std_logic;
signal \N__29293\ : std_logic;
signal \N__29290\ : std_logic;
signal \N__29287\ : std_logic;
signal \N__29282\ : std_logic;
signal \N__29279\ : std_logic;
signal \N__29278\ : std_logic;
signal \N__29275\ : std_logic;
signal \N__29272\ : std_logic;
signal \N__29269\ : std_logic;
signal \N__29264\ : std_logic;
signal \N__29261\ : std_logic;
signal \N__29258\ : std_logic;
signal \N__29255\ : std_logic;
signal \N__29254\ : std_logic;
signal \N__29251\ : std_logic;
signal \N__29248\ : std_logic;
signal \N__29245\ : std_logic;
signal \N__29242\ : std_logic;
signal \N__29237\ : std_logic;
signal \N__29234\ : std_logic;
signal \N__29231\ : std_logic;
signal \N__29228\ : std_logic;
signal \N__29225\ : std_logic;
signal \N__29222\ : std_logic;
signal \N__29221\ : std_logic;
signal \N__29218\ : std_logic;
signal \N__29215\ : std_logic;
signal \N__29212\ : std_logic;
signal \N__29207\ : std_logic;
signal \N__29204\ : std_logic;
signal \N__29201\ : std_logic;
signal \N__29198\ : std_logic;
signal \N__29195\ : std_logic;
signal \N__29194\ : std_logic;
signal \N__29191\ : std_logic;
signal \N__29188\ : std_logic;
signal \N__29185\ : std_logic;
signal \N__29180\ : std_logic;
signal \N__29177\ : std_logic;
signal \N__29174\ : std_logic;
signal \N__29171\ : std_logic;
signal \N__29168\ : std_logic;
signal \N__29167\ : std_logic;
signal \N__29164\ : std_logic;
signal \N__29161\ : std_logic;
signal \N__29158\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29150\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29141\ : std_logic;
signal \N__29140\ : std_logic;
signal \N__29137\ : std_logic;
signal \N__29134\ : std_logic;
signal \N__29131\ : std_logic;
signal \N__29126\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29120\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29113\ : std_logic;
signal \N__29110\ : std_logic;
signal \N__29107\ : std_logic;
signal \N__29104\ : std_logic;
signal \N__29099\ : std_logic;
signal \N__29096\ : std_logic;
signal \N__29093\ : std_logic;
signal \N__29090\ : std_logic;
signal \N__29087\ : std_logic;
signal \N__29084\ : std_logic;
signal \N__29081\ : std_logic;
signal \N__29078\ : std_logic;
signal \N__29075\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29063\ : std_logic;
signal \N__29060\ : std_logic;
signal \N__29057\ : std_logic;
signal \N__29054\ : std_logic;
signal \N__29051\ : std_logic;
signal \N__29048\ : std_logic;
signal \N__29045\ : std_logic;
signal \N__29042\ : std_logic;
signal \N__29041\ : std_logic;
signal \N__29038\ : std_logic;
signal \N__29035\ : std_logic;
signal \N__29030\ : std_logic;
signal \N__29027\ : std_logic;
signal \N__29024\ : std_logic;
signal \N__29021\ : std_logic;
signal \N__29018\ : std_logic;
signal \N__29015\ : std_logic;
signal \N__29012\ : std_logic;
signal \N__29009\ : std_logic;
signal \N__29008\ : std_logic;
signal \N__29005\ : std_logic;
signal \N__29002\ : std_logic;
signal \N__28997\ : std_logic;
signal \N__28994\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28988\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28979\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28972\ : std_logic;
signal \N__28967\ : std_logic;
signal \N__28964\ : std_logic;
signal \N__28961\ : std_logic;
signal \N__28958\ : std_logic;
signal \N__28955\ : std_logic;
signal \N__28952\ : std_logic;
signal \N__28949\ : std_logic;
signal \N__28946\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28939\ : std_logic;
signal \N__28936\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28928\ : std_logic;
signal \N__28925\ : std_logic;
signal \N__28922\ : std_logic;
signal \N__28919\ : std_logic;
signal \N__28916\ : std_logic;
signal \N__28915\ : std_logic;
signal \N__28912\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28906\ : std_logic;
signal \N__28903\ : std_logic;
signal \N__28900\ : std_logic;
signal \N__28895\ : std_logic;
signal \N__28892\ : std_logic;
signal \N__28889\ : std_logic;
signal \N__28886\ : std_logic;
signal \N__28885\ : std_logic;
signal \N__28882\ : std_logic;
signal \N__28879\ : std_logic;
signal \N__28876\ : std_logic;
signal \N__28873\ : std_logic;
signal \N__28870\ : std_logic;
signal \N__28865\ : std_logic;
signal \N__28862\ : std_logic;
signal \N__28859\ : std_logic;
signal \N__28856\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28854\ : std_logic;
signal \N__28853\ : std_logic;
signal \N__28852\ : std_logic;
signal \N__28851\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28849\ : std_logic;
signal \N__28848\ : std_logic;
signal \N__28847\ : std_logic;
signal \N__28846\ : std_logic;
signal \N__28845\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28843\ : std_logic;
signal \N__28842\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28840\ : std_logic;
signal \N__28839\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28837\ : std_logic;
signal \N__28836\ : std_logic;
signal \N__28835\ : std_logic;
signal \N__28834\ : std_logic;
signal \N__28833\ : std_logic;
signal \N__28832\ : std_logic;
signal \N__28831\ : std_logic;
signal \N__28830\ : std_logic;
signal \N__28829\ : std_logic;
signal \N__28828\ : std_logic;
signal \N__28827\ : std_logic;
signal \N__28824\ : std_logic;
signal \N__28823\ : std_logic;
signal \N__28822\ : std_logic;
signal \N__28821\ : std_logic;
signal \N__28820\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28818\ : std_logic;
signal \N__28817\ : std_logic;
signal \N__28810\ : std_logic;
signal \N__28801\ : std_logic;
signal \N__28800\ : std_logic;
signal \N__28797\ : std_logic;
signal \N__28796\ : std_logic;
signal \N__28793\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28786\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28780\ : std_logic;
signal \N__28777\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28771\ : std_logic;
signal \N__28768\ : std_logic;
signal \N__28765\ : std_logic;
signal \N__28762\ : std_logic;
signal \N__28759\ : std_logic;
signal \N__28756\ : std_logic;
signal \N__28753\ : std_logic;
signal \N__28750\ : std_logic;
signal \N__28747\ : std_logic;
signal \N__28744\ : std_logic;
signal \N__28741\ : std_logic;
signal \N__28738\ : std_logic;
signal \N__28735\ : std_logic;
signal \N__28732\ : std_logic;
signal \N__28731\ : std_logic;
signal \N__28728\ : std_logic;
signal \N__28721\ : std_logic;
signal \N__28712\ : std_logic;
signal \N__28707\ : std_logic;
signal \N__28700\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28698\ : std_logic;
signal \N__28697\ : std_logic;
signal \N__28696\ : std_logic;
signal \N__28695\ : std_logic;
signal \N__28694\ : std_logic;
signal \N__28693\ : std_logic;
signal \N__28682\ : std_logic;
signal \N__28675\ : std_logic;
signal \N__28666\ : std_logic;
signal \N__28657\ : std_logic;
signal \N__28656\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28642\ : std_logic;
signal \N__28639\ : std_logic;
signal \N__28632\ : std_logic;
signal \N__28627\ : std_logic;
signal \N__28624\ : std_logic;
signal \N__28621\ : std_logic;
signal \N__28618\ : std_logic;
signal \N__28615\ : std_logic;
signal \N__28612\ : std_logic;
signal \N__28609\ : std_logic;
signal \N__28606\ : std_logic;
signal \N__28603\ : std_logic;
signal \N__28600\ : std_logic;
signal \N__28595\ : std_logic;
signal \N__28592\ : std_logic;
signal \N__28587\ : std_logic;
signal \N__28582\ : std_logic;
signal \N__28579\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28558\ : std_logic;
signal \N__28555\ : std_logic;
signal \N__28552\ : std_logic;
signal \N__28549\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28547\ : std_logic;
signal \N__28544\ : std_logic;
signal \N__28537\ : std_logic;
signal \N__28532\ : std_logic;
signal \N__28529\ : std_logic;
signal \N__28528\ : std_logic;
signal \N__28525\ : std_logic;
signal \N__28522\ : std_logic;
signal \N__28519\ : std_logic;
signal \N__28516\ : std_logic;
signal \N__28513\ : std_logic;
signal \N__28510\ : std_logic;
signal \N__28507\ : std_logic;
signal \N__28504\ : std_logic;
signal \N__28501\ : std_logic;
signal \N__28496\ : std_logic;
signal \N__28493\ : std_logic;
signal \N__28486\ : std_logic;
signal \N__28483\ : std_logic;
signal \N__28478\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28466\ : std_logic;
signal \N__28463\ : std_logic;
signal \N__28460\ : std_logic;
signal \N__28457\ : std_logic;
signal \N__28454\ : std_logic;
signal \N__28451\ : std_logic;
signal \N__28448\ : std_logic;
signal \N__28445\ : std_logic;
signal \N__28442\ : std_logic;
signal \N__28439\ : std_logic;
signal \N__28436\ : std_logic;
signal \N__28433\ : std_logic;
signal \N__28430\ : std_logic;
signal \N__28427\ : std_logic;
signal \N__28424\ : std_logic;
signal \N__28421\ : std_logic;
signal \N__28418\ : std_logic;
signal \N__28415\ : std_logic;
signal \N__28412\ : std_logic;
signal \N__28409\ : std_logic;
signal \N__28406\ : std_logic;
signal \N__28403\ : std_logic;
signal \N__28400\ : std_logic;
signal \N__28397\ : std_logic;
signal \N__28394\ : std_logic;
signal \N__28391\ : std_logic;
signal \N__28388\ : std_logic;
signal \N__28387\ : std_logic;
signal \N__28384\ : std_logic;
signal \N__28381\ : std_logic;
signal \N__28378\ : std_logic;
signal \N__28377\ : std_logic;
signal \N__28374\ : std_logic;
signal \N__28371\ : std_logic;
signal \N__28368\ : std_logic;
signal \N__28361\ : std_logic;
signal \N__28358\ : std_logic;
signal \N__28355\ : std_logic;
signal \N__28354\ : std_logic;
signal \N__28351\ : std_logic;
signal \N__28348\ : std_logic;
signal \N__28343\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28334\ : std_logic;
signal \N__28331\ : std_logic;
signal \N__28328\ : std_logic;
signal \N__28325\ : std_logic;
signal \N__28322\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28316\ : std_logic;
signal \N__28313\ : std_logic;
signal \N__28312\ : std_logic;
signal \N__28309\ : std_logic;
signal \N__28306\ : std_logic;
signal \N__28301\ : std_logic;
signal \N__28298\ : std_logic;
signal \N__28295\ : std_logic;
signal \N__28292\ : std_logic;
signal \N__28289\ : std_logic;
signal \N__28286\ : std_logic;
signal \N__28283\ : std_logic;
signal \N__28280\ : std_logic;
signal \N__28279\ : std_logic;
signal \N__28276\ : std_logic;
signal \N__28273\ : std_logic;
signal \N__28268\ : std_logic;
signal \N__28265\ : std_logic;
signal \N__28262\ : std_logic;
signal \N__28259\ : std_logic;
signal \N__28256\ : std_logic;
signal \N__28253\ : std_logic;
signal \N__28250\ : std_logic;
signal \N__28249\ : std_logic;
signal \N__28248\ : std_logic;
signal \N__28247\ : std_logic;
signal \N__28240\ : std_logic;
signal \N__28237\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28231\ : std_logic;
signal \N__28226\ : std_logic;
signal \N__28223\ : std_logic;
signal \N__28220\ : std_logic;
signal \N__28217\ : std_logic;
signal \N__28214\ : std_logic;
signal \N__28211\ : std_logic;
signal \N__28208\ : std_logic;
signal \N__28205\ : std_logic;
signal \N__28202\ : std_logic;
signal \N__28199\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28193\ : std_logic;
signal \N__28190\ : std_logic;
signal \N__28187\ : std_logic;
signal \N__28184\ : std_logic;
signal \N__28181\ : std_logic;
signal \N__28178\ : std_logic;
signal \N__28175\ : std_logic;
signal \N__28172\ : std_logic;
signal \N__28169\ : std_logic;
signal \N__28166\ : std_logic;
signal \N__28163\ : std_logic;
signal \N__28160\ : std_logic;
signal \N__28157\ : std_logic;
signal \N__28154\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28144\ : std_logic;
signal \N__28141\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28139\ : std_logic;
signal \N__28136\ : std_logic;
signal \N__28131\ : std_logic;
signal \N__28128\ : std_logic;
signal \N__28123\ : std_logic;
signal \N__28120\ : std_logic;
signal \N__28115\ : std_logic;
signal \N__28112\ : std_logic;
signal \N__28109\ : std_logic;
signal \N__28106\ : std_logic;
signal \N__28103\ : std_logic;
signal \N__28100\ : std_logic;
signal \N__28097\ : std_logic;
signal \N__28094\ : std_logic;
signal \N__28091\ : std_logic;
signal \N__28088\ : std_logic;
signal \N__28085\ : std_logic;
signal \N__28082\ : std_logic;
signal \N__28079\ : std_logic;
signal \N__28076\ : std_logic;
signal \N__28073\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28067\ : std_logic;
signal \N__28064\ : std_logic;
signal \N__28061\ : std_logic;
signal \N__28058\ : std_logic;
signal \N__28055\ : std_logic;
signal \N__28052\ : std_logic;
signal \N__28049\ : std_logic;
signal \N__28046\ : std_logic;
signal \N__28043\ : std_logic;
signal \N__28040\ : std_logic;
signal \N__28037\ : std_logic;
signal \N__28034\ : std_logic;
signal \N__28031\ : std_logic;
signal \N__28028\ : std_logic;
signal \N__28025\ : std_logic;
signal \N__28022\ : std_logic;
signal \N__28019\ : std_logic;
signal \N__28016\ : std_logic;
signal \N__28013\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27997\ : std_logic;
signal \N__27994\ : std_logic;
signal \N__27993\ : std_logic;
signal \N__27992\ : std_logic;
signal \N__27989\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27976\ : std_logic;
signal \N__27973\ : std_logic;
signal \N__27968\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27959\ : std_logic;
signal \N__27956\ : std_logic;
signal \N__27953\ : std_logic;
signal \N__27950\ : std_logic;
signal \N__27949\ : std_logic;
signal \N__27948\ : std_logic;
signal \N__27945\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27939\ : std_logic;
signal \N__27934\ : std_logic;
signal \N__27931\ : std_logic;
signal \N__27928\ : std_logic;
signal \N__27925\ : std_logic;
signal \N__27920\ : std_logic;
signal \N__27917\ : std_logic;
signal \N__27914\ : std_logic;
signal \N__27911\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27905\ : std_logic;
signal \N__27902\ : std_logic;
signal \N__27899\ : std_logic;
signal \N__27896\ : std_logic;
signal \N__27893\ : std_logic;
signal \N__27890\ : std_logic;
signal \N__27887\ : std_logic;
signal \N__27884\ : std_logic;
signal \N__27881\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27875\ : std_logic;
signal \N__27872\ : std_logic;
signal \N__27869\ : std_logic;
signal \N__27866\ : std_logic;
signal \N__27863\ : std_logic;
signal \N__27860\ : std_logic;
signal \N__27857\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27853\ : std_logic;
signal \N__27852\ : std_logic;
signal \N__27849\ : std_logic;
signal \N__27846\ : std_logic;
signal \N__27843\ : std_logic;
signal \N__27842\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27829\ : std_logic;
signal \N__27826\ : std_logic;
signal \N__27821\ : std_logic;
signal \N__27818\ : std_logic;
signal \N__27815\ : std_logic;
signal \N__27812\ : std_logic;
signal \N__27809\ : std_logic;
signal \N__27806\ : std_logic;
signal \N__27803\ : std_logic;
signal \N__27800\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27798\ : std_logic;
signal \N__27797\ : std_logic;
signal \N__27794\ : std_logic;
signal \N__27789\ : std_logic;
signal \N__27786\ : std_logic;
signal \N__27783\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27773\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27764\ : std_logic;
signal \N__27761\ : std_logic;
signal \N__27758\ : std_logic;
signal \N__27757\ : std_logic;
signal \N__27756\ : std_logic;
signal \N__27753\ : std_logic;
signal \N__27752\ : std_logic;
signal \N__27749\ : std_logic;
signal \N__27746\ : std_logic;
signal \N__27741\ : std_logic;
signal \N__27738\ : std_logic;
signal \N__27735\ : std_logic;
signal \N__27732\ : std_logic;
signal \N__27729\ : std_logic;
signal \N__27722\ : std_logic;
signal \N__27719\ : std_logic;
signal \N__27716\ : std_logic;
signal \N__27713\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27701\ : std_logic;
signal \N__27698\ : std_logic;
signal \N__27695\ : std_logic;
signal \N__27692\ : std_logic;
signal \N__27689\ : std_logic;
signal \N__27686\ : std_logic;
signal \N__27683\ : std_logic;
signal \N__27680\ : std_logic;
signal \N__27677\ : std_logic;
signal \N__27676\ : std_logic;
signal \N__27675\ : std_logic;
signal \N__27674\ : std_logic;
signal \N__27669\ : std_logic;
signal \N__27666\ : std_logic;
signal \N__27663\ : std_logic;
signal \N__27660\ : std_logic;
signal \N__27655\ : std_logic;
signal \N__27650\ : std_logic;
signal \N__27647\ : std_logic;
signal \N__27644\ : std_logic;
signal \N__27641\ : std_logic;
signal \N__27638\ : std_logic;
signal \N__27635\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27626\ : std_logic;
signal \N__27623\ : std_logic;
signal \N__27620\ : std_logic;
signal \N__27617\ : std_logic;
signal \N__27614\ : std_logic;
signal \N__27611\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27598\ : std_logic;
signal \N__27597\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27595\ : std_logic;
signal \N__27592\ : std_logic;
signal \N__27591\ : std_logic;
signal \N__27582\ : std_logic;
signal \N__27579\ : std_logic;
signal \N__27576\ : std_logic;
signal \N__27569\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27565\ : std_logic;
signal \N__27564\ : std_logic;
signal \N__27563\ : std_logic;
signal \N__27560\ : std_logic;
signal \N__27555\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27533\ : std_logic;
signal \N__27530\ : std_logic;
signal \N__27527\ : std_logic;
signal \N__27526\ : std_logic;
signal \N__27521\ : std_logic;
signal \N__27520\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27509\ : std_logic;
signal \N__27506\ : std_logic;
signal \N__27503\ : std_logic;
signal \N__27500\ : std_logic;
signal \N__27497\ : std_logic;
signal \N__27494\ : std_logic;
signal \N__27491\ : std_logic;
signal \N__27488\ : std_logic;
signal \N__27487\ : std_logic;
signal \N__27486\ : std_logic;
signal \N__27485\ : std_logic;
signal \N__27480\ : std_logic;
signal \N__27477\ : std_logic;
signal \N__27474\ : std_logic;
signal \N__27469\ : std_logic;
signal \N__27466\ : std_logic;
signal \N__27461\ : std_logic;
signal \N__27458\ : std_logic;
signal \N__27455\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27446\ : std_logic;
signal \N__27443\ : std_logic;
signal \N__27440\ : std_logic;
signal \N__27437\ : std_logic;
signal \N__27434\ : std_logic;
signal \N__27431\ : std_logic;
signal \N__27428\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27419\ : std_logic;
signal \N__27416\ : std_logic;
signal \N__27413\ : std_logic;
signal \N__27410\ : std_logic;
signal \N__27407\ : std_logic;
signal \N__27404\ : std_logic;
signal \N__27401\ : std_logic;
signal \N__27398\ : std_logic;
signal \N__27397\ : std_logic;
signal \N__27394\ : std_logic;
signal \N__27393\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27389\ : std_logic;
signal \N__27386\ : std_logic;
signal \N__27383\ : std_logic;
signal \N__27380\ : std_logic;
signal \N__27377\ : std_logic;
signal \N__27368\ : std_logic;
signal \N__27365\ : std_logic;
signal \N__27362\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27356\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27350\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27346\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27339\ : std_logic;
signal \N__27336\ : std_logic;
signal \N__27329\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27325\ : std_logic;
signal \N__27324\ : std_logic;
signal \N__27321\ : std_logic;
signal \N__27318\ : std_logic;
signal \N__27315\ : std_logic;
signal \N__27308\ : std_logic;
signal \N__27305\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27303\ : std_logic;
signal \N__27300\ : std_logic;
signal \N__27297\ : std_logic;
signal \N__27294\ : std_logic;
signal \N__27291\ : std_logic;
signal \N__27284\ : std_logic;
signal \N__27281\ : std_logic;
signal \N__27280\ : std_logic;
signal \N__27279\ : std_logic;
signal \N__27278\ : std_logic;
signal \N__27277\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27275\ : std_logic;
signal \N__27274\ : std_logic;
signal \N__27273\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27269\ : std_logic;
signal \N__27266\ : std_logic;
signal \N__27257\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27242\ : std_logic;
signal \N__27233\ : std_logic;
signal \N__27230\ : std_logic;
signal \N__27229\ : std_logic;
signal \N__27228\ : std_logic;
signal \N__27225\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27219\ : std_logic;
signal \N__27216\ : std_logic;
signal \N__27209\ : std_logic;
signal \N__27206\ : std_logic;
signal \N__27203\ : std_logic;
signal \N__27200\ : std_logic;
signal \N__27197\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27195\ : std_logic;
signal \N__27192\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27186\ : std_logic;
signal \N__27179\ : std_logic;
signal \N__27176\ : std_logic;
signal \N__27175\ : std_logic;
signal \N__27174\ : std_logic;
signal \N__27171\ : std_logic;
signal \N__27168\ : std_logic;
signal \N__27165\ : std_logic;
signal \N__27158\ : std_logic;
signal \N__27155\ : std_logic;
signal \N__27154\ : std_logic;
signal \N__27153\ : std_logic;
signal \N__27150\ : std_logic;
signal \N__27147\ : std_logic;
signal \N__27144\ : std_logic;
signal \N__27137\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27133\ : std_logic;
signal \N__27132\ : std_logic;
signal \N__27129\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27112\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27108\ : std_logic;
signal \N__27105\ : std_logic;
signal \N__27102\ : std_logic;
signal \N__27095\ : std_logic;
signal \N__27092\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27090\ : std_logic;
signal \N__27087\ : std_logic;
signal \N__27084\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27071\ : std_logic;
signal \N__27070\ : std_logic;
signal \N__27067\ : std_logic;
signal \N__27064\ : std_logic;
signal \N__27063\ : std_logic;
signal \N__27058\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27052\ : std_logic;
signal \N__27047\ : std_logic;
signal \N__27044\ : std_logic;
signal \N__27043\ : std_logic;
signal \N__27040\ : std_logic;
signal \N__27037\ : std_logic;
signal \N__27036\ : std_logic;
signal \N__27031\ : std_logic;
signal \N__27028\ : std_logic;
signal \N__27025\ : std_logic;
signal \N__27020\ : std_logic;
signal \N__27017\ : std_logic;
signal \N__27016\ : std_logic;
signal \N__27013\ : std_logic;
signal \N__27010\ : std_logic;
signal \N__27005\ : std_logic;
signal \N__27004\ : std_logic;
signal \N__27001\ : std_logic;
signal \N__26998\ : std_logic;
signal \N__26995\ : std_logic;
signal \N__26990\ : std_logic;
signal \N__26987\ : std_logic;
signal \N__26986\ : std_logic;
signal \N__26983\ : std_logic;
signal \N__26980\ : std_logic;
signal \N__26979\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26968\ : std_logic;
signal \N__26963\ : std_logic;
signal \N__26960\ : std_logic;
signal \N__26957\ : std_logic;
signal \N__26956\ : std_logic;
signal \N__26953\ : std_logic;
signal \N__26950\ : std_logic;
signal \N__26947\ : std_logic;
signal \N__26942\ : std_logic;
signal \N__26939\ : std_logic;
signal \N__26936\ : std_logic;
signal \N__26935\ : std_logic;
signal \N__26932\ : std_logic;
signal \N__26929\ : std_logic;
signal \N__26926\ : std_logic;
signal \N__26921\ : std_logic;
signal \N__26918\ : std_logic;
signal \N__26915\ : std_logic;
signal \N__26914\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26908\ : std_logic;
signal \N__26907\ : std_logic;
signal \N__26902\ : std_logic;
signal \N__26899\ : std_logic;
signal \N__26896\ : std_logic;
signal \N__26891\ : std_logic;
signal \N__26888\ : std_logic;
signal \N__26887\ : std_logic;
signal \N__26884\ : std_logic;
signal \N__26881\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26875\ : std_logic;
signal \N__26872\ : std_logic;
signal \N__26869\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26861\ : std_logic;
signal \N__26860\ : std_logic;
signal \N__26857\ : std_logic;
signal \N__26854\ : std_logic;
signal \N__26849\ : std_logic;
signal \N__26848\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26834\ : std_logic;
signal \N__26831\ : std_logic;
signal \N__26830\ : std_logic;
signal \N__26827\ : std_logic;
signal \N__26824\ : std_logic;
signal \N__26819\ : std_logic;
signal \N__26818\ : std_logic;
signal \N__26815\ : std_logic;
signal \N__26812\ : std_logic;
signal \N__26809\ : std_logic;
signal \N__26804\ : std_logic;
signal \N__26801\ : std_logic;
signal \N__26800\ : std_logic;
signal \N__26795\ : std_logic;
signal \N__26794\ : std_logic;
signal \N__26791\ : std_logic;
signal \N__26788\ : std_logic;
signal \N__26785\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26776\ : std_logic;
signal \N__26771\ : std_logic;
signal \N__26770\ : std_logic;
signal \N__26767\ : std_logic;
signal \N__26764\ : std_logic;
signal \N__26761\ : std_logic;
signal \N__26756\ : std_logic;
signal \N__26753\ : std_logic;
signal \N__26752\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26746\ : std_logic;
signal \N__26741\ : std_logic;
signal \N__26740\ : std_logic;
signal \N__26737\ : std_logic;
signal \N__26734\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26726\ : std_logic;
signal \N__26723\ : std_logic;
signal \N__26722\ : std_logic;
signal \N__26719\ : std_logic;
signal \N__26716\ : std_logic;
signal \N__26715\ : std_logic;
signal \N__26710\ : std_logic;
signal \N__26707\ : std_logic;
signal \N__26704\ : std_logic;
signal \N__26699\ : std_logic;
signal \N__26696\ : std_logic;
signal \N__26695\ : std_logic;
signal \N__26692\ : std_logic;
signal \N__26689\ : std_logic;
signal \N__26686\ : std_logic;
signal \N__26685\ : std_logic;
signal \N__26680\ : std_logic;
signal \N__26677\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26669\ : std_logic;
signal \N__26666\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26662\ : std_logic;
signal \N__26659\ : std_logic;
signal \N__26658\ : std_logic;
signal \N__26653\ : std_logic;
signal \N__26650\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26642\ : std_logic;
signal \N__26639\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26635\ : std_logic;
signal \N__26632\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26626\ : std_logic;
signal \N__26623\ : std_logic;
signal \N__26620\ : std_logic;
signal \N__26617\ : std_logic;
signal \N__26612\ : std_logic;
signal \N__26609\ : std_logic;
signal \N__26608\ : std_logic;
signal \N__26605\ : std_logic;
signal \N__26602\ : std_logic;
signal \N__26601\ : std_logic;
signal \N__26596\ : std_logic;
signal \N__26593\ : std_logic;
signal \N__26590\ : std_logic;
signal \N__26585\ : std_logic;
signal \N__26582\ : std_logic;
signal \N__26581\ : std_logic;
signal \N__26580\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26572\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26560\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26554\ : std_logic;
signal \N__26551\ : std_logic;
signal \N__26548\ : std_logic;
signal \N__26545\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26533\ : std_logic;
signal \N__26530\ : std_logic;
signal \N__26529\ : std_logic;
signal \N__26524\ : std_logic;
signal \N__26521\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26513\ : std_logic;
signal \N__26510\ : std_logic;
signal \N__26509\ : std_logic;
signal \N__26506\ : std_logic;
signal \N__26503\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26497\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26488\ : std_logic;
signal \N__26483\ : std_logic;
signal \N__26480\ : std_logic;
signal \N__26477\ : std_logic;
signal \N__26476\ : std_logic;
signal \N__26475\ : std_logic;
signal \N__26474\ : std_logic;
signal \N__26473\ : std_logic;
signal \N__26462\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26452\ : std_logic;
signal \N__26449\ : std_logic;
signal \N__26446\ : std_logic;
signal \N__26443\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26439\ : std_logic;
signal \N__26436\ : std_logic;
signal \N__26433\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26423\ : std_logic;
signal \N__26422\ : std_logic;
signal \N__26419\ : std_logic;
signal \N__26416\ : std_logic;
signal \N__26415\ : std_logic;
signal \N__26410\ : std_logic;
signal \N__26407\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26398\ : std_logic;
signal \N__26395\ : std_logic;
signal \N__26392\ : std_logic;
signal \N__26391\ : std_logic;
signal \N__26386\ : std_logic;
signal \N__26383\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26371\ : std_logic;
signal \N__26368\ : std_logic;
signal \N__26365\ : std_logic;
signal \N__26360\ : std_logic;
signal \N__26359\ : std_logic;
signal \N__26356\ : std_logic;
signal \N__26353\ : std_logic;
signal \N__26350\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26342\ : std_logic;
signal \N__26341\ : std_logic;
signal \N__26340\ : std_logic;
signal \N__26335\ : std_logic;
signal \N__26332\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26324\ : std_logic;
signal \N__26321\ : std_logic;
signal \N__26320\ : std_logic;
signal \N__26315\ : std_logic;
signal \N__26314\ : std_logic;
signal \N__26311\ : std_logic;
signal \N__26308\ : std_logic;
signal \N__26305\ : std_logic;
signal \N__26300\ : std_logic;
signal \N__26297\ : std_logic;
signal \N__26296\ : std_logic;
signal \N__26293\ : std_logic;
signal \N__26290\ : std_logic;
signal \N__26287\ : std_logic;
signal \N__26286\ : std_logic;
signal \N__26283\ : std_logic;
signal \N__26280\ : std_logic;
signal \N__26277\ : std_logic;
signal \N__26272\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26263\ : std_logic;
signal \N__26260\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26256\ : std_logic;
signal \N__26251\ : std_logic;
signal \N__26248\ : std_logic;
signal \N__26245\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26237\ : std_logic;
signal \N__26234\ : std_logic;
signal \N__26231\ : std_logic;
signal \N__26228\ : std_logic;
signal \N__26225\ : std_logic;
signal \N__26222\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26216\ : std_logic;
signal \N__26213\ : std_logic;
signal \N__26210\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26198\ : std_logic;
signal \N__26195\ : std_logic;
signal \N__26192\ : std_logic;
signal \N__26189\ : std_logic;
signal \N__26186\ : std_logic;
signal \N__26183\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26177\ : std_logic;
signal \N__26174\ : std_logic;
signal \N__26171\ : std_logic;
signal \N__26168\ : std_logic;
signal \N__26165\ : std_logic;
signal \N__26162\ : std_logic;
signal \N__26159\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26150\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26144\ : std_logic;
signal \N__26141\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26135\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26129\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26123\ : std_logic;
signal \N__26120\ : std_logic;
signal \N__26117\ : std_logic;
signal \N__26114\ : std_logic;
signal \N__26111\ : std_logic;
signal \N__26108\ : std_logic;
signal \N__26105\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26096\ : std_logic;
signal \N__26093\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26084\ : std_logic;
signal \N__26081\ : std_logic;
signal \N__26078\ : std_logic;
signal \N__26075\ : std_logic;
signal \N__26072\ : std_logic;
signal \N__26069\ : std_logic;
signal \N__26066\ : std_logic;
signal \N__26063\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26054\ : std_logic;
signal \N__26051\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26033\ : std_logic;
signal \N__26030\ : std_logic;
signal \N__26027\ : std_logic;
signal \N__26024\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26015\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26006\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__26000\ : std_logic;
signal \N__25997\ : std_logic;
signal \N__25994\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25985\ : std_logic;
signal \N__25982\ : std_logic;
signal \N__25979\ : std_logic;
signal \N__25976\ : std_logic;
signal \N__25973\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25967\ : std_logic;
signal \N__25964\ : std_logic;
signal \N__25961\ : std_logic;
signal \N__25958\ : std_logic;
signal \N__25955\ : std_logic;
signal \N__25954\ : std_logic;
signal \N__25951\ : std_logic;
signal \N__25950\ : std_logic;
signal \N__25947\ : std_logic;
signal \N__25946\ : std_logic;
signal \N__25943\ : std_logic;
signal \N__25940\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25927\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25919\ : std_logic;
signal \N__25916\ : std_logic;
signal \N__25913\ : std_logic;
signal \N__25910\ : std_logic;
signal \N__25907\ : std_logic;
signal \N__25906\ : std_logic;
signal \N__25905\ : std_logic;
signal \N__25902\ : std_logic;
signal \N__25899\ : std_logic;
signal \N__25896\ : std_logic;
signal \N__25893\ : std_logic;
signal \N__25890\ : std_logic;
signal \N__25887\ : std_logic;
signal \N__25886\ : std_logic;
signal \N__25883\ : std_logic;
signal \N__25878\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25872\ : std_logic;
signal \N__25865\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25859\ : std_logic;
signal \N__25856\ : std_logic;
signal \N__25853\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25849\ : std_logic;
signal \N__25848\ : std_logic;
signal \N__25847\ : std_logic;
signal \N__25844\ : std_logic;
signal \N__25841\ : std_logic;
signal \N__25838\ : std_logic;
signal \N__25835\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25829\ : std_logic;
signal \N__25826\ : std_logic;
signal \N__25823\ : std_logic;
signal \N__25820\ : std_logic;
signal \N__25817\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25805\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25795\ : std_logic;
signal \N__25792\ : std_logic;
signal \N__25791\ : std_logic;
signal \N__25788\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25781\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25772\ : std_logic;
signal \N__25769\ : std_logic;
signal \N__25766\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25760\ : std_logic;
signal \N__25755\ : std_logic;
signal \N__25752\ : std_logic;
signal \N__25745\ : std_logic;
signal \N__25742\ : std_logic;
signal \N__25739\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25733\ : std_logic;
signal \N__25732\ : std_logic;
signal \N__25731\ : std_logic;
signal \N__25730\ : std_logic;
signal \N__25729\ : std_logic;
signal \N__25728\ : std_logic;
signal \N__25725\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25720\ : std_logic;
signal \N__25717\ : std_logic;
signal \N__25714\ : std_logic;
signal \N__25699\ : std_logic;
signal \N__25696\ : std_logic;
signal \N__25693\ : std_logic;
signal \N__25690\ : std_logic;
signal \N__25687\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25679\ : std_logic;
signal \N__25678\ : std_logic;
signal \N__25677\ : std_logic;
signal \N__25676\ : std_logic;
signal \N__25675\ : std_logic;
signal \N__25674\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25672\ : std_logic;
signal \N__25671\ : std_logic;
signal \N__25670\ : std_logic;
signal \N__25669\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25667\ : std_logic;
signal \N__25666\ : std_logic;
signal \N__25665\ : std_logic;
signal \N__25664\ : std_logic;
signal \N__25659\ : std_logic;
signal \N__25658\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25654\ : std_logic;
signal \N__25653\ : std_logic;
signal \N__25650\ : std_logic;
signal \N__25649\ : std_logic;
signal \N__25646\ : std_logic;
signal \N__25645\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25639\ : std_logic;
signal \N__25636\ : std_logic;
signal \N__25635\ : std_logic;
signal \N__25634\ : std_logic;
signal \N__25633\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25629\ : std_logic;
signal \N__25626\ : std_logic;
signal \N__25623\ : std_logic;
signal \N__25620\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25618\ : std_logic;
signal \N__25615\ : std_logic;
signal \N__25614\ : std_logic;
signal \N__25613\ : std_logic;
signal \N__25610\ : std_logic;
signal \N__25607\ : std_logic;
signal \N__25604\ : std_logic;
signal \N__25603\ : std_logic;
signal \N__25602\ : std_logic;
signal \N__25601\ : std_logic;
signal \N__25598\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25587\ : std_logic;
signal \N__25582\ : std_logic;
signal \N__25579\ : std_logic;
signal \N__25564\ : std_logic;
signal \N__25561\ : std_logic;
signal \N__25548\ : std_logic;
signal \N__25543\ : std_logic;
signal \N__25528\ : std_logic;
signal \N__25525\ : std_logic;
signal \N__25518\ : std_logic;
signal \N__25513\ : std_logic;
signal \N__25508\ : std_logic;
signal \N__25493\ : std_logic;
signal \N__25490\ : std_logic;
signal \N__25487\ : std_logic;
signal \N__25484\ : std_logic;
signal \N__25481\ : std_logic;
signal \N__25478\ : std_logic;
signal \N__25475\ : std_logic;
signal \N__25472\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25466\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25462\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25457\ : std_logic;
signal \N__25454\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25442\ : std_logic;
signal \N__25441\ : std_logic;
signal \N__25438\ : std_logic;
signal \N__25435\ : std_logic;
signal \N__25432\ : std_logic;
signal \N__25429\ : std_logic;
signal \N__25426\ : std_logic;
signal \N__25423\ : std_logic;
signal \N__25420\ : std_logic;
signal \N__25417\ : std_logic;
signal \N__25412\ : std_logic;
signal \N__25409\ : std_logic;
signal \N__25406\ : std_logic;
signal \N__25403\ : std_logic;
signal \N__25400\ : std_logic;
signal \N__25397\ : std_logic;
signal \N__25396\ : std_logic;
signal \N__25393\ : std_logic;
signal \N__25390\ : std_logic;
signal \N__25387\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25376\ : std_logic;
signal \N__25373\ : std_logic;
signal \N__25370\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25360\ : std_logic;
signal \N__25357\ : std_logic;
signal \N__25354\ : std_logic;
signal \N__25351\ : std_logic;
signal \N__25348\ : std_logic;
signal \N__25345\ : std_logic;
signal \N__25342\ : std_logic;
signal \N__25339\ : std_logic;
signal \N__25336\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25321\ : std_logic;
signal \N__25320\ : std_logic;
signal \N__25317\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25304\ : std_logic;
signal \N__25299\ : std_logic;
signal \N__25292\ : std_logic;
signal \N__25289\ : std_logic;
signal \N__25288\ : std_logic;
signal \N__25285\ : std_logic;
signal \N__25282\ : std_logic;
signal \N__25279\ : std_logic;
signal \N__25274\ : std_logic;
signal \N__25271\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25265\ : std_logic;
signal \N__25262\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25258\ : std_logic;
signal \N__25257\ : std_logic;
signal \N__25254\ : std_logic;
signal \N__25251\ : std_logic;
signal \N__25250\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25244\ : std_logic;
signal \N__25241\ : std_logic;
signal \N__25238\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25226\ : std_logic;
signal \N__25223\ : std_logic;
signal \N__25222\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25216\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25193\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25184\ : std_logic;
signal \N__25181\ : std_logic;
signal \N__25180\ : std_logic;
signal \N__25177\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25173\ : std_logic;
signal \N__25170\ : std_logic;
signal \N__25167\ : std_logic;
signal \N__25166\ : std_logic;
signal \N__25163\ : std_logic;
signal \N__25158\ : std_logic;
signal \N__25155\ : std_logic;
signal \N__25152\ : std_logic;
signal \N__25145\ : std_logic;
signal \N__25144\ : std_logic;
signal \N__25141\ : std_logic;
signal \N__25138\ : std_logic;
signal \N__25135\ : std_logic;
signal \N__25132\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25123\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25115\ : std_logic;
signal \N__25112\ : std_logic;
signal \N__25109\ : std_logic;
signal \N__25106\ : std_logic;
signal \N__25105\ : std_logic;
signal \N__25102\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25098\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25092\ : std_logic;
signal \N__25091\ : std_logic;
signal \N__25088\ : std_logic;
signal \N__25083\ : std_logic;
signal \N__25080\ : std_logic;
signal \N__25077\ : std_logic;
signal \N__25070\ : std_logic;
signal \N__25067\ : std_logic;
signal \N__25064\ : std_logic;
signal \N__25061\ : std_logic;
signal \N__25058\ : std_logic;
signal \N__25055\ : std_logic;
signal \N__25054\ : std_logic;
signal \N__25051\ : std_logic;
signal \N__25050\ : std_logic;
signal \N__25047\ : std_logic;
signal \N__25044\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25040\ : std_logic;
signal \N__25037\ : std_logic;
signal \N__25034\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25028\ : std_logic;
signal \N__25025\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25014\ : std_logic;
signal \N__25007\ : std_logic;
signal \N__25004\ : std_logic;
signal \N__25001\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24982\ : std_logic;
signal \N__24979\ : std_logic;
signal \N__24976\ : std_logic;
signal \N__24973\ : std_logic;
signal \N__24972\ : std_logic;
signal \N__24971\ : std_logic;
signal \N__24968\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24962\ : std_logic;
signal \N__24959\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24947\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24940\ : std_logic;
signal \N__24937\ : std_logic;
signal \N__24934\ : std_logic;
signal \N__24931\ : std_logic;
signal \N__24926\ : std_logic;
signal \N__24923\ : std_logic;
signal \N__24920\ : std_logic;
signal \N__24917\ : std_logic;
signal \N__24914\ : std_logic;
signal \N__24911\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24907\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24898\ : std_logic;
signal \N__24895\ : std_logic;
signal \N__24892\ : std_logic;
signal \N__24887\ : std_logic;
signal \N__24884\ : std_logic;
signal \N__24881\ : std_logic;
signal \N__24880\ : std_logic;
signal \N__24879\ : std_logic;
signal \N__24876\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24869\ : std_logic;
signal \N__24866\ : std_logic;
signal \N__24863\ : std_logic;
signal \N__24860\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24852\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24842\ : std_logic;
signal \N__24839\ : std_logic;
signal \N__24836\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24832\ : std_logic;
signal \N__24829\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24822\ : std_logic;
signal \N__24821\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24796\ : std_logic;
signal \N__24793\ : std_logic;
signal \N__24790\ : std_logic;
signal \N__24787\ : std_logic;
signal \N__24784\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24773\ : std_logic;
signal \N__24770\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24761\ : std_logic;
signal \N__24758\ : std_logic;
signal \N__24755\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24753\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24747\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24734\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24728\ : std_logic;
signal \N__24719\ : std_logic;
signal \N__24718\ : std_logic;
signal \N__24715\ : std_logic;
signal \N__24712\ : std_logic;
signal \N__24709\ : std_logic;
signal \N__24706\ : std_logic;
signal \N__24703\ : std_logic;
signal \N__24700\ : std_logic;
signal \N__24697\ : std_logic;
signal \N__24692\ : std_logic;
signal \N__24689\ : std_logic;
signal \N__24686\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24679\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24666\ : std_logic;
signal \N__24659\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24655\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24646\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24640\ : std_logic;
signal \N__24637\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24629\ : std_logic;
signal \N__24626\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24620\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24613\ : std_logic;
signal \N__24612\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24610\ : std_logic;
signal \N__24607\ : std_logic;
signal \N__24600\ : std_logic;
signal \N__24599\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24593\ : std_logic;
signal \N__24590\ : std_logic;
signal \N__24587\ : std_logic;
signal \N__24578\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24571\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24565\ : std_logic;
signal \N__24562\ : std_logic;
signal \N__24559\ : std_logic;
signal \N__24556\ : std_logic;
signal \N__24551\ : std_logic;
signal \N__24548\ : std_logic;
signal \N__24545\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24539\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24535\ : std_logic;
signal \N__24534\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24522\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24511\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24505\ : std_logic;
signal \N__24502\ : std_logic;
signal \N__24499\ : std_logic;
signal \N__24496\ : std_logic;
signal \N__24493\ : std_logic;
signal \N__24490\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24482\ : std_logic;
signal \N__24479\ : std_logic;
signal \N__24476\ : std_logic;
signal \N__24473\ : std_logic;
signal \N__24472\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24465\ : std_logic;
signal \N__24460\ : std_logic;
signal \N__24459\ : std_logic;
signal \N__24456\ : std_logic;
signal \N__24453\ : std_logic;
signal \N__24448\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24442\ : std_logic;
signal \N__24439\ : std_logic;
signal \N__24436\ : std_logic;
signal \N__24433\ : std_logic;
signal \N__24430\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24424\ : std_logic;
signal \N__24421\ : std_logic;
signal \N__24418\ : std_logic;
signal \N__24413\ : std_logic;
signal \N__24410\ : std_logic;
signal \N__24407\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24395\ : std_logic;
signal \N__24394\ : std_logic;
signal \N__24391\ : std_logic;
signal \N__24388\ : std_logic;
signal \N__24387\ : std_logic;
signal \N__24386\ : std_logic;
signal \N__24381\ : std_logic;
signal \N__24376\ : std_logic;
signal \N__24373\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24365\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24355\ : std_logic;
signal \N__24352\ : std_logic;
signal \N__24349\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24341\ : std_logic;
signal \N__24338\ : std_logic;
signal \N__24335\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24316\ : std_logic;
signal \N__24313\ : std_logic;
signal \N__24310\ : std_logic;
signal \N__24307\ : std_logic;
signal \N__24302\ : std_logic;
signal \N__24299\ : std_logic;
signal \N__24298\ : std_logic;
signal \N__24295\ : std_logic;
signal \N__24292\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24290\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24284\ : std_logic;
signal \N__24279\ : std_logic;
signal \N__24272\ : std_logic;
signal \N__24269\ : std_logic;
signal \N__24266\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24260\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24256\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24248\ : std_logic;
signal \N__24243\ : std_logic;
signal \N__24236\ : std_logic;
signal \N__24235\ : std_logic;
signal \N__24232\ : std_logic;
signal \N__24229\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24217\ : std_logic;
signal \N__24214\ : std_logic;
signal \N__24211\ : std_logic;
signal \N__24206\ : std_logic;
signal \N__24203\ : std_logic;
signal \N__24200\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24190\ : std_logic;
signal \N__24189\ : std_logic;
signal \N__24188\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24180\ : std_logic;
signal \N__24177\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24169\ : std_logic;
signal \N__24166\ : std_logic;
signal \N__24163\ : std_logic;
signal \N__24160\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24154\ : std_logic;
signal \N__24151\ : std_logic;
signal \N__24148\ : std_logic;
signal \N__24145\ : std_logic;
signal \N__24140\ : std_logic;
signal \N__24137\ : std_logic;
signal \N__24134\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24128\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24126\ : std_logic;
signal \N__24123\ : std_logic;
signal \N__24120\ : std_logic;
signal \N__24119\ : std_logic;
signal \N__24116\ : std_logic;
signal \N__24111\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24097\ : std_logic;
signal \N__24094\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24088\ : std_logic;
signal \N__24085\ : std_logic;
signal \N__24080\ : std_logic;
signal \N__24077\ : std_logic;
signal \N__24074\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24065\ : std_logic;
signal \N__24064\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24060\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24050\ : std_logic;
signal \N__24047\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24039\ : std_logic;
signal \N__24032\ : std_logic;
signal \N__24031\ : std_logic;
signal \N__24028\ : std_logic;
signal \N__24025\ : std_logic;
signal \N__24022\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24016\ : std_logic;
signal \N__24013\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24007\ : std_logic;
signal \N__24002\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23996\ : std_logic;
signal \N__23993\ : std_logic;
signal \N__23990\ : std_logic;
signal \N__23989\ : std_logic;
signal \N__23988\ : std_logic;
signal \N__23985\ : std_logic;
signal \N__23982\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23975\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23964\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23953\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23947\ : std_logic;
signal \N__23944\ : std_logic;
signal \N__23941\ : std_logic;
signal \N__23938\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23930\ : std_logic;
signal \N__23927\ : std_logic;
signal \N__23924\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23918\ : std_logic;
signal \N__23915\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23911\ : std_logic;
signal \N__23908\ : std_logic;
signal \N__23905\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23899\ : std_logic;
signal \N__23896\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23888\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23881\ : std_logic;
signal \N__23880\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23863\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23854\ : std_logic;
signal \N__23851\ : std_logic;
signal \N__23848\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23829\ : std_logic;
signal \N__23826\ : std_logic;
signal \N__23823\ : std_logic;
signal \N__23820\ : std_logic;
signal \N__23815\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23806\ : std_logic;
signal \N__23803\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23797\ : std_logic;
signal \N__23794\ : std_logic;
signal \N__23791\ : std_logic;
signal \N__23786\ : std_logic;
signal \N__23783\ : std_logic;
signal \N__23780\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23778\ : std_logic;
signal \N__23775\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23769\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23756\ : std_logic;
signal \N__23755\ : std_logic;
signal \N__23754\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23750\ : std_logic;
signal \N__23743\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23735\ : std_logic;
signal \N__23734\ : std_logic;
signal \N__23731\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23725\ : std_logic;
signal \N__23722\ : std_logic;
signal \N__23719\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23710\ : std_logic;
signal \N__23709\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23700\ : std_logic;
signal \N__23697\ : std_logic;
signal \N__23692\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23684\ : std_logic;
signal \N__23683\ : std_logic;
signal \N__23680\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23677\ : std_logic;
signal \N__23676\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23674\ : std_logic;
signal \N__23673\ : std_logic;
signal \N__23672\ : std_logic;
signal \N__23671\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23665\ : std_logic;
signal \N__23662\ : std_logic;
signal \N__23659\ : std_logic;
signal \N__23656\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23649\ : std_logic;
signal \N__23648\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23642\ : std_logic;
signal \N__23641\ : std_logic;
signal \N__23638\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23636\ : std_logic;
signal \N__23635\ : std_logic;
signal \N__23632\ : std_logic;
signal \N__23631\ : std_logic;
signal \N__23628\ : std_logic;
signal \N__23623\ : std_logic;
signal \N__23616\ : std_logic;
signal \N__23613\ : std_logic;
signal \N__23610\ : std_logic;
signal \N__23607\ : std_logic;
signal \N__23604\ : std_logic;
signal \N__23601\ : std_logic;
signal \N__23598\ : std_logic;
signal \N__23595\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23586\ : std_logic;
signal \N__23585\ : std_logic;
signal \N__23582\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23578\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23566\ : std_logic;
signal \N__23563\ : std_logic;
signal \N__23560\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23526\ : std_logic;
signal \N__23517\ : std_logic;
signal \N__23514\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23497\ : std_logic;
signal \N__23494\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23490\ : std_logic;
signal \N__23489\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23462\ : std_logic;
signal \N__23461\ : std_logic;
signal \N__23458\ : std_logic;
signal \N__23455\ : std_logic;
signal \N__23452\ : std_logic;
signal \N__23449\ : std_logic;
signal \N__23446\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23426\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23420\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23414\ : std_logic;
signal \N__23411\ : std_logic;
signal \N__23408\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23402\ : std_logic;
signal \N__23399\ : std_logic;
signal \N__23396\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23384\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23357\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23309\ : std_logic;
signal \N__23306\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23291\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23270\ : std_logic;
signal \N__23267\ : std_logic;
signal \N__23264\ : std_logic;
signal \N__23261\ : std_logic;
signal \N__23258\ : std_logic;
signal \N__23255\ : std_logic;
signal \N__23252\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23243\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23237\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23219\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23213\ : std_logic;
signal \N__23210\ : std_logic;
signal \N__23207\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23198\ : std_logic;
signal \N__23195\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23186\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23180\ : std_logic;
signal \N__23177\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23165\ : std_logic;
signal \N__23162\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23156\ : std_logic;
signal \N__23153\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23147\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23135\ : std_logic;
signal \N__23132\ : std_logic;
signal \N__23129\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23120\ : std_logic;
signal \N__23117\ : std_logic;
signal \N__23114\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23102\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23084\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23063\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23038\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23028\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23026\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23018\ : std_logic;
signal \N__23015\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__23002\ : std_logic;
signal \N__22999\ : std_logic;
signal \N__22996\ : std_logic;
signal \N__22993\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22976\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22967\ : std_logic;
signal \N__22964\ : std_logic;
signal \N__22961\ : std_logic;
signal \N__22958\ : std_logic;
signal \N__22955\ : std_logic;
signal \N__22952\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22940\ : std_logic;
signal \N__22937\ : std_logic;
signal \N__22934\ : std_logic;
signal \N__22931\ : std_logic;
signal \N__22928\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22889\ : std_logic;
signal \N__22886\ : std_logic;
signal \N__22883\ : std_logic;
signal \N__22880\ : std_logic;
signal \N__22877\ : std_logic;
signal \N__22874\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22844\ : std_logic;
signal \N__22841\ : std_logic;
signal \N__22838\ : std_logic;
signal \N__22835\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22829\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22811\ : std_logic;
signal \N__22808\ : std_logic;
signal \N__22805\ : std_logic;
signal \N__22802\ : std_logic;
signal \N__22799\ : std_logic;
signal \N__22796\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22790\ : std_logic;
signal \N__22787\ : std_logic;
signal \N__22784\ : std_logic;
signal \N__22781\ : std_logic;
signal \N__22778\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22757\ : std_logic;
signal \N__22754\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22741\ : std_logic;
signal \N__22740\ : std_logic;
signal \N__22739\ : std_logic;
signal \N__22738\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22732\ : std_logic;
signal \N__22727\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22725\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22722\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22719\ : std_logic;
signal \N__22714\ : std_logic;
signal \N__22699\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22689\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22687\ : std_logic;
signal \N__22686\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22684\ : std_logic;
signal \N__22683\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22669\ : std_logic;
signal \N__22666\ : std_logic;
signal \N__22663\ : std_logic;
signal \N__22658\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22638\ : std_logic;
signal \N__22625\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22623\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22613\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22608\ : std_logic;
signal \N__22605\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22595\ : std_logic;
signal \N__22592\ : std_logic;
signal \N__22591\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22581\ : std_logic;
signal \N__22578\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22576\ : std_logic;
signal \N__22575\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22554\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22552\ : std_logic;
signal \N__22551\ : std_logic;
signal \N__22546\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22523\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22495\ : std_logic;
signal \N__22490\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22479\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22465\ : std_logic;
signal \N__22462\ : std_logic;
signal \N__22459\ : std_logic;
signal \N__22456\ : std_logic;
signal \N__22453\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22447\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22441\ : std_logic;
signal \N__22436\ : std_logic;
signal \N__22433\ : std_logic;
signal \N__22430\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22424\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22394\ : std_logic;
signal \N__22391\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22292\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22268\ : std_logic;
signal \N__22265\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22238\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22214\ : std_logic;
signal \N__22211\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22181\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22148\ : std_logic;
signal \N__22145\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22136\ : std_logic;
signal \N__22133\ : std_logic;
signal \N__22130\ : std_logic;
signal \N__22127\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22103\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22082\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22012\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21988\ : std_logic;
signal \N__21985\ : std_logic;
signal \N__21982\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21907\ : std_logic;
signal \N__21906\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21901\ : std_logic;
signal \N__21900\ : std_logic;
signal \N__21897\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21878\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21859\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21842\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21836\ : std_logic;
signal \N__21833\ : std_logic;
signal \N__21830\ : std_logic;
signal \N__21827\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21809\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21743\ : std_logic;
signal \N__21740\ : std_logic;
signal \N__21737\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21705\ : std_logic;
signal \N__21702\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21694\ : std_logic;
signal \N__21685\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21655\ : std_logic;
signal \N__21652\ : std_logic;
signal \N__21649\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21586\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21575\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21560\ : std_logic;
signal \N__21557\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21536\ : std_logic;
signal \N__21533\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21515\ : std_logic;
signal \N__21512\ : std_logic;
signal \N__21509\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21503\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21488\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21472\ : std_logic;
signal \N__21467\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21462\ : std_logic;
signal \N__21459\ : std_logic;
signal \N__21456\ : std_logic;
signal \N__21453\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21443\ : std_logic;
signal \N__21442\ : std_logic;
signal \N__21439\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21426\ : std_logic;
signal \N__21425\ : std_logic;
signal \N__21422\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21411\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21385\ : std_logic;
signal \N__21382\ : std_logic;
signal \N__21377\ : std_logic;
signal \N__21374\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21370\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21358\ : std_logic;
signal \N__21355\ : std_logic;
signal \N__21352\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21346\ : std_logic;
signal \N__21343\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21334\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21328\ : std_logic;
signal \N__21323\ : std_logic;
signal \N__21320\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21316\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21308\ : std_logic;
signal \N__21305\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21298\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21286\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21275\ : std_logic;
signal \N__21272\ : std_logic;
signal \N__21269\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21267\ : std_logic;
signal \N__21266\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21262\ : std_logic;
signal \N__21259\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21257\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21242\ : std_logic;
signal \N__21237\ : std_logic;
signal \N__21226\ : std_logic;
signal \N__21223\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21217\ : std_logic;
signal \N__21214\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21201\ : std_logic;
signal \N__21198\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21192\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21178\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21166\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21154\ : std_logic;
signal \N__21151\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21133\ : std_logic;
signal \N__21130\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21121\ : std_logic;
signal \N__21118\ : std_logic;
signal \N__21115\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21094\ : std_logic;
signal \N__21091\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21068\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21062\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21058\ : std_logic;
signal \N__21057\ : std_logic;
signal \N__21054\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21045\ : std_logic;
signal \N__21042\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21025\ : std_logic;
signal \N__21024\ : std_logic;
signal \N__21021\ : std_logic;
signal \N__21018\ : std_logic;
signal \N__21015\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21009\ : std_logic;
signal \N__21006\ : std_logic;
signal \N__21001\ : std_logic;
signal \N__20998\ : std_logic;
signal \N__20995\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20980\ : std_logic;
signal \N__20977\ : std_logic;
signal \N__20976\ : std_logic;
signal \N__20973\ : std_logic;
signal \N__20970\ : std_logic;
signal \N__20967\ : std_logic;
signal \N__20964\ : std_logic;
signal \N__20961\ : std_logic;
signal \N__20956\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20947\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20920\ : std_logic;
signal \N__20917\ : std_logic;
signal \N__20914\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20905\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20891\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20887\ : std_logic;
signal \N__20884\ : std_logic;
signal \N__20881\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20872\ : std_logic;
signal \N__20869\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20861\ : std_logic;
signal \N__20860\ : std_logic;
signal \N__20859\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20857\ : std_logic;
signal \N__20856\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20854\ : std_logic;
signal \N__20851\ : std_logic;
signal \N__20848\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20843\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20820\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20795\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20784\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20776\ : std_logic;
signal \N__20775\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20773\ : std_logic;
signal \N__20772\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20769\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20763\ : std_logic;
signal \N__20754\ : std_logic;
signal \N__20747\ : std_logic;
signal \N__20744\ : std_logic;
signal \N__20737\ : std_logic;
signal \N__20734\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20726\ : std_logic;
signal \N__20725\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20723\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20721\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20712\ : std_logic;
signal \N__20709\ : std_logic;
signal \N__20706\ : std_logic;
signal \N__20703\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20680\ : std_logic;
signal \N__20677\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20662\ : std_logic;
signal \N__20657\ : std_logic;
signal \N__20654\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20648\ : std_logic;
signal \N__20645\ : std_logic;
signal \N__20642\ : std_logic;
signal \N__20639\ : std_logic;
signal \N__20636\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20630\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20618\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20603\ : std_logic;
signal \N__20600\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20590\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20584\ : std_logic;
signal \N__20583\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20563\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20541\ : std_logic;
signal \N__20540\ : std_logic;
signal \N__20537\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20523\ : std_logic;
signal \N__20520\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20509\ : std_logic;
signal \N__20504\ : std_logic;
signal \N__20501\ : std_logic;
signal \N__20498\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20493\ : std_logic;
signal \N__20490\ : std_logic;
signal \N__20487\ : std_logic;
signal \N__20484\ : std_logic;
signal \N__20477\ : std_logic;
signal \N__20474\ : std_logic;
signal \N__20471\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20464\ : std_logic;
signal \N__20463\ : std_logic;
signal \N__20460\ : std_logic;
signal \N__20457\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20451\ : std_logic;
signal \N__20448\ : std_logic;
signal \N__20443\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20431\ : std_logic;
signal \N__20428\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20410\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20402\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20387\ : std_logic;
signal \N__20384\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20356\ : std_logic;
signal \N__20353\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20335\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20326\ : std_logic;
signal \N__20323\ : std_logic;
signal \N__20320\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20311\ : std_logic;
signal \N__20308\ : std_logic;
signal \N__20305\ : std_logic;
signal \N__20302\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20290\ : std_logic;
signal \N__20287\ : std_logic;
signal \N__20284\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20272\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20261\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20243\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20231\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20201\ : std_logic;
signal \N__20198\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20194\ : std_logic;
signal \N__20191\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20175\ : std_logic;
signal \N__20172\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20149\ : std_logic;
signal \N__20146\ : std_logic;
signal \N__20143\ : std_logic;
signal \N__20140\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20136\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20133\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20127\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20108\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20094\ : std_logic;
signal \N__20091\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20080\ : std_logic;
signal \N__20077\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20038\ : std_logic;
signal \N__20035\ : std_logic;
signal \N__20032\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20018\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20009\ : std_logic;
signal \N__20006\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__20001\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19986\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19978\ : std_logic;
signal \N__19975\ : std_logic;
signal \N__19972\ : std_logic;
signal \N__19969\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19943\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19882\ : std_logic;
signal \N__19879\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19865\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19859\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19832\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19820\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19795\ : std_logic;
signal \N__19792\ : std_logic;
signal \N__19789\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19780\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19776\ : std_logic;
signal \N__19773\ : std_logic;
signal \N__19770\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19738\ : std_logic;
signal \N__19737\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19726\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19720\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19714\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19708\ : std_logic;
signal \N__19705\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19686\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19662\ : std_logic;
signal \N__19659\ : std_logic;
signal \N__19654\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19621\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19609\ : std_logic;
signal \N__19606\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19585\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19574\ : std_logic;
signal \N__19571\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19567\ : std_logic;
signal \N__19566\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19558\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19546\ : std_logic;
signal \N__19543\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19536\ : std_logic;
signal \N__19533\ : std_logic;
signal \N__19530\ : std_logic;
signal \N__19527\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19514\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19498\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19489\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19485\ : std_logic;
signal \N__19482\ : std_logic;
signal \N__19479\ : std_logic;
signal \N__19476\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19444\ : std_logic;
signal \N__19443\ : std_logic;
signal \N__19440\ : std_logic;
signal \N__19437\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19426\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19406\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19400\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19321\ : std_logic;
signal \N__19318\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19312\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19304\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19280\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19262\ : std_logic;
signal \N__19259\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19244\ : std_logic;
signal \N__19241\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19223\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19196\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19169\ : std_logic;
signal \N__19166\ : std_logic;
signal \N__19163\ : std_logic;
signal \N__19160\ : std_logic;
signal \N__19157\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19145\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19138\ : std_logic;
signal \N__19137\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19129\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19117\ : std_logic;
signal \N__19116\ : std_logic;
signal \N__19113\ : std_logic;
signal \N__19108\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19100\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19096\ : std_logic;
signal \N__19095\ : std_logic;
signal \N__19092\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19086\ : std_logic;
signal \N__19083\ : std_logic;
signal \N__19080\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19063\ : std_logic;
signal \N__19062\ : std_logic;
signal \N__19059\ : std_logic;
signal \N__19056\ : std_logic;
signal \N__19053\ : std_logic;
signal \N__19050\ : std_logic;
signal \N__19043\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19034\ : std_logic;
signal \N__19031\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19027\ : std_logic;
signal \N__19026\ : std_logic;
signal \N__19019\ : std_logic;
signal \N__19016\ : std_logic;
signal \N__19015\ : std_logic;
signal \N__19012\ : std_logic;
signal \N__19009\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__19003\ : std_logic;
signal \N__19002\ : std_logic;
signal \N__18999\ : std_logic;
signal \N__18996\ : std_logic;
signal \N__18993\ : std_logic;
signal \N__18986\ : std_logic;
signal \N__18983\ : std_logic;
signal \N__18982\ : std_logic;
signal \N__18979\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18971\ : std_logic;
signal \N__18970\ : std_logic;
signal \N__18967\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18956\ : std_logic;
signal \N__18953\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18951\ : std_logic;
signal \N__18950\ : std_logic;
signal \N__18949\ : std_logic;
signal \N__18948\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18946\ : std_logic;
signal \N__18945\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18943\ : std_logic;
signal \N__18942\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18940\ : std_logic;
signal \N__18939\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18915\ : std_logic;
signal \N__18900\ : std_logic;
signal \N__18897\ : std_logic;
signal \N__18892\ : std_logic;
signal \N__18891\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18889\ : std_logic;
signal \N__18888\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18886\ : std_logic;
signal \N__18885\ : std_logic;
signal \N__18880\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18868\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18856\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18848\ : std_logic;
signal \N__18847\ : std_logic;
signal \N__18846\ : std_logic;
signal \N__18843\ : std_logic;
signal \N__18840\ : std_logic;
signal \N__18837\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18824\ : std_logic;
signal \N__18821\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18803\ : std_logic;
signal \N__18800\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18770\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18755\ : std_logic;
signal \N__18752\ : std_logic;
signal \N__18749\ : std_logic;
signal \N__18746\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18734\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18728\ : std_logic;
signal \N__18725\ : std_logic;
signal \N__18722\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18707\ : std_logic;
signal \N__18704\ : std_logic;
signal \N__18701\ : std_logic;
signal \N__18698\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18689\ : std_logic;
signal \N__18688\ : std_logic;
signal \N__18687\ : std_logic;
signal \N__18686\ : std_logic;
signal \N__18685\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18681\ : std_logic;
signal \N__18678\ : std_logic;
signal \N__18677\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18668\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18647\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18638\ : std_logic;
signal \N__18635\ : std_logic;
signal \N__18632\ : std_logic;
signal \N__18629\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18620\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18614\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18608\ : std_logic;
signal \N__18605\ : std_logic;
signal \N__18602\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18596\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18587\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18581\ : std_logic;
signal \N__18578\ : std_logic;
signal \N__18575\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18569\ : std_logic;
signal \N__18566\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18548\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18542\ : std_logic;
signal \N__18539\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18470\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18458\ : std_logic;
signal \N__18455\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18425\ : std_logic;
signal \N__18422\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18416\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18350\ : std_logic;
signal \N__18347\ : std_logic;
signal \N__18344\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18329\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18323\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18319\ : std_logic;
signal \N__18314\ : std_logic;
signal \N__18311\ : std_logic;
signal \N__18308\ : std_logic;
signal \N__18305\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18293\ : std_logic;
signal \N__18290\ : std_logic;
signal \N__18287\ : std_logic;
signal \N__18284\ : std_logic;
signal \N__18281\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18275\ : std_logic;
signal \N__18272\ : std_logic;
signal \N__18269\ : std_logic;
signal \N__18266\ : std_logic;
signal \N__18263\ : std_logic;
signal \N__18260\ : std_logic;
signal \N__18257\ : std_logic;
signal \N__18254\ : std_logic;
signal \N__18251\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18245\ : std_logic;
signal \N__18242\ : std_logic;
signal \N__18239\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18233\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18224\ : std_logic;
signal \N__18221\ : std_logic;
signal \N__18218\ : std_logic;
signal \N__18215\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18206\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18191\ : std_logic;
signal \N__18188\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18182\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18176\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18164\ : std_logic;
signal \N__18161\ : std_logic;
signal \N__18158\ : std_logic;
signal \N__18155\ : std_logic;
signal \N__18152\ : std_logic;
signal \N__18149\ : std_logic;
signal \N__18146\ : std_logic;
signal \N__18145\ : std_logic;
signal \N__18144\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18134\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_97\ : std_logic;
signal \bfn_1_9_0_\ : std_logic;
signal \pwm_generator_inst.O_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_0\ : std_logic;
signal \pwm_generator_inst.O_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_1\ : std_logic;
signal \pwm_generator_inst.O_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_2\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_3\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_4\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_5\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_6\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_7\ : std_logic;
signal \bfn_1_10_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_9\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_10\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_15\ : std_logic;
signal \bfn_1_11_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_16\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_17\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_18\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_19\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_1_15\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4\ : std_logic;
signal \bfn_1_12_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_17\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_18\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_19\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_20\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_21\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_22\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_23\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0\ : std_logic;
signal \bfn_1_13_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_24\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_25\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_15\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO\ : std_logic;
signal \bfn_1_14_0_\ : std_logic;
signal \N_110_i_i\ : std_logic;
signal un7_start_stop : std_logic;
signal pwm_duty_input_5 : std_logic;
signal pwm_duty_input_9 : std_logic;
signal pwm_duty_input_8 : std_logic;
signal \current_shift_inst.PI_CTRL.m7_2\ : std_logic;
signal pwm_duty_input_7 : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_0_3\ : std_logic;
signal pwm_duty_input_1 : std_logic;
signal pwm_duty_input_3 : std_logic;
signal pwm_duty_input_0 : std_logic;
signal pwm_duty_input_2 : std_logic;
signal \current_shift_inst.PI_CTRL.m14_2\ : std_logic;
signal pwm_duty_input_10 : std_logic;
signal \current_shift_inst.PI_CTRL.N_19_cascade_\ : std_logic;
signal pwm_duty_input_4 : std_logic;
signal \pwm_generator_inst.O_0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_0\ : std_logic;
signal \bfn_2_7_0_\ : std_logic;
signal \pwm_generator_inst.O_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_0\ : std_logic;
signal \pwm_generator_inst.O_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_1\ : std_logic;
signal \pwm_generator_inst.O_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_2\ : std_logic;
signal \pwm_generator_inst.O_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_3\ : std_logic;
signal \pwm_generator_inst.O_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_4\ : std_logic;
signal \pwm_generator_inst.O_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_5\ : std_logic;
signal \pwm_generator_inst.O_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_7\ : std_logic;
signal \pwm_generator_inst.O_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_8\ : std_logic;
signal \bfn_2_8_0_\ : std_logic;
signal \pwm_generator_inst.O_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_15\ : std_logic;
signal \bfn_2_9_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_18\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_17\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_18\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_18_cascade_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_16\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_13\ : std_logic;
signal \pwm_generator_inst.O_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_98_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_96\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_178\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_91\ : std_logic;
signal \un2_counter_7_cascade_\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_0\ : std_logic;
signal \bfn_3_9_0_\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_2\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_7\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_7\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_8\ : std_logic;
signal \bfn_3_10_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_8\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_9_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_118\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\ : std_logic;
signal \bfn_4_7_0_\ : std_logic;
signal un5_counter_cry_1 : std_logic;
signal \counterZ0Z_3\ : std_logic;
signal un5_counter_cry_2 : std_logic;
signal \counterZ0Z_4\ : std_logic;
signal un5_counter_cry_3 : std_logic;
signal \counterZ0Z_5\ : std_logic;
signal un5_counter_cry_4 : std_logic;
signal \counterZ0Z_6\ : std_logic;
signal un5_counter_cry_5 : std_logic;
signal un5_counter_cry_6 : std_logic;
signal \counterZ0Z_8\ : std_logic;
signal un5_counter_cry_7 : std_logic;
signal un5_counter_cry_8 : std_logic;
signal \counterZ0Z_9\ : std_logic;
signal \bfn_4_8_0_\ : std_logic;
signal un5_counter_cry_9 : std_logic;
signal \counterZ0Z_11\ : std_logic;
signal un5_counter_cry_10 : std_logic;
signal \counterZ0Z_12\ : std_logic;
signal un5_counter_cry_11 : std_logic;
signal \counter_RNO_0Z0Z_12\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5\ : std_logic;
signal pwm_duty_input_6 : std_logic;
signal \N_28_mux\ : std_logic;
signal i8_mux : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\ : std_logic;
signal \bfn_4_13_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\ : std_logic;
signal \bfn_4_14_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\ : std_logic;
signal \bfn_4_15_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\ : std_logic;
signal \bfn_4_16_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un8_enablelto31\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_12\ : std_logic;
signal \counter_RNO_0Z0Z_7\ : std_logic;
signal \counterZ0Z_7\ : std_logic;
signal \counterZ0Z_1\ : std_logic;
signal \counterZ0Z_2\ : std_logic;
signal \un2_counter_5_cascade_\ : std_logic;
signal \counterZ0Z_0\ : std_logic;
signal \un2_counter_9_cascade_\ : std_logic;
signal \clk_10khz_RNIIENAZ0Z2_cascade_\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_2\ : std_logic;
signal un2_counter_8 : std_logic;
signal \counter_RNO_0Z0Z_10\ : std_logic;
signal un2_counter_9 : std_logic;
signal un2_counter_7 : std_logic;
signal \counterZ0Z_10\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_10_31_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_11_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_9_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_8_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_25\ : std_logic;
signal clk_10khz_i : std_logic;
signal \clk_10khz_RNIIENAZ0Z2\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_7\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_1\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_4\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_2_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_47_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_43\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_46_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_46_21_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_44\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_7\ : std_logic;
signal \bfn_7_17_0_\ : std_logic;
signal \current_shift_inst.control_input_1_cry_0\ : std_logic;
signal \current_shift_inst.control_input_1_cry_1\ : std_logic;
signal \current_shift_inst.control_input_1_cry_2\ : std_logic;
signal \current_shift_inst.control_input_1_cry_3\ : std_logic;
signal \current_shift_inst.control_input_1_cry_4\ : std_logic;
signal \current_shift_inst.control_input_1_cry_5\ : std_logic;
signal \current_shift_inst.control_input_1_cry_6\ : std_logic;
signal \current_shift_inst.control_input_1_cry_7\ : std_logic;
signal \bfn_7_18_0_\ : std_logic;
signal \current_shift_inst.control_input_1_cry_8\ : std_logic;
signal \current_shift_inst.control_input_1_cry_9\ : std_logic;
signal \current_shift_inst.control_input_1_cry_10\ : std_logic;
signal \current_shift_inst.control_input_1_cry_11\ : std_logic;
signal \current_shift_inst.control_input_1_cry_12\ : std_logic;
signal \current_shift_inst.control_input_1_cry_13\ : std_logic;
signal \current_shift_inst.control_input_1_cry_14\ : std_logic;
signal \current_shift_inst.control_input_1_cry_15\ : std_logic;
signal \bfn_7_19_0_\ : std_logic;
signal \current_shift_inst.control_input_1_cry_16\ : std_logic;
signal \current_shift_inst.control_input_1_cry_17\ : std_logic;
signal \current_shift_inst.control_input_1_cry_18\ : std_logic;
signal \current_shift_inst.control_input_1_cry_19\ : std_logic;
signal \current_shift_inst.control_input_1_cry_20\ : std_logic;
signal \current_shift_inst.control_input_1_cry_21\ : std_logic;
signal \current_shift_inst.control_input_1_cry_22\ : std_logic;
signal \current_shift_inst.control_input_1_cry_23\ : std_logic;
signal \bfn_7_20_0_\ : std_logic;
signal \current_shift_inst.control_input_1_cry_24\ : std_logic;
signal il_min_comp2_c : std_logic;
signal il_max_comp2_c : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_0\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_6\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_3\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_5\ : std_logic;
signal \bfn_8_11_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ1Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \bfn_8_12_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_16\ : std_logic;
signal \bfn_8_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_enablelt3_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_47_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_46_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_76\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_75\ : std_logic;
signal \bfn_8_17_0_\ : std_logic;
signal \current_shift_inst.z_i_0_31\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CO\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_3_c_invZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_2\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_3\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0Z_0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_4\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIVQKU1_5\ : std_logic;
signal \current_shift_inst.control_input_1_axb_0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_5\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_6\ : std_logic;
signal \current_shift_inst.control_input_1_axb_1\ : std_logic;
signal \bfn_8_18_0_\ : std_logic;
signal \current_shift_inst.control_input_1_axb_2\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_7\ : std_logic;
signal \current_shift_inst.control_input_1_axb_3\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_8\ : std_logic;
signal \current_shift_inst.control_input_1_axb_4\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_9\ : std_logic;
signal \current_shift_inst.control_input_1_axb_5\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_10\ : std_logic;
signal \current_shift_inst.control_input_1_axb_6\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_11\ : std_logic;
signal \current_shift_inst.control_input_1_axb_7\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIR0UI_13\ : std_logic;
signal \current_shift_inst.control_input_1_axb_8\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_13\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_14\ : std_logic;
signal \current_shift_inst.control_input_1_axb_9\ : std_logic;
signal \bfn_8_19_0_\ : std_logic;
signal \current_shift_inst.control_input_1_axb_10\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_15\ : std_logic;
signal \current_shift_inst.control_input_1_axb_11\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIH6661_17\ : std_logic;
signal \current_shift_inst.control_input_1_axb_12\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIAL3J_18\ : std_logic;
signal \current_shift_inst.control_input_1_axb_13\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI4H5J_19\ : std_logic;
signal \current_shift_inst.control_input_1_axb_14\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_19\ : std_logic;
signal \current_shift_inst.control_input_1_axb_15\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_20\ : std_logic;
signal \current_shift_inst.control_input_1_axb_16\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_21\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_22\ : std_logic;
signal \current_shift_inst.control_input_1_axb_17\ : std_logic;
signal \bfn_8_20_0_\ : std_logic;
signal \current_shift_inst.control_input_1_axb_18\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_23\ : std_logic;
signal \current_shift_inst.control_input_1_axb_19\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_24\ : std_logic;
signal \current_shift_inst.control_input_1_axb_20\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_25\ : std_logic;
signal \current_shift_inst.control_input_1_axb_21\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_26\ : std_logic;
signal \current_shift_inst.control_input_1_axb_22\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_27\ : std_logic;
signal \current_shift_inst.control_input_1_axb_23\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_28\ : std_logic;
signal \current_shift_inst.control_input_1_axb_24\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_29\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_30\ : std_logic;
signal \current_shift_inst.control_input_1_cry_24_THRU_CO\ : std_logic;
signal \bfn_8_21_0_\ : std_logic;
signal \current_shift_inst.phase_valid_RNISLORZ0Z2\ : std_logic;
signal \il_min_comp2_D1\ : std_logic;
signal il_max_comp1_c : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_0\ : std_logic;
signal \pwm_generator_inst.counter_i_0\ : std_logic;
signal \bfn_9_8_0_\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_1\ : std_logic;
signal \pwm_generator_inst.counter_i_1\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_0\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counter_i_2\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_1\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_3\ : std_logic;
signal \pwm_generator_inst.counter_i_3\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_2\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_4\ : std_logic;
signal \pwm_generator_inst.counter_i_4\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_3\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_5\ : std_logic;
signal \pwm_generator_inst.counter_i_5\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_4\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_6\ : std_logic;
signal \pwm_generator_inst.counter_i_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_5\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_7\ : std_logic;
signal \pwm_generator_inst.counter_i_7\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_7\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_8\ : std_logic;
signal \pwm_generator_inst.counter_i_8\ : std_logic;
signal \bfn_9_9_0_\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_9\ : std_logic;
signal \pwm_generator_inst.counter_i_9\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_8\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_9\ : std_logic;
signal pwm_output_c : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_0\ : std_logic;
signal \bfn_9_13_0_\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_0\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_2\ : std_logic;
signal \N_702_g\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_4\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_5\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_6\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_5\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_8\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\ : std_logic;
signal \bfn_9_14_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_9\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_10\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_11\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_12\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_13\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_12\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_15\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_16\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\ : std_logic;
signal \bfn_9_15_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_17\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_18\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_19\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_20\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_21\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_22\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_23\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_24\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\ : std_logic;
signal \bfn_9_16_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_29\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.N_1717_i\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_2_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3_cascade_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_4_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIK3CV_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIP5T51_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIER9V_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJDBL1_10\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIE6961_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIHVAV_6\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI7DM51_10\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI53NU1_6\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI7H2J_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIIKQI_10\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIU4VI_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIBU361_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIBBPU1_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI1PG21_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNINKG81_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIR32K_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPB581_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJ3381_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIVQF91_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIAO7K_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI4D1J_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIKKJ81_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIHCE81_26\ : std_logic;
signal \bfn_9_21_0_\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \bfn_9_22_0_\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \bfn_9_23_0_\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \bfn_9_24_0_\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \current_shift_inst.timer_phase.N_188_i_g\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_0\ : std_logic;
signal \bfn_9_25_0_\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_1\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_0\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_2\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_1\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_3\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_2\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_4\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_3\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_5\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_4\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_6\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_5\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_7\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_6\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_7\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_8\ : std_logic;
signal \bfn_9_26_0_\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_9\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_8\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_10\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_9\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_11\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_10\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_12\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_11\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_13\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_12\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_14\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_13\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_15\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_14\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_15\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_16\ : std_logic;
signal \bfn_9_27_0_\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_17\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_16\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_18\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_17\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_19\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_18\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_20\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_19\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_21\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_20\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_22\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_21\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_23\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_22\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_23\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_24\ : std_logic;
signal \bfn_9_28_0_\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_25\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_24\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_26\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_25\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_27\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_26\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_28\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_27\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_28\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_29\ : std_logic;
signal \il_max_comp1_D1\ : std_logic;
signal \pwm_generator_inst.un1_counterlto2_0_cascade_\ : std_logic;
signal \pwm_generator_inst.un1_counterlt9_cascade_\ : std_logic;
signal \pwm_generator_inst.un1_counterlto9_2\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_0\ : std_logic;
signal \bfn_10_9_0_\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_1\ : std_logic;
signal \pwm_generator_inst.counter_cry_0\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counter_cry_1\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_3\ : std_logic;
signal \pwm_generator_inst.counter_cry_2\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_4\ : std_logic;
signal \pwm_generator_inst.counter_cry_3\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_5\ : std_logic;
signal \pwm_generator_inst.counter_cry_4\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_6\ : std_logic;
signal \pwm_generator_inst.counter_cry_5\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_7\ : std_logic;
signal \pwm_generator_inst.counter_cry_6\ : std_logic;
signal \pwm_generator_inst.counter_cry_7\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_8\ : std_logic;
signal \bfn_10_10_0_\ : std_logic;
signal \pwm_generator_inst.un1_counter_0\ : std_logic;
signal \pwm_generator_inst.counter_cry_8\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.time_passed11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa\ : std_logic;
signal \G_407\ : std_logic;
signal \bfn_10_14_0_\ : std_logic;
signal \G_406\ : std_logic;
signal \current_shift_inst.z_cry_0\ : std_logic;
signal \current_shift_inst.z_cry_1\ : std_logic;
signal \current_shift_inst.z_cry_2\ : std_logic;
signal \current_shift_inst.z_cry_3\ : std_logic;
signal \current_shift_inst.z_cry_4\ : std_logic;
signal \current_shift_inst.z_cry_5\ : std_logic;
signal \current_shift_inst.z_cry_6\ : std_logic;
signal \current_shift_inst.z_cry_7\ : std_logic;
signal \bfn_10_15_0_\ : std_logic;
signal \current_shift_inst.z_cry_8\ : std_logic;
signal \current_shift_inst.z_cry_9\ : std_logic;
signal \current_shift_inst.z_cry_10\ : std_logic;
signal \current_shift_inst.z_cry_11\ : std_logic;
signal \current_shift_inst.z_cry_12\ : std_logic;
signal \current_shift_inst.z_cry_13\ : std_logic;
signal \current_shift_inst.z_cry_14\ : std_logic;
signal \current_shift_inst.z_cry_15\ : std_logic;
signal \bfn_10_16_0_\ : std_logic;
signal \current_shift_inst.z_cry_16\ : std_logic;
signal \current_shift_inst.z_cry_17\ : std_logic;
signal \current_shift_inst.z_cry_18\ : std_logic;
signal \current_shift_inst.z_cry_19\ : std_logic;
signal \current_shift_inst.z_cry_20\ : std_logic;
signal \current_shift_inst.z_cry_21\ : std_logic;
signal \current_shift_inst.z_cry_22\ : std_logic;
signal \current_shift_inst.z_cry_23\ : std_logic;
signal \bfn_10_17_0_\ : std_logic;
signal \current_shift_inst.z_cry_24\ : std_logic;
signal \current_shift_inst.z_cry_25\ : std_logic;
signal \current_shift_inst.z_cry_26\ : std_logic;
signal \current_shift_inst.z_cry_27\ : std_logic;
signal \current_shift_inst.z_cry_28\ : std_logic;
signal \current_shift_inst.z_cry_29\ : std_logic;
signal \current_shift_inst.z_cry_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_1\ : std_logic;
signal \bfn_10_18_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_2\ : std_logic;
signal \current_shift_inst.z_5_2\ : std_logic;
signal \current_shift_inst.z_5_cry_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_3\ : std_logic;
signal \current_shift_inst.z_5_3\ : std_logic;
signal \current_shift_inst.z_5_cry_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_4\ : std_logic;
signal \current_shift_inst.z_5_4\ : std_logic;
signal \current_shift_inst.z_5_cry_3\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_5\ : std_logic;
signal \current_shift_inst.z_5_5\ : std_logic;
signal \current_shift_inst.z_5_cry_4\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_6\ : std_logic;
signal \current_shift_inst.z_5_6\ : std_logic;
signal \current_shift_inst.z_5_cry_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_7\ : std_logic;
signal \current_shift_inst.z_5_7\ : std_logic;
signal \current_shift_inst.z_5_cry_6\ : std_logic;
signal \current_shift_inst.z_5_8\ : std_logic;
signal \current_shift_inst.z_5_cry_7\ : std_logic;
signal \current_shift_inst.z_5_cry_8\ : std_logic;
signal \current_shift_inst.z_5_9\ : std_logic;
signal \bfn_10_19_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_10\ : std_logic;
signal \current_shift_inst.z_5_10\ : std_logic;
signal \current_shift_inst.z_5_cry_9\ : std_logic;
signal \current_shift_inst.z_5_11\ : std_logic;
signal \current_shift_inst.z_5_cry_10\ : std_logic;
signal \current_shift_inst.z_5_12\ : std_logic;
signal \current_shift_inst.z_5_cry_11\ : std_logic;
signal \current_shift_inst.z_5_13\ : std_logic;
signal \current_shift_inst.z_5_cry_12\ : std_logic;
signal \current_shift_inst.z_5_14\ : std_logic;
signal \current_shift_inst.z_5_cry_13\ : std_logic;
signal \current_shift_inst.z_5_15\ : std_logic;
signal \current_shift_inst.z_5_cry_14\ : std_logic;
signal \current_shift_inst.z_5_16\ : std_logic;
signal \current_shift_inst.z_5_cry_15\ : std_logic;
signal \current_shift_inst.z_5_cry_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_17\ : std_logic;
signal \current_shift_inst.z_5_17\ : std_logic;
signal \bfn_10_20_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_18\ : std_logic;
signal \current_shift_inst.z_5_18\ : std_logic;
signal \current_shift_inst.z_5_cry_17\ : std_logic;
signal \current_shift_inst.z_5_19\ : std_logic;
signal \current_shift_inst.z_5_cry_18\ : std_logic;
signal \current_shift_inst.z_5_20\ : std_logic;
signal \current_shift_inst.z_5_cry_19\ : std_logic;
signal \current_shift_inst.z_5_21\ : std_logic;
signal \current_shift_inst.z_5_cry_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_22\ : std_logic;
signal \current_shift_inst.z_5_22\ : std_logic;
signal \current_shift_inst.z_5_cry_21\ : std_logic;
signal \current_shift_inst.z_5_23\ : std_logic;
signal \current_shift_inst.z_5_cry_22\ : std_logic;
signal \current_shift_inst.z_5_24\ : std_logic;
signal \current_shift_inst.z_5_cry_23\ : std_logic;
signal \current_shift_inst.z_5_cry_24\ : std_logic;
signal \current_shift_inst.z_5_25\ : std_logic;
signal \bfn_10_21_0_\ : std_logic;
signal \current_shift_inst.z_5_26\ : std_logic;
signal \current_shift_inst.z_5_cry_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_27\ : std_logic;
signal \current_shift_inst.z_5_27\ : std_logic;
signal \current_shift_inst.z_5_cry_26\ : std_logic;
signal \current_shift_inst.z_5_28\ : std_logic;
signal \current_shift_inst.z_5_cry_27\ : std_logic;
signal \current_shift_inst.z_5_29\ : std_logic;
signal \current_shift_inst.z_5_cry_28\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \current_shift_inst.z_5_30\ : std_logic;
signal \current_shift_inst.z_5_cry_29\ : std_logic;
signal \current_shift_inst.z_5_cry_30\ : std_logic;
signal \current_shift_inst.z_5_cry_30_THRU_CO\ : std_logic;
signal s4_phy_c : std_logic;
signal il_min_comp1_c : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_11_8_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7\ : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17\ : std_logic;
signal \bfn_11_10_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19\ : std_logic;
signal \il_min_comp1_D1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_fast_31\ : std_logic;
signal \current_shift_inst.un38_control_input_0\ : std_logic;
signal \bfn_11_14_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_1\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_2\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_3_c_RNINL4GZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_3\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_4\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_5\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_6\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_7\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_8\ : std_logic;
signal \bfn_11_15_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_9\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_10_c_RNIJLTGZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_10\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_11\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_12\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_13\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_14\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_15\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_16\ : std_logic;
signal \bfn_11_16_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_17\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_18\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_19\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_20\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_21\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_22\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_23\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_24\ : std_logic;
signal \bfn_11_17_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_25\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_26\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_27\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_28\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_29\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_9\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_9_c_RNIALDJZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIO0U12_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNILORI_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIOSSI_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_13\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJTQ51_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_8\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIN7DV_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_28\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIDS8K_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5S981_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_11\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIDLO51_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_31\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_axb_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_19\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPC571_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI190J_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_16\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5M161_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_14\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIVDV51_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIDR081_20\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNILRVJ_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_21\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIOV0K_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIU73K_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI7K6K_26\ : std_logic;
signal \il_max_comp2_D1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.start_timer_hc_0_sqmuxa_cascade_\ : std_logic;
signal \phase_controller_inst1.N_88\ : std_logic;
signal \phase_controller_inst1.hc_time_passed\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_5\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_6\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_3\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_4\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_1\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_1\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_2\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_2\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_24\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_15\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_11\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_19\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_10\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_12\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_14\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_18\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_29\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_22\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_26\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_27\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_30\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_21\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_25\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_20\ : std_logic;
signal \current_shift_inst.z_31\ : std_logic;
signal \current_shift_inst.z_i_31\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI1C4K_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_26\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIB4C81_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_25\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI4G5K_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_29\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI7OAK_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_24\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_23\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIVJ781_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1Z0Z_6_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6_cascade_\ : std_logic;
signal \phase_controller_slave.start_timer_hc_0_sqmuxa_cascade_\ : std_logic;
signal s3_phy_c : std_logic;
signal \phase_controller_slave.stateZ0Z_1\ : std_logic;
signal \il_min_comp2_D2\ : std_logic;
signal \il_max_comp2_D2\ : std_logic;
signal \phase_controller_slave.stateZ0Z_3\ : std_logic;
signal \current_shift_inst.timer_phase.N_192_i\ : std_logic;
signal \current_shift_inst.timer_phase.running_i\ : std_logic;
signal clk_12mhz : std_logic;
signal \GB_BUFFER_clk_12mhz_THRU_CO\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_321_i\ : std_logic;
signal \current_shift_inst.N_199_cascade_\ : std_logic;
signal \current_shift_inst.timer_s1.N_187_i\ : std_logic;
signal \current_shift_inst.phase_validZ0\ : std_logic;
signal \current_shift_inst.start_timer_sZ0Z1\ : std_logic;
signal \current_shift_inst.stop_timer_sZ0Z1\ : std_logic;
signal \current_shift_inst.meas_stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto5Z0Z_3_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlt8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_13\ : std_logic;
signal \il_max_comp1_D2\ : std_logic;
signal \phase_controller_inst1.N_86_cascade_\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_3\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_3\ : std_logic;
signal \bfn_13_13_0_\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_4\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_5\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_6\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_7\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_10\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_11\ : std_logic;
signal \bfn_13_14_0_\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_12\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_14\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_15\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_18\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_19\ : std_logic;
signal \bfn_13_15_0_\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_20\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_21\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_22\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_24\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_25\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_26\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_27\ : std_logic;
signal \bfn_13_16_0_\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_28\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_29\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_30\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.N_187_i_g\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.S1_riseZ0\ : std_logic;
signal s1_phy_c : std_logic;
signal \current_shift_inst.S1_syncZ0Z0\ : std_logic;
signal \current_shift_inst.S3_sync_prevZ0\ : std_logic;
signal \current_shift_inst.S3_riseZ0\ : std_logic;
signal \current_shift_inst.S1_syncZ0Z1\ : std_logic;
signal \current_shift_inst.S1_sync_prevZ0\ : std_logic;
signal \current_shift_inst.S3_syncZ0Z0\ : std_logic;
signal \current_shift_inst.S3_syncZ0Z1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13_cascade_\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_13_19_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_13_20_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_17\ : std_logic;
signal \bfn_13_21_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_19\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_slave.stateZ0Z_0\ : std_logic;
signal \phase_controller_slave.stateZ0Z_4\ : std_logic;
signal \phase_controller_slave.start_timer_tr_0_sqmuxa\ : std_logic;
signal \phase_controller_slave.N_210_cascade_\ : std_logic;
signal \phase_controller_slave.stoper_tr.time_passed11_cascade_\ : std_logic;
signal \phase_controller_slave.tr_time_passed\ : std_logic;
signal \phase_controller_slave.stoper_tr.time_passed_1_sqmuxa\ : std_logic;
signal \bfn_13_23_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7\ : std_logic;
signal \bfn_13_24_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15\ : std_logic;
signal \bfn_13_25_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19\ : std_logic;
signal \current_shift_inst.start_timer_phaseZ0\ : std_logic;
signal \current_shift_inst.timer_phase.runningZ0\ : std_logic;
signal \current_shift_inst.stop_timer_phaseZ0\ : std_logic;
signal \current_shift_inst.timer_phase.N_188_i\ : std_logic;
signal s2_phy_c : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_3_cascade_\ : std_logic;
signal \delay_measurement_inst.stop_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt14_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt30_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_2_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_2_tz\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a1_1_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_1_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto13_3Z0Z_1_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto13\ : std_logic;
signal measured_delay_hc_20 : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto30_2_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlt15\ : std_logic;
signal \delay_measurement_inst.tr_stateZ0Z_0\ : std_logic;
signal \delay_measurement_inst.prev_tr_sigZ0\ : std_logic;
signal \delay_measurement_inst.tr_state_RNIMR6LZ0Z_0_cascade_\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_2\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_8\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_8\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_23\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_23\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_9\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_9\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_16\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_16\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_17\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_17\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_13\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_13\ : std_logic;
signal measured_delay_hc_15 : std_logic;
signal measured_delay_hc_14 : std_logic;
signal measured_delay_hc_6 : std_logic;
signal measured_delay_hc_2 : std_logic;
signal measured_delay_hc_9 : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.time_passed_1_sqmuxa\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3Z0Z_3_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_5Z0Z_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.time_passed11_cascade_\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0\ : std_logic;
signal start_stop_c : std_logic;
signal shift_flag_start : std_logic;
signal \phase_controller_slave.un1_startZ0\ : std_logic;
signal \phase_controller_slave.stoper_tr.time_passed11\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_14_22_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7\ : std_logic;
signal \bfn_14_23_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15\ : std_logic;
signal \bfn_14_24_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18\ : std_logic;
signal delay_tr_input_c : std_logic;
signal delay_tr_d1 : std_logic;
signal delay_tr_d2 : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_4\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_1\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6\ : std_logic;
signal \bfn_15_7_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_11\ : std_logic;
signal \bfn_15_8_0_\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \bfn_15_9_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \bfn_15_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_321_i_g\ : std_logic;
signal measured_delay_hc_10 : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2\ : std_logic;
signal \current_shift_inst.timer_s1.runningZ0\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_3\ : std_logic;
signal measured_delay_hc_3 : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_4\ : std_logic;
signal measured_delay_hc_4 : std_logic;
signal \delay_measurement_inst.hc_stateZ0Z_0\ : std_logic;
signal \delay_measurement_inst.start_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.prev_hc_sigZ0\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_0\ : std_logic;
signal \bfn_15_13_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_1\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_0\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_2\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_1\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_3\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_4\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_5\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_7\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_8\ : std_logic;
signal \bfn_15_14_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_9\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_10\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_9\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_11\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_12\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_13\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_15\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_16\ : std_logic;
signal \bfn_15_15_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_17\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_18\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_17\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_19\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_20\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_21\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_23\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_24\ : std_logic;
signal \bfn_15_16_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_25\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_26\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_25\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_27\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_28\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.running_i\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_29\ : std_logic;
signal \current_shift_inst.timer_s1.N_191_i\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_0\ : std_logic;
signal \bfn_15_17_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ1Z_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \bfn_15_18_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_16\ : std_logic;
signal \bfn_15_19_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_18\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_19\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_slave.stoper_hc.time_passed11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_20_li\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3\ : std_logic;
signal \delay_measurement_inst.stop_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6\ : std_logic;
signal measured_delay_tr_7 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6\ : std_logic;
signal measured_delay_tr_8 : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_slave.start_timer_trZ0\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19\ : std_logic;
signal \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\ : std_logic;
signal \bfn_16_7_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\ : std_logic;
signal \bfn_16_8_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\ : std_logic;
signal \bfn_16_9_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\ : std_logic;
signal \bfn_16_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_322_i\ : std_logic;
signal measured_delay_hc_12 : std_logic;
signal measured_delay_hc_11 : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_6_cascade_\ : std_logic;
signal \delay_measurement_inst.tr_state_RNIMR6LZ0Z_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_375_cascade_\ : std_logic;
signal \delay_measurement_inst.N_265_i_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_6_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_364\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_6_19_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_0_19\ : std_logic;
signal \delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_409\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_400_cascade_\ : std_logic;
signal \delay_measurement_inst.N_394_1_cascade_\ : std_logic;
signal \delay_measurement_inst.N_394_1\ : std_logic;
signal measured_delay_tr_12 : std_logic;
signal measured_delay_tr_10 : std_logic;
signal measured_delay_tr_6 : std_logic;
signal measured_delay_tr_3 : std_logic;
signal measured_delay_tr_5 : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_1\ : std_logic;
signal measured_delay_tr_1 : std_logic;
signal measured_delay_tr_2 : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst1.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_slave.start_timer_hcZ0\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\ : std_logic;
signal red_c_i : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal measured_delay_hc_16 : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlt31\ : std_logic;
signal measured_delay_hc_1 : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_16_19_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_16_20_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_17\ : std_logic;
signal \bfn_16_21_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal measured_delay_tr_19 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal measured_delay_tr_11 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal measured_delay_tr_13 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal delay_hc_input_c : std_logic;
signal delay_hc_d1 : std_logic;
signal delay_hc_d2 : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_2\ : std_logic;
signal measured_delay_hc_25 : std_logic;
signal measured_delay_hc_26 : std_logic;
signal measured_delay_hc_23 : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_8\ : std_logic;
signal measured_delay_hc_8 : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_7\ : std_logic;
signal measured_delay_hc_7 : std_logic;
signal measured_delay_hc_24 : std_logic;
signal measured_delay_hc_0 : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_18\ : std_logic;
signal measured_delay_hc_18 : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto31_0_0\ : std_logic;
signal measured_delay_hc_19 : std_logic;
signal measured_delay_hc_21 : std_logic;
signal measured_delay_hc_22 : std_logic;
signal \delay_measurement_inst.un1_elapsed_time_hc\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3\ : std_logic;
signal measured_delay_hc_17 : std_logic;
signal \bfn_17_11_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_7\ : std_logic;
signal \bfn_17_12_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_15\ : std_logic;
signal \bfn_17_13_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_23\ : std_logic;
signal \bfn_17_14_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_324_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_7_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_4\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16\ : std_logic;
signal measured_delay_tr_17 : std_logic;
signal \delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20\ : std_logic;
signal measured_delay_tr_18 : std_logic;
signal \phase_controller_inst1.N_83\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_4\ : std_logic;
signal \phase_controller_inst1.N_83_cascade_\ : std_logic;
signal \phase_controller_inst1.T01_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa_cascade_\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_1\ : std_logic;
signal \phase_controller_inst1.tr_time_passed\ : std_logic;
signal \il_min_comp1_D2\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.time_passed11_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.time_passed11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa\ : std_logic;
signal measured_delay_tr_16 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal measured_delay_hc_29 : std_logic;
signal measured_delay_hc_28 : std_logic;
signal measured_delay_hc_30 : std_logic;
signal measured_delay_hc_27 : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_4\ : std_logic;
signal measured_delay_hc_13 : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal measured_delay_hc_31 : std_logic;
signal measured_delay_hc_5 : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlt31_0\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa\ : std_logic;
signal \delay_measurement_inst.N_410\ : std_logic;
signal \delay_measurement_inst.N_358\ : std_logic;
signal \delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15\ : std_logic;
signal measured_delay_tr_4 : std_logic;
signal \delay_measurement_inst.N_265_i_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_3\ : std_logic;
signal \bfn_18_13_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_11\ : std_logic;
signal \bfn_18_14_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_19\ : std_logic;
signal \bfn_18_15_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\ : std_logic;
signal \bfn_18_16_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_31\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_323_i\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_18_17_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7\ : std_logic;
signal \bfn_18_18_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17\ : std_logic;
signal \bfn_18_19_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_21\ : std_logic;
signal \delay_measurement_inst.N_271_1\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_14\ : std_logic;
signal \delay_measurement_inst.N_265_i\ : std_logic;
signal measured_delay_tr_14 : std_logic;
signal \phase_controller_slave.hc_time_passed\ : std_logic;
signal \phase_controller_slave.stateZ0Z_2\ : std_logic;
signal \phase_controller_slave.N_211\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13\ : std_logic;
signal measured_delay_tr_15 : std_logic;
signal measured_delay_tr_9 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_100mhz_0 : std_logic;
signal \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\ : std_logic;
signal red_c_g : std_logic;

signal reset_wire : std_logic;
signal start_stop_wire : std_logic;
signal il_max_comp2_wire : std_logic;
signal pwm_output_wire : std_logic;
signal il_max_comp1_wire : std_logic;
signal s2_phy_wire : std_logic;
signal delay_hc_input_wire : std_logic;
signal delay_tr_input_wire : std_logic;
signal il_min_comp2_wire : std_logic;
signal s1_phy_wire : std_logic;
signal s4_phy_wire : std_logic;
signal il_min_comp1_wire : std_logic;
signal s3_phy_wire : std_logic;
signal rgb_b_wire : std_logic;
signal rgb_g_wire : std_logic;
signal rgb_r_wire : std_logic;
signal \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);

begin
    reset_wire <= reset;
    start_stop_wire <= start_stop;
    il_max_comp2_wire <= il_max_comp2;
    pwm_output <= pwm_output_wire;
    il_max_comp1_wire <= il_max_comp1;
    s2_phy <= s2_phy_wire;
    delay_hc_input_wire <= delay_hc_input;
    delay_tr_input_wire <= delay_tr_input;
    il_min_comp2_wire <= il_min_comp2;
    s1_phy <= s1_phy_wire;
    s4_phy <= s4_phy_wire;
    il_min_comp1_wire <= il_min_comp1;
    s3_phy <= s3_phy_wire;
    rgb_b <= rgb_b_wire;
    rgb_g <= rgb_g_wire;
    rgb_r <= rgb_r_wire;
    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_A_wire\ <= '0'&\N__18887\&\N__18890\&\N__18888\&\N__18891\&\N__18889\&\N__19120\&\N__19100\&\N__19064\&\N__20811\&\N__19139\&\N__18846\&\N__19002\&\N__18970\&\N__19015\&\N__18982\;
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__28855\&\N__28852\&'0'&'0'&'0'&\N__28850\&\N__28854\&\N__28851\&\N__28853\;
    \pwm_generator_inst.un2_threshold_acc_1_25\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(25);
    \pwm_generator_inst.un2_threshold_acc_1_24\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(24);
    \pwm_generator_inst.un2_threshold_acc_1_23\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(23);
    \pwm_generator_inst.un2_threshold_acc_1_22\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(22);
    \pwm_generator_inst.un2_threshold_acc_1_21\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(21);
    \pwm_generator_inst.un2_threshold_acc_1_20\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(20);
    \pwm_generator_inst.un2_threshold_acc_1_19\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(19);
    \pwm_generator_inst.un2_threshold_acc_1_18\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(18);
    \pwm_generator_inst.un2_threshold_acc_1_17\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(17);
    \pwm_generator_inst.un2_threshold_acc_1_16\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_acc_1_15\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.O_14\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.O_13\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.O_12\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un3_threshold_acc\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.O_10\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.O_9\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.O_8\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.O_7\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.O_6\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.O_5\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.O_4\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.O_3\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.O_2\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.O_1\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.O_0\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_A_wire\ <= '0'&\N__18950\&\N__18943\&\N__18948\&\N__18942\&\N__18949\&\N__18941\&\N__18951\&\N__18938\&\N__18944\&\N__18937\&\N__18945\&\N__18939\&\N__18946\&\N__18940\&\N__18947\;
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__28823\&\N__28820\&'0'&'0'&'0'&\N__28818\&\N__28822\&\N__28819\&\N__28821\;
    \pwm_generator_inst.un2_threshold_acc_2_1_16\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_acc_2_1_15\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.un2_threshold_acc_2_14\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.un2_threshold_acc_2_13\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.un2_threshold_acc_2_12\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un2_threshold_acc_2_11\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.un2_threshold_acc_2_10\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.un2_threshold_acc_2_9\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.un2_threshold_acc_2_8\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.un2_threshold_acc_2_7\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.un2_threshold_acc_2_6\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.un2_threshold_acc_2_5\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.un2_threshold_acc_2_4\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.un2_threshold_acc_2_3\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.un2_threshold_acc_2_2\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.un2_threshold_acc_2_1\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.un2_threshold_acc_2_0\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(0);

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__31943\,
            RESETB => \N__40529\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => clk_100mhz_0
        );

    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__28856\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__28849\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__28731\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__28817\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\
        );

    \reset_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__48351\,
            GLOBALBUFFEROUTPUT => red_c_g
        );

    \reset_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48353\,
            DIN => \N__48352\,
            DOUT => \N__48351\,
            PACKAGEPIN => reset_wire
        );

    \reset_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48353\,
            PADOUT => \N__48352\,
            PADIN => \N__48351\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \start_stop_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48342\,
            DIN => \N__48341\,
            DOUT => \N__48340\,
            PACKAGEPIN => start_stop_wire
        );

    \start_stop_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48342\,
            PADOUT => \N__48341\,
            PADIN => \N__48340\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => start_stop_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48333\,
            DIN => \N__48332\,
            DOUT => \N__48331\,
            PACKAGEPIN => il_max_comp2_wire
        );

    \il_max_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48333\,
            PADOUT => \N__48332\,
            PADIN => \N__48331\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48324\,
            DIN => \N__48323\,
            DOUT => \N__48322\,
            PACKAGEPIN => pwm_output_wire
        );

    \pwm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48324\,
            PADOUT => \N__48323\,
            PADIN => \N__48322\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23270\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48315\,
            DIN => \N__48314\,
            DOUT => \N__48313\,
            PACKAGEPIN => il_max_comp1_wire
        );

    \il_max_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48315\,
            PADOUT => \N__48314\,
            PADIN => \N__48313\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s2_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48306\,
            DIN => \N__48305\,
            DOUT => \N__48304\,
            PACKAGEPIN => s2_phy_wire
        );

    \s2_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48306\,
            PADOUT => \N__48305\,
            PADIN => \N__48304\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__33443\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_hc_input_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48297\,
            DIN => \N__48296\,
            DOUT => \N__48295\,
            PACKAGEPIN => delay_hc_input_wire
        );

    \delay_hc_input_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48297\,
            PADOUT => \N__48296\,
            PADIN => \N__48295\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_hc_input_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_tr_input_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48288\,
            DIN => \N__48287\,
            DOUT => \N__48286\,
            PACKAGEPIN => delay_tr_input_wire
        );

    \delay_tr_input_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48288\,
            PADOUT => \N__48287\,
            PADIN => \N__48286\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_tr_input_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48279\,
            DIN => \N__48278\,
            DOUT => \N__48277\,
            PACKAGEPIN => il_min_comp2_wire
        );

    \il_min_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48279\,
            PADOUT => \N__48278\,
            PADIN => \N__48277\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s1_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48270\,
            DIN => \N__48269\,
            DOUT => \N__48268\,
            PACKAGEPIN => s1_phy_wire
        );

    \s1_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48270\,
            PADOUT => \N__48269\,
            PADIN => \N__48268\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__32888\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s4_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48261\,
            DIN => \N__48260\,
            DOUT => \N__48259\,
            PACKAGEPIN => s4_phy_wire
        );

    \s4_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48261\,
            PADOUT => \N__48260\,
            PADIN => \N__48259\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__28436\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48252\,
            DIN => \N__48251\,
            DOUT => \N__48250\,
            PACKAGEPIN => il_min_comp1_wire
        );

    \il_min_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48252\,
            PADOUT => \N__48251\,
            PADIN => \N__48250\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s3_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48243\,
            DIN => \N__48242\,
            DOUT => \N__48241\,
            PACKAGEPIN => s3_phy_wire
        );

    \s3_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48243\,
            PADOUT => \N__48242\,
            PADIN => \N__48241\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__31913\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__11547\ : InMux
    port map (
            O => \N__48224\,
            I => \N__48221\
        );

    \I__11546\ : LocalMux
    port map (
            O => \N__48221\,
            I => \N__48218\
        );

    \I__11545\ : Odrv4
    port map (
            O => \N__48218\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9\
        );

    \I__11544\ : InMux
    port map (
            O => \N__48215\,
            I => \N__48211\
        );

    \I__11543\ : InMux
    port map (
            O => \N__48214\,
            I => \N__48208\
        );

    \I__11542\ : LocalMux
    port map (
            O => \N__48211\,
            I => \N__48205\
        );

    \I__11541\ : LocalMux
    port map (
            O => \N__48208\,
            I => \N__48202\
        );

    \I__11540\ : Odrv4
    port map (
            O => \N__48205\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__11539\ : Odrv4
    port map (
            O => \N__48202\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__11538\ : CascadeMux
    port map (
            O => \N__48197\,
            I => \N__48192\
        );

    \I__11537\ : CascadeMux
    port map (
            O => \N__48196\,
            I => \N__48189\
        );

    \I__11536\ : CascadeMux
    port map (
            O => \N__48195\,
            I => \N__48186\
        );

    \I__11535\ : InMux
    port map (
            O => \N__48192\,
            I => \N__48164\
        );

    \I__11534\ : InMux
    port map (
            O => \N__48189\,
            I => \N__48164\
        );

    \I__11533\ : InMux
    port map (
            O => \N__48186\,
            I => \N__48164\
        );

    \I__11532\ : InMux
    port map (
            O => \N__48185\,
            I => \N__48164\
        );

    \I__11531\ : InMux
    port map (
            O => \N__48184\,
            I => \N__48159\
        );

    \I__11530\ : InMux
    port map (
            O => \N__48183\,
            I => \N__48159\
        );

    \I__11529\ : CascadeMux
    port map (
            O => \N__48182\,
            I => \N__48150\
        );

    \I__11528\ : CascadeMux
    port map (
            O => \N__48181\,
            I => \N__48146\
        );

    \I__11527\ : CascadeMux
    port map (
            O => \N__48180\,
            I => \N__48142\
        );

    \I__11526\ : CascadeMux
    port map (
            O => \N__48179\,
            I => \N__48139\
        );

    \I__11525\ : InMux
    port map (
            O => \N__48178\,
            I => \N__48126\
        );

    \I__11524\ : InMux
    port map (
            O => \N__48177\,
            I => \N__48126\
        );

    \I__11523\ : InMux
    port map (
            O => \N__48176\,
            I => \N__48126\
        );

    \I__11522\ : InMux
    port map (
            O => \N__48175\,
            I => \N__48126\
        );

    \I__11521\ : InMux
    port map (
            O => \N__48174\,
            I => \N__48126\
        );

    \I__11520\ : InMux
    port map (
            O => \N__48173\,
            I => \N__48126\
        );

    \I__11519\ : LocalMux
    port map (
            O => \N__48164\,
            I => \N__48121\
        );

    \I__11518\ : LocalMux
    port map (
            O => \N__48159\,
            I => \N__48121\
        );

    \I__11517\ : InMux
    port map (
            O => \N__48158\,
            I => \N__48118\
        );

    \I__11516\ : InMux
    port map (
            O => \N__48157\,
            I => \N__48115\
        );

    \I__11515\ : InMux
    port map (
            O => \N__48156\,
            I => \N__48110\
        );

    \I__11514\ : InMux
    port map (
            O => \N__48155\,
            I => \N__48110\
        );

    \I__11513\ : InMux
    port map (
            O => \N__48154\,
            I => \N__48093\
        );

    \I__11512\ : InMux
    port map (
            O => \N__48153\,
            I => \N__48093\
        );

    \I__11511\ : InMux
    port map (
            O => \N__48150\,
            I => \N__48093\
        );

    \I__11510\ : InMux
    port map (
            O => \N__48149\,
            I => \N__48093\
        );

    \I__11509\ : InMux
    port map (
            O => \N__48146\,
            I => \N__48093\
        );

    \I__11508\ : InMux
    port map (
            O => \N__48145\,
            I => \N__48093\
        );

    \I__11507\ : InMux
    port map (
            O => \N__48142\,
            I => \N__48093\
        );

    \I__11506\ : InMux
    port map (
            O => \N__48139\,
            I => \N__48093\
        );

    \I__11505\ : LocalMux
    port map (
            O => \N__48126\,
            I => \N__48088\
        );

    \I__11504\ : Span4Mux_v
    port map (
            O => \N__48121\,
            I => \N__48088\
        );

    \I__11503\ : LocalMux
    port map (
            O => \N__48118\,
            I => \N__48085\
        );

    \I__11502\ : LocalMux
    port map (
            O => \N__48115\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__11501\ : LocalMux
    port map (
            O => \N__48110\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__11500\ : LocalMux
    port map (
            O => \N__48093\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__11499\ : Odrv4
    port map (
            O => \N__48088\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__11498\ : Odrv4
    port map (
            O => \N__48085\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__11497\ : CascadeMux
    port map (
            O => \N__48074\,
            I => \N__48068\
        );

    \I__11496\ : CascadeMux
    port map (
            O => \N__48073\,
            I => \N__48056\
        );

    \I__11495\ : CascadeMux
    port map (
            O => \N__48072\,
            I => \N__48053\
        );

    \I__11494\ : CascadeMux
    port map (
            O => \N__48071\,
            I => \N__48050\
        );

    \I__11493\ : InMux
    port map (
            O => \N__48068\,
            I => \N__48042\
        );

    \I__11492\ : InMux
    port map (
            O => \N__48067\,
            I => \N__48042\
        );

    \I__11491\ : CascadeMux
    port map (
            O => \N__48066\,
            I => \N__48039\
        );

    \I__11490\ : CascadeMux
    port map (
            O => \N__48065\,
            I => \N__48036\
        );

    \I__11489\ : CascadeMux
    port map (
            O => \N__48064\,
            I => \N__48033\
        );

    \I__11488\ : CascadeMux
    port map (
            O => \N__48063\,
            I => \N__48030\
        );

    \I__11487\ : InMux
    port map (
            O => \N__48062\,
            I => \N__48015\
        );

    \I__11486\ : InMux
    port map (
            O => \N__48061\,
            I => \N__48015\
        );

    \I__11485\ : InMux
    port map (
            O => \N__48060\,
            I => \N__48015\
        );

    \I__11484\ : InMux
    port map (
            O => \N__48059\,
            I => \N__48015\
        );

    \I__11483\ : InMux
    port map (
            O => \N__48056\,
            I => \N__48002\
        );

    \I__11482\ : InMux
    port map (
            O => \N__48053\,
            I => \N__48002\
        );

    \I__11481\ : InMux
    port map (
            O => \N__48050\,
            I => \N__48002\
        );

    \I__11480\ : InMux
    port map (
            O => \N__48049\,
            I => \N__48002\
        );

    \I__11479\ : InMux
    port map (
            O => \N__48048\,
            I => \N__48002\
        );

    \I__11478\ : InMux
    port map (
            O => \N__48047\,
            I => \N__48002\
        );

    \I__11477\ : LocalMux
    port map (
            O => \N__48042\,
            I => \N__47999\
        );

    \I__11476\ : InMux
    port map (
            O => \N__48039\,
            I => \N__47988\
        );

    \I__11475\ : InMux
    port map (
            O => \N__48036\,
            I => \N__47988\
        );

    \I__11474\ : InMux
    port map (
            O => \N__48033\,
            I => \N__47988\
        );

    \I__11473\ : InMux
    port map (
            O => \N__48030\,
            I => \N__47988\
        );

    \I__11472\ : InMux
    port map (
            O => \N__48029\,
            I => \N__47983\
        );

    \I__11471\ : InMux
    port map (
            O => \N__48028\,
            I => \N__47983\
        );

    \I__11470\ : InMux
    port map (
            O => \N__48027\,
            I => \N__47974\
        );

    \I__11469\ : InMux
    port map (
            O => \N__48026\,
            I => \N__47974\
        );

    \I__11468\ : InMux
    port map (
            O => \N__48025\,
            I => \N__47974\
        );

    \I__11467\ : InMux
    port map (
            O => \N__48024\,
            I => \N__47974\
        );

    \I__11466\ : LocalMux
    port map (
            O => \N__48015\,
            I => \N__47969\
        );

    \I__11465\ : LocalMux
    port map (
            O => \N__48002\,
            I => \N__47969\
        );

    \I__11464\ : Span4Mux_h
    port map (
            O => \N__47999\,
            I => \N__47966\
        );

    \I__11463\ : InMux
    port map (
            O => \N__47998\,
            I => \N__47961\
        );

    \I__11462\ : InMux
    port map (
            O => \N__47997\,
            I => \N__47961\
        );

    \I__11461\ : LocalMux
    port map (
            O => \N__47988\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__11460\ : LocalMux
    port map (
            O => \N__47983\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__11459\ : LocalMux
    port map (
            O => \N__47974\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__11458\ : Odrv4
    port map (
            O => \N__47969\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__11457\ : Odrv4
    port map (
            O => \N__47966\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__11456\ : LocalMux
    port map (
            O => \N__47961\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__11455\ : CascadeMux
    port map (
            O => \N__47948\,
            I => \N__47943\
        );

    \I__11454\ : CascadeMux
    port map (
            O => \N__47947\,
            I => \N__47937\
        );

    \I__11453\ : CascadeMux
    port map (
            O => \N__47946\,
            I => \N__47934\
        );

    \I__11452\ : InMux
    port map (
            O => \N__47943\,
            I => \N__47930\
        );

    \I__11451\ : InMux
    port map (
            O => \N__47942\,
            I => \N__47923\
        );

    \I__11450\ : InMux
    port map (
            O => \N__47941\,
            I => \N__47923\
        );

    \I__11449\ : InMux
    port map (
            O => \N__47940\,
            I => \N__47923\
        );

    \I__11448\ : InMux
    port map (
            O => \N__47937\,
            I => \N__47916\
        );

    \I__11447\ : InMux
    port map (
            O => \N__47934\,
            I => \N__47916\
        );

    \I__11446\ : InMux
    port map (
            O => \N__47933\,
            I => \N__47916\
        );

    \I__11445\ : LocalMux
    port map (
            O => \N__47930\,
            I => \N__47903\
        );

    \I__11444\ : LocalMux
    port map (
            O => \N__47923\,
            I => \N__47903\
        );

    \I__11443\ : LocalMux
    port map (
            O => \N__47916\,
            I => \N__47903\
        );

    \I__11442\ : InMux
    port map (
            O => \N__47915\,
            I => \N__47898\
        );

    \I__11441\ : InMux
    port map (
            O => \N__47914\,
            I => \N__47898\
        );

    \I__11440\ : CascadeMux
    port map (
            O => \N__47913\,
            I => \N__47895\
        );

    \I__11439\ : InMux
    port map (
            O => \N__47912\,
            I => \N__47879\
        );

    \I__11438\ : InMux
    port map (
            O => \N__47911\,
            I => \N__47879\
        );

    \I__11437\ : InMux
    port map (
            O => \N__47910\,
            I => \N__47879\
        );

    \I__11436\ : Span4Mux_v
    port map (
            O => \N__47903\,
            I => \N__47874\
        );

    \I__11435\ : LocalMux
    port map (
            O => \N__47898\,
            I => \N__47874\
        );

    \I__11434\ : InMux
    port map (
            O => \N__47895\,
            I => \N__47867\
        );

    \I__11433\ : InMux
    port map (
            O => \N__47894\,
            I => \N__47867\
        );

    \I__11432\ : InMux
    port map (
            O => \N__47893\,
            I => \N__47850\
        );

    \I__11431\ : InMux
    port map (
            O => \N__47892\,
            I => \N__47850\
        );

    \I__11430\ : InMux
    port map (
            O => \N__47891\,
            I => \N__47850\
        );

    \I__11429\ : InMux
    port map (
            O => \N__47890\,
            I => \N__47850\
        );

    \I__11428\ : InMux
    port map (
            O => \N__47889\,
            I => \N__47850\
        );

    \I__11427\ : InMux
    port map (
            O => \N__47888\,
            I => \N__47850\
        );

    \I__11426\ : InMux
    port map (
            O => \N__47887\,
            I => \N__47850\
        );

    \I__11425\ : InMux
    port map (
            O => \N__47886\,
            I => \N__47850\
        );

    \I__11424\ : LocalMux
    port map (
            O => \N__47879\,
            I => \N__47845\
        );

    \I__11423\ : Span4Mux_h
    port map (
            O => \N__47874\,
            I => \N__47845\
        );

    \I__11422\ : InMux
    port map (
            O => \N__47873\,
            I => \N__47840\
        );

    \I__11421\ : InMux
    port map (
            O => \N__47872\,
            I => \N__47840\
        );

    \I__11420\ : LocalMux
    port map (
            O => \N__47867\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__11419\ : LocalMux
    port map (
            O => \N__47850\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__11418\ : Odrv4
    port map (
            O => \N__47845\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__11417\ : LocalMux
    port map (
            O => \N__47840\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__11416\ : InMux
    port map (
            O => \N__47831\,
            I => \N__47828\
        );

    \I__11415\ : LocalMux
    port map (
            O => \N__47828\,
            I => \N__47825\
        );

    \I__11414\ : Span4Mux_v
    port map (
            O => \N__47825\,
            I => \N__47821\
        );

    \I__11413\ : InMux
    port map (
            O => \N__47824\,
            I => \N__47818\
        );

    \I__11412\ : Sp12to4
    port map (
            O => \N__47821\,
            I => \N__47813\
        );

    \I__11411\ : LocalMux
    port map (
            O => \N__47818\,
            I => \N__47813\
        );

    \I__11410\ : Odrv12
    port map (
            O => \N__47813\,
            I => \phase_controller_inst1.stoper_tr.N_21\
        );

    \I__11409\ : InMux
    port map (
            O => \N__47810\,
            I => \N__47807\
        );

    \I__11408\ : LocalMux
    port map (
            O => \N__47807\,
            I => \N__47803\
        );

    \I__11407\ : CascadeMux
    port map (
            O => \N__47806\,
            I => \N__47800\
        );

    \I__11406\ : Span4Mux_h
    port map (
            O => \N__47803\,
            I => \N__47797\
        );

    \I__11405\ : InMux
    port map (
            O => \N__47800\,
            I => \N__47794\
        );

    \I__11404\ : Span4Mux_v
    port map (
            O => \N__47797\,
            I => \N__47791\
        );

    \I__11403\ : LocalMux
    port map (
            O => \N__47794\,
            I => \N__47788\
        );

    \I__11402\ : Odrv4
    port map (
            O => \N__47791\,
            I => \delay_measurement_inst.N_271_1\
        );

    \I__11401\ : Odrv4
    port map (
            O => \N__47788\,
            I => \delay_measurement_inst.N_271_1\
        );

    \I__11400\ : InMux
    port map (
            O => \N__47783\,
            I => \N__47776\
        );

    \I__11399\ : InMux
    port map (
            O => \N__47782\,
            I => \N__47773\
        );

    \I__11398\ : InMux
    port map (
            O => \N__47781\,
            I => \N__47770\
        );

    \I__11397\ : InMux
    port map (
            O => \N__47780\,
            I => \N__47767\
        );

    \I__11396\ : InMux
    port map (
            O => \N__47779\,
            I => \N__47764\
        );

    \I__11395\ : LocalMux
    port map (
            O => \N__47776\,
            I => \N__47761\
        );

    \I__11394\ : LocalMux
    port map (
            O => \N__47773\,
            I => \N__47756\
        );

    \I__11393\ : LocalMux
    port map (
            O => \N__47770\,
            I => \N__47756\
        );

    \I__11392\ : LocalMux
    port map (
            O => \N__47767\,
            I => \N__47753\
        );

    \I__11391\ : LocalMux
    port map (
            O => \N__47764\,
            I => \N__47750\
        );

    \I__11390\ : Span4Mux_v
    port map (
            O => \N__47761\,
            I => \N__47745\
        );

    \I__11389\ : Span4Mux_v
    port map (
            O => \N__47756\,
            I => \N__47745\
        );

    \I__11388\ : Span4Mux_h
    port map (
            O => \N__47753\,
            I => \N__47742\
        );

    \I__11387\ : Odrv12
    port map (
            O => \N__47750\,
            I => \delay_measurement_inst.elapsed_time_tr_14\
        );

    \I__11386\ : Odrv4
    port map (
            O => \N__47745\,
            I => \delay_measurement_inst.elapsed_time_tr_14\
        );

    \I__11385\ : Odrv4
    port map (
            O => \N__47742\,
            I => \delay_measurement_inst.elapsed_time_tr_14\
        );

    \I__11384\ : InMux
    port map (
            O => \N__47735\,
            I => \N__47732\
        );

    \I__11383\ : LocalMux
    port map (
            O => \N__47732\,
            I => \N__47729\
        );

    \I__11382\ : Span4Mux_v
    port map (
            O => \N__47729\,
            I => \N__47726\
        );

    \I__11381\ : Span4Mux_v
    port map (
            O => \N__47726\,
            I => \N__47720\
        );

    \I__11380\ : InMux
    port map (
            O => \N__47725\,
            I => \N__47713\
        );

    \I__11379\ : InMux
    port map (
            O => \N__47724\,
            I => \N__47713\
        );

    \I__11378\ : InMux
    port map (
            O => \N__47723\,
            I => \N__47713\
        );

    \I__11377\ : Odrv4
    port map (
            O => \N__47720\,
            I => \delay_measurement_inst.N_265_i\
        );

    \I__11376\ : LocalMux
    port map (
            O => \N__47713\,
            I => \delay_measurement_inst.N_265_i\
        );

    \I__11375\ : InMux
    port map (
            O => \N__47708\,
            I => \N__47701\
        );

    \I__11374\ : InMux
    port map (
            O => \N__47707\,
            I => \N__47701\
        );

    \I__11373\ : InMux
    port map (
            O => \N__47706\,
            I => \N__47698\
        );

    \I__11372\ : LocalMux
    port map (
            O => \N__47701\,
            I => \N__47695\
        );

    \I__11371\ : LocalMux
    port map (
            O => \N__47698\,
            I => \N__47691\
        );

    \I__11370\ : Span4Mux_h
    port map (
            O => \N__47695\,
            I => \N__47688\
        );

    \I__11369\ : CascadeMux
    port map (
            O => \N__47694\,
            I => \N__47685\
        );

    \I__11368\ : Span4Mux_h
    port map (
            O => \N__47691\,
            I => \N__47681\
        );

    \I__11367\ : Span4Mux_h
    port map (
            O => \N__47688\,
            I => \N__47678\
        );

    \I__11366\ : InMux
    port map (
            O => \N__47685\,
            I => \N__47673\
        );

    \I__11365\ : InMux
    port map (
            O => \N__47684\,
            I => \N__47673\
        );

    \I__11364\ : Odrv4
    port map (
            O => \N__47681\,
            I => measured_delay_tr_14
        );

    \I__11363\ : Odrv4
    port map (
            O => \N__47678\,
            I => measured_delay_tr_14
        );

    \I__11362\ : LocalMux
    port map (
            O => \N__47673\,
            I => measured_delay_tr_14
        );

    \I__11361\ : InMux
    port map (
            O => \N__47666\,
            I => \N__47660\
        );

    \I__11360\ : InMux
    port map (
            O => \N__47665\,
            I => \N__47657\
        );

    \I__11359\ : InMux
    port map (
            O => \N__47664\,
            I => \N__47652\
        );

    \I__11358\ : InMux
    port map (
            O => \N__47663\,
            I => \N__47652\
        );

    \I__11357\ : LocalMux
    port map (
            O => \N__47660\,
            I => \N__47649\
        );

    \I__11356\ : LocalMux
    port map (
            O => \N__47657\,
            I => \phase_controller_slave.hc_time_passed\
        );

    \I__11355\ : LocalMux
    port map (
            O => \N__47652\,
            I => \phase_controller_slave.hc_time_passed\
        );

    \I__11354\ : Odrv12
    port map (
            O => \N__47649\,
            I => \phase_controller_slave.hc_time_passed\
        );

    \I__11353\ : InMux
    port map (
            O => \N__47642\,
            I => \N__47638\
        );

    \I__11352\ : CascadeMux
    port map (
            O => \N__47641\,
            I => \N__47634\
        );

    \I__11351\ : LocalMux
    port map (
            O => \N__47638\,
            I => \N__47631\
        );

    \I__11350\ : InMux
    port map (
            O => \N__47637\,
            I => \N__47628\
        );

    \I__11349\ : InMux
    port map (
            O => \N__47634\,
            I => \N__47625\
        );

    \I__11348\ : Span4Mux_h
    port map (
            O => \N__47631\,
            I => \N__47622\
        );

    \I__11347\ : LocalMux
    port map (
            O => \N__47628\,
            I => \phase_controller_slave.stateZ0Z_2\
        );

    \I__11346\ : LocalMux
    port map (
            O => \N__47625\,
            I => \phase_controller_slave.stateZ0Z_2\
        );

    \I__11345\ : Odrv4
    port map (
            O => \N__47622\,
            I => \phase_controller_slave.stateZ0Z_2\
        );

    \I__11344\ : InMux
    port map (
            O => \N__47615\,
            I => \N__47612\
        );

    \I__11343\ : LocalMux
    port map (
            O => \N__47612\,
            I => \N__47609\
        );

    \I__11342\ : Odrv12
    port map (
            O => \N__47609\,
            I => \phase_controller_slave.N_211\
        );

    \I__11341\ : InMux
    port map (
            O => \N__47606\,
            I => \N__47599\
        );

    \I__11340\ : InMux
    port map (
            O => \N__47605\,
            I => \N__47599\
        );

    \I__11339\ : InMux
    port map (
            O => \N__47604\,
            I => \N__47590\
        );

    \I__11338\ : LocalMux
    port map (
            O => \N__47599\,
            I => \N__47587\
        );

    \I__11337\ : InMux
    port map (
            O => \N__47598\,
            I => \N__47578\
        );

    \I__11336\ : InMux
    port map (
            O => \N__47597\,
            I => \N__47578\
        );

    \I__11335\ : InMux
    port map (
            O => \N__47596\,
            I => \N__47578\
        );

    \I__11334\ : InMux
    port map (
            O => \N__47595\,
            I => \N__47578\
        );

    \I__11333\ : InMux
    port map (
            O => \N__47594\,
            I => \N__47573\
        );

    \I__11332\ : InMux
    port map (
            O => \N__47593\,
            I => \N__47573\
        );

    \I__11331\ : LocalMux
    port map (
            O => \N__47590\,
            I => \N__47570\
        );

    \I__11330\ : Span4Mux_v
    port map (
            O => \N__47587\,
            I => \N__47567\
        );

    \I__11329\ : LocalMux
    port map (
            O => \N__47578\,
            I => \N__47564\
        );

    \I__11328\ : LocalMux
    port map (
            O => \N__47573\,
            I => \N__47561\
        );

    \I__11327\ : Span4Mux_v
    port map (
            O => \N__47570\,
            I => \N__47558\
        );

    \I__11326\ : Span4Mux_h
    port map (
            O => \N__47567\,
            I => \N__47555\
        );

    \I__11325\ : Span4Mux_v
    port map (
            O => \N__47564\,
            I => \N__47552\
        );

    \I__11324\ : Span4Mux_v
    port map (
            O => \N__47561\,
            I => \N__47547\
        );

    \I__11323\ : Span4Mux_h
    port map (
            O => \N__47558\,
            I => \N__47547\
        );

    \I__11322\ : Odrv4
    port map (
            O => \N__47555\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13\
        );

    \I__11321\ : Odrv4
    port map (
            O => \N__47552\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13\
        );

    \I__11320\ : Odrv4
    port map (
            O => \N__47547\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13\
        );

    \I__11319\ : InMux
    port map (
            O => \N__47540\,
            I => \N__47531\
        );

    \I__11318\ : InMux
    port map (
            O => \N__47539\,
            I => \N__47527\
        );

    \I__11317\ : InMux
    port map (
            O => \N__47538\,
            I => \N__47524\
        );

    \I__11316\ : InMux
    port map (
            O => \N__47537\,
            I => \N__47521\
        );

    \I__11315\ : InMux
    port map (
            O => \N__47536\,
            I => \N__47513\
        );

    \I__11314\ : InMux
    port map (
            O => \N__47535\,
            I => \N__47513\
        );

    \I__11313\ : InMux
    port map (
            O => \N__47534\,
            I => \N__47513\
        );

    \I__11312\ : LocalMux
    port map (
            O => \N__47531\,
            I => \N__47510\
        );

    \I__11311\ : InMux
    port map (
            O => \N__47530\,
            I => \N__47507\
        );

    \I__11310\ : LocalMux
    port map (
            O => \N__47527\,
            I => \N__47502\
        );

    \I__11309\ : LocalMux
    port map (
            O => \N__47524\,
            I => \N__47502\
        );

    \I__11308\ : LocalMux
    port map (
            O => \N__47521\,
            I => \N__47499\
        );

    \I__11307\ : InMux
    port map (
            O => \N__47520\,
            I => \N__47496\
        );

    \I__11306\ : LocalMux
    port map (
            O => \N__47513\,
            I => \N__47493\
        );

    \I__11305\ : Span4Mux_h
    port map (
            O => \N__47510\,
            I => \N__47488\
        );

    \I__11304\ : LocalMux
    port map (
            O => \N__47507\,
            I => \N__47488\
        );

    \I__11303\ : Span4Mux_v
    port map (
            O => \N__47502\,
            I => \N__47484\
        );

    \I__11302\ : Span4Mux_h
    port map (
            O => \N__47499\,
            I => \N__47481\
        );

    \I__11301\ : LocalMux
    port map (
            O => \N__47496\,
            I => \N__47478\
        );

    \I__11300\ : Span4Mux_v
    port map (
            O => \N__47493\,
            I => \N__47475\
        );

    \I__11299\ : Span4Mux_v
    port map (
            O => \N__47488\,
            I => \N__47472\
        );

    \I__11298\ : InMux
    port map (
            O => \N__47487\,
            I => \N__47469\
        );

    \I__11297\ : Span4Mux_v
    port map (
            O => \N__47484\,
            I => \N__47466\
        );

    \I__11296\ : Span4Mux_v
    port map (
            O => \N__47481\,
            I => \N__47463\
        );

    \I__11295\ : Span4Mux_h
    port map (
            O => \N__47478\,
            I => \N__47456\
        );

    \I__11294\ : Span4Mux_v
    port map (
            O => \N__47475\,
            I => \N__47456\
        );

    \I__11293\ : Span4Mux_v
    port map (
            O => \N__47472\,
            I => \N__47456\
        );

    \I__11292\ : LocalMux
    port map (
            O => \N__47469\,
            I => measured_delay_tr_15
        );

    \I__11291\ : Odrv4
    port map (
            O => \N__47466\,
            I => measured_delay_tr_15
        );

    \I__11290\ : Odrv4
    port map (
            O => \N__47463\,
            I => measured_delay_tr_15
        );

    \I__11289\ : Odrv4
    port map (
            O => \N__47456\,
            I => measured_delay_tr_15
        );

    \I__11288\ : CascadeMux
    port map (
            O => \N__47447\,
            I => \N__47444\
        );

    \I__11287\ : InMux
    port map (
            O => \N__47444\,
            I => \N__47439\
        );

    \I__11286\ : InMux
    port map (
            O => \N__47443\,
            I => \N__47436\
        );

    \I__11285\ : CascadeMux
    port map (
            O => \N__47442\,
            I => \N__47432\
        );

    \I__11284\ : LocalMux
    port map (
            O => \N__47439\,
            I => \N__47429\
        );

    \I__11283\ : LocalMux
    port map (
            O => \N__47436\,
            I => \N__47426\
        );

    \I__11282\ : InMux
    port map (
            O => \N__47435\,
            I => \N__47421\
        );

    \I__11281\ : InMux
    port map (
            O => \N__47432\,
            I => \N__47421\
        );

    \I__11280\ : Span4Mux_v
    port map (
            O => \N__47429\,
            I => \N__47418\
        );

    \I__11279\ : Span4Mux_h
    port map (
            O => \N__47426\,
            I => \N__47413\
        );

    \I__11278\ : LocalMux
    port map (
            O => \N__47421\,
            I => \N__47413\
        );

    \I__11277\ : Span4Mux_h
    port map (
            O => \N__47418\,
            I => \N__47410\
        );

    \I__11276\ : Span4Mux_v
    port map (
            O => \N__47413\,
            I => \N__47407\
        );

    \I__11275\ : Odrv4
    port map (
            O => \N__47410\,
            I => measured_delay_tr_9
        );

    \I__11274\ : Odrv4
    port map (
            O => \N__47407\,
            I => measured_delay_tr_9
        );

    \I__11273\ : InMux
    port map (
            O => \N__47402\,
            I => \N__47397\
        );

    \I__11272\ : InMux
    port map (
            O => \N__47401\,
            I => \N__47392\
        );

    \I__11271\ : InMux
    port map (
            O => \N__47400\,
            I => \N__47392\
        );

    \I__11270\ : LocalMux
    port map (
            O => \N__47397\,
            I => \N__47387\
        );

    \I__11269\ : LocalMux
    port map (
            O => \N__47392\,
            I => \N__47384\
        );

    \I__11268\ : InMux
    port map (
            O => \N__47391\,
            I => \N__47379\
        );

    \I__11267\ : InMux
    port map (
            O => \N__47390\,
            I => \N__47379\
        );

    \I__11266\ : Span4Mux_v
    port map (
            O => \N__47387\,
            I => \N__47376\
        );

    \I__11265\ : Span4Mux_v
    port map (
            O => \N__47384\,
            I => \N__47371\
        );

    \I__11264\ : LocalMux
    port map (
            O => \N__47379\,
            I => \N__47371\
        );

    \I__11263\ : Span4Mux_h
    port map (
            O => \N__47376\,
            I => \N__47366\
        );

    \I__11262\ : Span4Mux_h
    port map (
            O => \N__47371\,
            I => \N__47366\
        );

    \I__11261\ : Odrv4
    port map (
            O => \N__47366\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0Z0Z_6\
        );

    \I__11260\ : CascadeMux
    port map (
            O => \N__47363\,
            I => \N__47360\
        );

    \I__11259\ : InMux
    port map (
            O => \N__47360\,
            I => \N__47357\
        );

    \I__11258\ : LocalMux
    port map (
            O => \N__47357\,
            I => \N__47354\
        );

    \I__11257\ : Odrv12
    port map (
            O => \N__47354\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\
        );

    \I__11256\ : ClkMux
    port map (
            O => \N__47351\,
            I => \N__46862\
        );

    \I__11255\ : ClkMux
    port map (
            O => \N__47350\,
            I => \N__46862\
        );

    \I__11254\ : ClkMux
    port map (
            O => \N__47349\,
            I => \N__46862\
        );

    \I__11253\ : ClkMux
    port map (
            O => \N__47348\,
            I => \N__46862\
        );

    \I__11252\ : ClkMux
    port map (
            O => \N__47347\,
            I => \N__46862\
        );

    \I__11251\ : ClkMux
    port map (
            O => \N__47346\,
            I => \N__46862\
        );

    \I__11250\ : ClkMux
    port map (
            O => \N__47345\,
            I => \N__46862\
        );

    \I__11249\ : ClkMux
    port map (
            O => \N__47344\,
            I => \N__46862\
        );

    \I__11248\ : ClkMux
    port map (
            O => \N__47343\,
            I => \N__46862\
        );

    \I__11247\ : ClkMux
    port map (
            O => \N__47342\,
            I => \N__46862\
        );

    \I__11246\ : ClkMux
    port map (
            O => \N__47341\,
            I => \N__46862\
        );

    \I__11245\ : ClkMux
    port map (
            O => \N__47340\,
            I => \N__46862\
        );

    \I__11244\ : ClkMux
    port map (
            O => \N__47339\,
            I => \N__46862\
        );

    \I__11243\ : ClkMux
    port map (
            O => \N__47338\,
            I => \N__46862\
        );

    \I__11242\ : ClkMux
    port map (
            O => \N__47337\,
            I => \N__46862\
        );

    \I__11241\ : ClkMux
    port map (
            O => \N__47336\,
            I => \N__46862\
        );

    \I__11240\ : ClkMux
    port map (
            O => \N__47335\,
            I => \N__46862\
        );

    \I__11239\ : ClkMux
    port map (
            O => \N__47334\,
            I => \N__46862\
        );

    \I__11238\ : ClkMux
    port map (
            O => \N__47333\,
            I => \N__46862\
        );

    \I__11237\ : ClkMux
    port map (
            O => \N__47332\,
            I => \N__46862\
        );

    \I__11236\ : ClkMux
    port map (
            O => \N__47331\,
            I => \N__46862\
        );

    \I__11235\ : ClkMux
    port map (
            O => \N__47330\,
            I => \N__46862\
        );

    \I__11234\ : ClkMux
    port map (
            O => \N__47329\,
            I => \N__46862\
        );

    \I__11233\ : ClkMux
    port map (
            O => \N__47328\,
            I => \N__46862\
        );

    \I__11232\ : ClkMux
    port map (
            O => \N__47327\,
            I => \N__46862\
        );

    \I__11231\ : ClkMux
    port map (
            O => \N__47326\,
            I => \N__46862\
        );

    \I__11230\ : ClkMux
    port map (
            O => \N__47325\,
            I => \N__46862\
        );

    \I__11229\ : ClkMux
    port map (
            O => \N__47324\,
            I => \N__46862\
        );

    \I__11228\ : ClkMux
    port map (
            O => \N__47323\,
            I => \N__46862\
        );

    \I__11227\ : ClkMux
    port map (
            O => \N__47322\,
            I => \N__46862\
        );

    \I__11226\ : ClkMux
    port map (
            O => \N__47321\,
            I => \N__46862\
        );

    \I__11225\ : ClkMux
    port map (
            O => \N__47320\,
            I => \N__46862\
        );

    \I__11224\ : ClkMux
    port map (
            O => \N__47319\,
            I => \N__46862\
        );

    \I__11223\ : ClkMux
    port map (
            O => \N__47318\,
            I => \N__46862\
        );

    \I__11222\ : ClkMux
    port map (
            O => \N__47317\,
            I => \N__46862\
        );

    \I__11221\ : ClkMux
    port map (
            O => \N__47316\,
            I => \N__46862\
        );

    \I__11220\ : ClkMux
    port map (
            O => \N__47315\,
            I => \N__46862\
        );

    \I__11219\ : ClkMux
    port map (
            O => \N__47314\,
            I => \N__46862\
        );

    \I__11218\ : ClkMux
    port map (
            O => \N__47313\,
            I => \N__46862\
        );

    \I__11217\ : ClkMux
    port map (
            O => \N__47312\,
            I => \N__46862\
        );

    \I__11216\ : ClkMux
    port map (
            O => \N__47311\,
            I => \N__46862\
        );

    \I__11215\ : ClkMux
    port map (
            O => \N__47310\,
            I => \N__46862\
        );

    \I__11214\ : ClkMux
    port map (
            O => \N__47309\,
            I => \N__46862\
        );

    \I__11213\ : ClkMux
    port map (
            O => \N__47308\,
            I => \N__46862\
        );

    \I__11212\ : ClkMux
    port map (
            O => \N__47307\,
            I => \N__46862\
        );

    \I__11211\ : ClkMux
    port map (
            O => \N__47306\,
            I => \N__46862\
        );

    \I__11210\ : ClkMux
    port map (
            O => \N__47305\,
            I => \N__46862\
        );

    \I__11209\ : ClkMux
    port map (
            O => \N__47304\,
            I => \N__46862\
        );

    \I__11208\ : ClkMux
    port map (
            O => \N__47303\,
            I => \N__46862\
        );

    \I__11207\ : ClkMux
    port map (
            O => \N__47302\,
            I => \N__46862\
        );

    \I__11206\ : ClkMux
    port map (
            O => \N__47301\,
            I => \N__46862\
        );

    \I__11205\ : ClkMux
    port map (
            O => \N__47300\,
            I => \N__46862\
        );

    \I__11204\ : ClkMux
    port map (
            O => \N__47299\,
            I => \N__46862\
        );

    \I__11203\ : ClkMux
    port map (
            O => \N__47298\,
            I => \N__46862\
        );

    \I__11202\ : ClkMux
    port map (
            O => \N__47297\,
            I => \N__46862\
        );

    \I__11201\ : ClkMux
    port map (
            O => \N__47296\,
            I => \N__46862\
        );

    \I__11200\ : ClkMux
    port map (
            O => \N__47295\,
            I => \N__46862\
        );

    \I__11199\ : ClkMux
    port map (
            O => \N__47294\,
            I => \N__46862\
        );

    \I__11198\ : ClkMux
    port map (
            O => \N__47293\,
            I => \N__46862\
        );

    \I__11197\ : ClkMux
    port map (
            O => \N__47292\,
            I => \N__46862\
        );

    \I__11196\ : ClkMux
    port map (
            O => \N__47291\,
            I => \N__46862\
        );

    \I__11195\ : ClkMux
    port map (
            O => \N__47290\,
            I => \N__46862\
        );

    \I__11194\ : ClkMux
    port map (
            O => \N__47289\,
            I => \N__46862\
        );

    \I__11193\ : ClkMux
    port map (
            O => \N__47288\,
            I => \N__46862\
        );

    \I__11192\ : ClkMux
    port map (
            O => \N__47287\,
            I => \N__46862\
        );

    \I__11191\ : ClkMux
    port map (
            O => \N__47286\,
            I => \N__46862\
        );

    \I__11190\ : ClkMux
    port map (
            O => \N__47285\,
            I => \N__46862\
        );

    \I__11189\ : ClkMux
    port map (
            O => \N__47284\,
            I => \N__46862\
        );

    \I__11188\ : ClkMux
    port map (
            O => \N__47283\,
            I => \N__46862\
        );

    \I__11187\ : ClkMux
    port map (
            O => \N__47282\,
            I => \N__46862\
        );

    \I__11186\ : ClkMux
    port map (
            O => \N__47281\,
            I => \N__46862\
        );

    \I__11185\ : ClkMux
    port map (
            O => \N__47280\,
            I => \N__46862\
        );

    \I__11184\ : ClkMux
    port map (
            O => \N__47279\,
            I => \N__46862\
        );

    \I__11183\ : ClkMux
    port map (
            O => \N__47278\,
            I => \N__46862\
        );

    \I__11182\ : ClkMux
    port map (
            O => \N__47277\,
            I => \N__46862\
        );

    \I__11181\ : ClkMux
    port map (
            O => \N__47276\,
            I => \N__46862\
        );

    \I__11180\ : ClkMux
    port map (
            O => \N__47275\,
            I => \N__46862\
        );

    \I__11179\ : ClkMux
    port map (
            O => \N__47274\,
            I => \N__46862\
        );

    \I__11178\ : ClkMux
    port map (
            O => \N__47273\,
            I => \N__46862\
        );

    \I__11177\ : ClkMux
    port map (
            O => \N__47272\,
            I => \N__46862\
        );

    \I__11176\ : ClkMux
    port map (
            O => \N__47271\,
            I => \N__46862\
        );

    \I__11175\ : ClkMux
    port map (
            O => \N__47270\,
            I => \N__46862\
        );

    \I__11174\ : ClkMux
    port map (
            O => \N__47269\,
            I => \N__46862\
        );

    \I__11173\ : ClkMux
    port map (
            O => \N__47268\,
            I => \N__46862\
        );

    \I__11172\ : ClkMux
    port map (
            O => \N__47267\,
            I => \N__46862\
        );

    \I__11171\ : ClkMux
    port map (
            O => \N__47266\,
            I => \N__46862\
        );

    \I__11170\ : ClkMux
    port map (
            O => \N__47265\,
            I => \N__46862\
        );

    \I__11169\ : ClkMux
    port map (
            O => \N__47264\,
            I => \N__46862\
        );

    \I__11168\ : ClkMux
    port map (
            O => \N__47263\,
            I => \N__46862\
        );

    \I__11167\ : ClkMux
    port map (
            O => \N__47262\,
            I => \N__46862\
        );

    \I__11166\ : ClkMux
    port map (
            O => \N__47261\,
            I => \N__46862\
        );

    \I__11165\ : ClkMux
    port map (
            O => \N__47260\,
            I => \N__46862\
        );

    \I__11164\ : ClkMux
    port map (
            O => \N__47259\,
            I => \N__46862\
        );

    \I__11163\ : ClkMux
    port map (
            O => \N__47258\,
            I => \N__46862\
        );

    \I__11162\ : ClkMux
    port map (
            O => \N__47257\,
            I => \N__46862\
        );

    \I__11161\ : ClkMux
    port map (
            O => \N__47256\,
            I => \N__46862\
        );

    \I__11160\ : ClkMux
    port map (
            O => \N__47255\,
            I => \N__46862\
        );

    \I__11159\ : ClkMux
    port map (
            O => \N__47254\,
            I => \N__46862\
        );

    \I__11158\ : ClkMux
    port map (
            O => \N__47253\,
            I => \N__46862\
        );

    \I__11157\ : ClkMux
    port map (
            O => \N__47252\,
            I => \N__46862\
        );

    \I__11156\ : ClkMux
    port map (
            O => \N__47251\,
            I => \N__46862\
        );

    \I__11155\ : ClkMux
    port map (
            O => \N__47250\,
            I => \N__46862\
        );

    \I__11154\ : ClkMux
    port map (
            O => \N__47249\,
            I => \N__46862\
        );

    \I__11153\ : ClkMux
    port map (
            O => \N__47248\,
            I => \N__46862\
        );

    \I__11152\ : ClkMux
    port map (
            O => \N__47247\,
            I => \N__46862\
        );

    \I__11151\ : ClkMux
    port map (
            O => \N__47246\,
            I => \N__46862\
        );

    \I__11150\ : ClkMux
    port map (
            O => \N__47245\,
            I => \N__46862\
        );

    \I__11149\ : ClkMux
    port map (
            O => \N__47244\,
            I => \N__46862\
        );

    \I__11148\ : ClkMux
    port map (
            O => \N__47243\,
            I => \N__46862\
        );

    \I__11147\ : ClkMux
    port map (
            O => \N__47242\,
            I => \N__46862\
        );

    \I__11146\ : ClkMux
    port map (
            O => \N__47241\,
            I => \N__46862\
        );

    \I__11145\ : ClkMux
    port map (
            O => \N__47240\,
            I => \N__46862\
        );

    \I__11144\ : ClkMux
    port map (
            O => \N__47239\,
            I => \N__46862\
        );

    \I__11143\ : ClkMux
    port map (
            O => \N__47238\,
            I => \N__46862\
        );

    \I__11142\ : ClkMux
    port map (
            O => \N__47237\,
            I => \N__46862\
        );

    \I__11141\ : ClkMux
    port map (
            O => \N__47236\,
            I => \N__46862\
        );

    \I__11140\ : ClkMux
    port map (
            O => \N__47235\,
            I => \N__46862\
        );

    \I__11139\ : ClkMux
    port map (
            O => \N__47234\,
            I => \N__46862\
        );

    \I__11138\ : ClkMux
    port map (
            O => \N__47233\,
            I => \N__46862\
        );

    \I__11137\ : ClkMux
    port map (
            O => \N__47232\,
            I => \N__46862\
        );

    \I__11136\ : ClkMux
    port map (
            O => \N__47231\,
            I => \N__46862\
        );

    \I__11135\ : ClkMux
    port map (
            O => \N__47230\,
            I => \N__46862\
        );

    \I__11134\ : ClkMux
    port map (
            O => \N__47229\,
            I => \N__46862\
        );

    \I__11133\ : ClkMux
    port map (
            O => \N__47228\,
            I => \N__46862\
        );

    \I__11132\ : ClkMux
    port map (
            O => \N__47227\,
            I => \N__46862\
        );

    \I__11131\ : ClkMux
    port map (
            O => \N__47226\,
            I => \N__46862\
        );

    \I__11130\ : ClkMux
    port map (
            O => \N__47225\,
            I => \N__46862\
        );

    \I__11129\ : ClkMux
    port map (
            O => \N__47224\,
            I => \N__46862\
        );

    \I__11128\ : ClkMux
    port map (
            O => \N__47223\,
            I => \N__46862\
        );

    \I__11127\ : ClkMux
    port map (
            O => \N__47222\,
            I => \N__46862\
        );

    \I__11126\ : ClkMux
    port map (
            O => \N__47221\,
            I => \N__46862\
        );

    \I__11125\ : ClkMux
    port map (
            O => \N__47220\,
            I => \N__46862\
        );

    \I__11124\ : ClkMux
    port map (
            O => \N__47219\,
            I => \N__46862\
        );

    \I__11123\ : ClkMux
    port map (
            O => \N__47218\,
            I => \N__46862\
        );

    \I__11122\ : ClkMux
    port map (
            O => \N__47217\,
            I => \N__46862\
        );

    \I__11121\ : ClkMux
    port map (
            O => \N__47216\,
            I => \N__46862\
        );

    \I__11120\ : ClkMux
    port map (
            O => \N__47215\,
            I => \N__46862\
        );

    \I__11119\ : ClkMux
    port map (
            O => \N__47214\,
            I => \N__46862\
        );

    \I__11118\ : ClkMux
    port map (
            O => \N__47213\,
            I => \N__46862\
        );

    \I__11117\ : ClkMux
    port map (
            O => \N__47212\,
            I => \N__46862\
        );

    \I__11116\ : ClkMux
    port map (
            O => \N__47211\,
            I => \N__46862\
        );

    \I__11115\ : ClkMux
    port map (
            O => \N__47210\,
            I => \N__46862\
        );

    \I__11114\ : ClkMux
    port map (
            O => \N__47209\,
            I => \N__46862\
        );

    \I__11113\ : ClkMux
    port map (
            O => \N__47208\,
            I => \N__46862\
        );

    \I__11112\ : ClkMux
    port map (
            O => \N__47207\,
            I => \N__46862\
        );

    \I__11111\ : ClkMux
    port map (
            O => \N__47206\,
            I => \N__46862\
        );

    \I__11110\ : ClkMux
    port map (
            O => \N__47205\,
            I => \N__46862\
        );

    \I__11109\ : ClkMux
    port map (
            O => \N__47204\,
            I => \N__46862\
        );

    \I__11108\ : ClkMux
    port map (
            O => \N__47203\,
            I => \N__46862\
        );

    \I__11107\ : ClkMux
    port map (
            O => \N__47202\,
            I => \N__46862\
        );

    \I__11106\ : ClkMux
    port map (
            O => \N__47201\,
            I => \N__46862\
        );

    \I__11105\ : ClkMux
    port map (
            O => \N__47200\,
            I => \N__46862\
        );

    \I__11104\ : ClkMux
    port map (
            O => \N__47199\,
            I => \N__46862\
        );

    \I__11103\ : ClkMux
    port map (
            O => \N__47198\,
            I => \N__46862\
        );

    \I__11102\ : ClkMux
    port map (
            O => \N__47197\,
            I => \N__46862\
        );

    \I__11101\ : ClkMux
    port map (
            O => \N__47196\,
            I => \N__46862\
        );

    \I__11100\ : ClkMux
    port map (
            O => \N__47195\,
            I => \N__46862\
        );

    \I__11099\ : ClkMux
    port map (
            O => \N__47194\,
            I => \N__46862\
        );

    \I__11098\ : ClkMux
    port map (
            O => \N__47193\,
            I => \N__46862\
        );

    \I__11097\ : ClkMux
    port map (
            O => \N__47192\,
            I => \N__46862\
        );

    \I__11096\ : ClkMux
    port map (
            O => \N__47191\,
            I => \N__46862\
        );

    \I__11095\ : ClkMux
    port map (
            O => \N__47190\,
            I => \N__46862\
        );

    \I__11094\ : ClkMux
    port map (
            O => \N__47189\,
            I => \N__46862\
        );

    \I__11093\ : GlobalMux
    port map (
            O => \N__46862\,
            I => clk_100mhz_0
        );

    \I__11092\ : CEMux
    port map (
            O => \N__46859\,
            I => \N__46853\
        );

    \I__11091\ : CEMux
    port map (
            O => \N__46858\,
            I => \N__46849\
        );

    \I__11090\ : CEMux
    port map (
            O => \N__46857\,
            I => \N__46846\
        );

    \I__11089\ : CEMux
    port map (
            O => \N__46856\,
            I => \N__46843\
        );

    \I__11088\ : LocalMux
    port map (
            O => \N__46853\,
            I => \N__46840\
        );

    \I__11087\ : CEMux
    port map (
            O => \N__46852\,
            I => \N__46837\
        );

    \I__11086\ : LocalMux
    port map (
            O => \N__46849\,
            I => \N__46834\
        );

    \I__11085\ : LocalMux
    port map (
            O => \N__46846\,
            I => \N__46831\
        );

    \I__11084\ : LocalMux
    port map (
            O => \N__46843\,
            I => \N__46828\
        );

    \I__11083\ : Span4Mux_v
    port map (
            O => \N__46840\,
            I => \N__46823\
        );

    \I__11082\ : LocalMux
    port map (
            O => \N__46837\,
            I => \N__46820\
        );

    \I__11081\ : Span4Mux_v
    port map (
            O => \N__46834\,
            I => \N__46817\
        );

    \I__11080\ : Span4Mux_h
    port map (
            O => \N__46831\,
            I => \N__46812\
        );

    \I__11079\ : Span4Mux_h
    port map (
            O => \N__46828\,
            I => \N__46812\
        );

    \I__11078\ : CEMux
    port map (
            O => \N__46827\,
            I => \N__46809\
        );

    \I__11077\ : CEMux
    port map (
            O => \N__46826\,
            I => \N__46806\
        );

    \I__11076\ : Span4Mux_h
    port map (
            O => \N__46823\,
            I => \N__46801\
        );

    \I__11075\ : Span4Mux_v
    port map (
            O => \N__46820\,
            I => \N__46801\
        );

    \I__11074\ : Span4Mux_h
    port map (
            O => \N__46817\,
            I => \N__46796\
        );

    \I__11073\ : Span4Mux_h
    port map (
            O => \N__46812\,
            I => \N__46796\
        );

    \I__11072\ : LocalMux
    port map (
            O => \N__46809\,
            I => \N__46793\
        );

    \I__11071\ : LocalMux
    port map (
            O => \N__46806\,
            I => \N__46790\
        );

    \I__11070\ : Odrv4
    port map (
            O => \N__46801\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__11069\ : Odrv4
    port map (
            O => \N__46796\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__11068\ : Odrv4
    port map (
            O => \N__46793\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__11067\ : Odrv12
    port map (
            O => \N__46790\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__11066\ : CascadeMux
    port map (
            O => \N__46781\,
            I => \N__46774\
        );

    \I__11065\ : InMux
    port map (
            O => \N__46780\,
            I => \N__46770\
        );

    \I__11064\ : InMux
    port map (
            O => \N__46779\,
            I => \N__46767\
        );

    \I__11063\ : InMux
    port map (
            O => \N__46778\,
            I => \N__46764\
        );

    \I__11062\ : InMux
    port map (
            O => \N__46777\,
            I => \N__46761\
        );

    \I__11061\ : InMux
    port map (
            O => \N__46774\,
            I => \N__46758\
        );

    \I__11060\ : InMux
    port map (
            O => \N__46773\,
            I => \N__46755\
        );

    \I__11059\ : LocalMux
    port map (
            O => \N__46770\,
            I => \N__46752\
        );

    \I__11058\ : LocalMux
    port map (
            O => \N__46767\,
            I => \N__46749\
        );

    \I__11057\ : LocalMux
    port map (
            O => \N__46764\,
            I => \N__46746\
        );

    \I__11056\ : LocalMux
    port map (
            O => \N__46761\,
            I => \N__46698\
        );

    \I__11055\ : LocalMux
    port map (
            O => \N__46758\,
            I => \N__46624\
        );

    \I__11054\ : LocalMux
    port map (
            O => \N__46755\,
            I => \N__46621\
        );

    \I__11053\ : Glb2LocalMux
    port map (
            O => \N__46752\,
            I => \N__46298\
        );

    \I__11052\ : Glb2LocalMux
    port map (
            O => \N__46749\,
            I => \N__46298\
        );

    \I__11051\ : Glb2LocalMux
    port map (
            O => \N__46746\,
            I => \N__46298\
        );

    \I__11050\ : SRMux
    port map (
            O => \N__46745\,
            I => \N__46298\
        );

    \I__11049\ : SRMux
    port map (
            O => \N__46744\,
            I => \N__46298\
        );

    \I__11048\ : SRMux
    port map (
            O => \N__46743\,
            I => \N__46298\
        );

    \I__11047\ : SRMux
    port map (
            O => \N__46742\,
            I => \N__46298\
        );

    \I__11046\ : SRMux
    port map (
            O => \N__46741\,
            I => \N__46298\
        );

    \I__11045\ : SRMux
    port map (
            O => \N__46740\,
            I => \N__46298\
        );

    \I__11044\ : SRMux
    port map (
            O => \N__46739\,
            I => \N__46298\
        );

    \I__11043\ : SRMux
    port map (
            O => \N__46738\,
            I => \N__46298\
        );

    \I__11042\ : SRMux
    port map (
            O => \N__46737\,
            I => \N__46298\
        );

    \I__11041\ : SRMux
    port map (
            O => \N__46736\,
            I => \N__46298\
        );

    \I__11040\ : SRMux
    port map (
            O => \N__46735\,
            I => \N__46298\
        );

    \I__11039\ : SRMux
    port map (
            O => \N__46734\,
            I => \N__46298\
        );

    \I__11038\ : SRMux
    port map (
            O => \N__46733\,
            I => \N__46298\
        );

    \I__11037\ : SRMux
    port map (
            O => \N__46732\,
            I => \N__46298\
        );

    \I__11036\ : SRMux
    port map (
            O => \N__46731\,
            I => \N__46298\
        );

    \I__11035\ : SRMux
    port map (
            O => \N__46730\,
            I => \N__46298\
        );

    \I__11034\ : SRMux
    port map (
            O => \N__46729\,
            I => \N__46298\
        );

    \I__11033\ : SRMux
    port map (
            O => \N__46728\,
            I => \N__46298\
        );

    \I__11032\ : SRMux
    port map (
            O => \N__46727\,
            I => \N__46298\
        );

    \I__11031\ : SRMux
    port map (
            O => \N__46726\,
            I => \N__46298\
        );

    \I__11030\ : SRMux
    port map (
            O => \N__46725\,
            I => \N__46298\
        );

    \I__11029\ : SRMux
    port map (
            O => \N__46724\,
            I => \N__46298\
        );

    \I__11028\ : SRMux
    port map (
            O => \N__46723\,
            I => \N__46298\
        );

    \I__11027\ : SRMux
    port map (
            O => \N__46722\,
            I => \N__46298\
        );

    \I__11026\ : SRMux
    port map (
            O => \N__46721\,
            I => \N__46298\
        );

    \I__11025\ : SRMux
    port map (
            O => \N__46720\,
            I => \N__46298\
        );

    \I__11024\ : SRMux
    port map (
            O => \N__46719\,
            I => \N__46298\
        );

    \I__11023\ : SRMux
    port map (
            O => \N__46718\,
            I => \N__46298\
        );

    \I__11022\ : SRMux
    port map (
            O => \N__46717\,
            I => \N__46298\
        );

    \I__11021\ : SRMux
    port map (
            O => \N__46716\,
            I => \N__46298\
        );

    \I__11020\ : SRMux
    port map (
            O => \N__46715\,
            I => \N__46298\
        );

    \I__11019\ : SRMux
    port map (
            O => \N__46714\,
            I => \N__46298\
        );

    \I__11018\ : SRMux
    port map (
            O => \N__46713\,
            I => \N__46298\
        );

    \I__11017\ : SRMux
    port map (
            O => \N__46712\,
            I => \N__46298\
        );

    \I__11016\ : SRMux
    port map (
            O => \N__46711\,
            I => \N__46298\
        );

    \I__11015\ : SRMux
    port map (
            O => \N__46710\,
            I => \N__46298\
        );

    \I__11014\ : SRMux
    port map (
            O => \N__46709\,
            I => \N__46298\
        );

    \I__11013\ : SRMux
    port map (
            O => \N__46708\,
            I => \N__46298\
        );

    \I__11012\ : SRMux
    port map (
            O => \N__46707\,
            I => \N__46298\
        );

    \I__11011\ : SRMux
    port map (
            O => \N__46706\,
            I => \N__46298\
        );

    \I__11010\ : SRMux
    port map (
            O => \N__46705\,
            I => \N__46298\
        );

    \I__11009\ : SRMux
    port map (
            O => \N__46704\,
            I => \N__46298\
        );

    \I__11008\ : SRMux
    port map (
            O => \N__46703\,
            I => \N__46298\
        );

    \I__11007\ : SRMux
    port map (
            O => \N__46702\,
            I => \N__46298\
        );

    \I__11006\ : SRMux
    port map (
            O => \N__46701\,
            I => \N__46298\
        );

    \I__11005\ : Glb2LocalMux
    port map (
            O => \N__46698\,
            I => \N__46298\
        );

    \I__11004\ : SRMux
    port map (
            O => \N__46697\,
            I => \N__46298\
        );

    \I__11003\ : SRMux
    port map (
            O => \N__46696\,
            I => \N__46298\
        );

    \I__11002\ : SRMux
    port map (
            O => \N__46695\,
            I => \N__46298\
        );

    \I__11001\ : SRMux
    port map (
            O => \N__46694\,
            I => \N__46298\
        );

    \I__11000\ : SRMux
    port map (
            O => \N__46693\,
            I => \N__46298\
        );

    \I__10999\ : SRMux
    port map (
            O => \N__46692\,
            I => \N__46298\
        );

    \I__10998\ : SRMux
    port map (
            O => \N__46691\,
            I => \N__46298\
        );

    \I__10997\ : SRMux
    port map (
            O => \N__46690\,
            I => \N__46298\
        );

    \I__10996\ : SRMux
    port map (
            O => \N__46689\,
            I => \N__46298\
        );

    \I__10995\ : SRMux
    port map (
            O => \N__46688\,
            I => \N__46298\
        );

    \I__10994\ : SRMux
    port map (
            O => \N__46687\,
            I => \N__46298\
        );

    \I__10993\ : SRMux
    port map (
            O => \N__46686\,
            I => \N__46298\
        );

    \I__10992\ : SRMux
    port map (
            O => \N__46685\,
            I => \N__46298\
        );

    \I__10991\ : SRMux
    port map (
            O => \N__46684\,
            I => \N__46298\
        );

    \I__10990\ : SRMux
    port map (
            O => \N__46683\,
            I => \N__46298\
        );

    \I__10989\ : SRMux
    port map (
            O => \N__46682\,
            I => \N__46298\
        );

    \I__10988\ : SRMux
    port map (
            O => \N__46681\,
            I => \N__46298\
        );

    \I__10987\ : SRMux
    port map (
            O => \N__46680\,
            I => \N__46298\
        );

    \I__10986\ : SRMux
    port map (
            O => \N__46679\,
            I => \N__46298\
        );

    \I__10985\ : SRMux
    port map (
            O => \N__46678\,
            I => \N__46298\
        );

    \I__10984\ : SRMux
    port map (
            O => \N__46677\,
            I => \N__46298\
        );

    \I__10983\ : SRMux
    port map (
            O => \N__46676\,
            I => \N__46298\
        );

    \I__10982\ : SRMux
    port map (
            O => \N__46675\,
            I => \N__46298\
        );

    \I__10981\ : SRMux
    port map (
            O => \N__46674\,
            I => \N__46298\
        );

    \I__10980\ : SRMux
    port map (
            O => \N__46673\,
            I => \N__46298\
        );

    \I__10979\ : SRMux
    port map (
            O => \N__46672\,
            I => \N__46298\
        );

    \I__10978\ : SRMux
    port map (
            O => \N__46671\,
            I => \N__46298\
        );

    \I__10977\ : SRMux
    port map (
            O => \N__46670\,
            I => \N__46298\
        );

    \I__10976\ : SRMux
    port map (
            O => \N__46669\,
            I => \N__46298\
        );

    \I__10975\ : SRMux
    port map (
            O => \N__46668\,
            I => \N__46298\
        );

    \I__10974\ : SRMux
    port map (
            O => \N__46667\,
            I => \N__46298\
        );

    \I__10973\ : SRMux
    port map (
            O => \N__46666\,
            I => \N__46298\
        );

    \I__10972\ : SRMux
    port map (
            O => \N__46665\,
            I => \N__46298\
        );

    \I__10971\ : SRMux
    port map (
            O => \N__46664\,
            I => \N__46298\
        );

    \I__10970\ : SRMux
    port map (
            O => \N__46663\,
            I => \N__46298\
        );

    \I__10969\ : SRMux
    port map (
            O => \N__46662\,
            I => \N__46298\
        );

    \I__10968\ : SRMux
    port map (
            O => \N__46661\,
            I => \N__46298\
        );

    \I__10967\ : SRMux
    port map (
            O => \N__46660\,
            I => \N__46298\
        );

    \I__10966\ : SRMux
    port map (
            O => \N__46659\,
            I => \N__46298\
        );

    \I__10965\ : SRMux
    port map (
            O => \N__46658\,
            I => \N__46298\
        );

    \I__10964\ : SRMux
    port map (
            O => \N__46657\,
            I => \N__46298\
        );

    \I__10963\ : SRMux
    port map (
            O => \N__46656\,
            I => \N__46298\
        );

    \I__10962\ : SRMux
    port map (
            O => \N__46655\,
            I => \N__46298\
        );

    \I__10961\ : SRMux
    port map (
            O => \N__46654\,
            I => \N__46298\
        );

    \I__10960\ : SRMux
    port map (
            O => \N__46653\,
            I => \N__46298\
        );

    \I__10959\ : SRMux
    port map (
            O => \N__46652\,
            I => \N__46298\
        );

    \I__10958\ : SRMux
    port map (
            O => \N__46651\,
            I => \N__46298\
        );

    \I__10957\ : SRMux
    port map (
            O => \N__46650\,
            I => \N__46298\
        );

    \I__10956\ : SRMux
    port map (
            O => \N__46649\,
            I => \N__46298\
        );

    \I__10955\ : SRMux
    port map (
            O => \N__46648\,
            I => \N__46298\
        );

    \I__10954\ : SRMux
    port map (
            O => \N__46647\,
            I => \N__46298\
        );

    \I__10953\ : SRMux
    port map (
            O => \N__46646\,
            I => \N__46298\
        );

    \I__10952\ : SRMux
    port map (
            O => \N__46645\,
            I => \N__46298\
        );

    \I__10951\ : SRMux
    port map (
            O => \N__46644\,
            I => \N__46298\
        );

    \I__10950\ : SRMux
    port map (
            O => \N__46643\,
            I => \N__46298\
        );

    \I__10949\ : SRMux
    port map (
            O => \N__46642\,
            I => \N__46298\
        );

    \I__10948\ : SRMux
    port map (
            O => \N__46641\,
            I => \N__46298\
        );

    \I__10947\ : SRMux
    port map (
            O => \N__46640\,
            I => \N__46298\
        );

    \I__10946\ : SRMux
    port map (
            O => \N__46639\,
            I => \N__46298\
        );

    \I__10945\ : SRMux
    port map (
            O => \N__46638\,
            I => \N__46298\
        );

    \I__10944\ : SRMux
    port map (
            O => \N__46637\,
            I => \N__46298\
        );

    \I__10943\ : SRMux
    port map (
            O => \N__46636\,
            I => \N__46298\
        );

    \I__10942\ : SRMux
    port map (
            O => \N__46635\,
            I => \N__46298\
        );

    \I__10941\ : SRMux
    port map (
            O => \N__46634\,
            I => \N__46298\
        );

    \I__10940\ : SRMux
    port map (
            O => \N__46633\,
            I => \N__46298\
        );

    \I__10939\ : SRMux
    port map (
            O => \N__46632\,
            I => \N__46298\
        );

    \I__10938\ : SRMux
    port map (
            O => \N__46631\,
            I => \N__46298\
        );

    \I__10937\ : SRMux
    port map (
            O => \N__46630\,
            I => \N__46298\
        );

    \I__10936\ : SRMux
    port map (
            O => \N__46629\,
            I => \N__46298\
        );

    \I__10935\ : SRMux
    port map (
            O => \N__46628\,
            I => \N__46298\
        );

    \I__10934\ : SRMux
    port map (
            O => \N__46627\,
            I => \N__46298\
        );

    \I__10933\ : Glb2LocalMux
    port map (
            O => \N__46624\,
            I => \N__46298\
        );

    \I__10932\ : Glb2LocalMux
    port map (
            O => \N__46621\,
            I => \N__46298\
        );

    \I__10931\ : SRMux
    port map (
            O => \N__46620\,
            I => \N__46298\
        );

    \I__10930\ : SRMux
    port map (
            O => \N__46619\,
            I => \N__46298\
        );

    \I__10929\ : SRMux
    port map (
            O => \N__46618\,
            I => \N__46298\
        );

    \I__10928\ : SRMux
    port map (
            O => \N__46617\,
            I => \N__46298\
        );

    \I__10927\ : SRMux
    port map (
            O => \N__46616\,
            I => \N__46298\
        );

    \I__10926\ : SRMux
    port map (
            O => \N__46615\,
            I => \N__46298\
        );

    \I__10925\ : SRMux
    port map (
            O => \N__46614\,
            I => \N__46298\
        );

    \I__10924\ : SRMux
    port map (
            O => \N__46613\,
            I => \N__46298\
        );

    \I__10923\ : SRMux
    port map (
            O => \N__46612\,
            I => \N__46298\
        );

    \I__10922\ : SRMux
    port map (
            O => \N__46611\,
            I => \N__46298\
        );

    \I__10921\ : SRMux
    port map (
            O => \N__46610\,
            I => \N__46298\
        );

    \I__10920\ : SRMux
    port map (
            O => \N__46609\,
            I => \N__46298\
        );

    \I__10919\ : SRMux
    port map (
            O => \N__46608\,
            I => \N__46298\
        );

    \I__10918\ : SRMux
    port map (
            O => \N__46607\,
            I => \N__46298\
        );

    \I__10917\ : SRMux
    port map (
            O => \N__46606\,
            I => \N__46298\
        );

    \I__10916\ : SRMux
    port map (
            O => \N__46605\,
            I => \N__46298\
        );

    \I__10915\ : SRMux
    port map (
            O => \N__46604\,
            I => \N__46298\
        );

    \I__10914\ : SRMux
    port map (
            O => \N__46603\,
            I => \N__46298\
        );

    \I__10913\ : SRMux
    port map (
            O => \N__46602\,
            I => \N__46298\
        );

    \I__10912\ : SRMux
    port map (
            O => \N__46601\,
            I => \N__46298\
        );

    \I__10911\ : SRMux
    port map (
            O => \N__46600\,
            I => \N__46298\
        );

    \I__10910\ : SRMux
    port map (
            O => \N__46599\,
            I => \N__46298\
        );

    \I__10909\ : SRMux
    port map (
            O => \N__46598\,
            I => \N__46298\
        );

    \I__10908\ : SRMux
    port map (
            O => \N__46597\,
            I => \N__46298\
        );

    \I__10907\ : SRMux
    port map (
            O => \N__46596\,
            I => \N__46298\
        );

    \I__10906\ : SRMux
    port map (
            O => \N__46595\,
            I => \N__46298\
        );

    \I__10905\ : GlobalMux
    port map (
            O => \N__46298\,
            I => \N__46295\
        );

    \I__10904\ : gio2CtrlBuf
    port map (
            O => \N__46295\,
            I => red_c_g
        );

    \I__10903\ : InMux
    port map (
            O => \N__46292\,
            I => \N__46288\
        );

    \I__10902\ : InMux
    port map (
            O => \N__46291\,
            I => \N__46285\
        );

    \I__10901\ : LocalMux
    port map (
            O => \N__46288\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__10900\ : LocalMux
    port map (
            O => \N__46285\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__10899\ : InMux
    port map (
            O => \N__46280\,
            I => \N__46277\
        );

    \I__10898\ : LocalMux
    port map (
            O => \N__46277\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12\
        );

    \I__10897\ : InMux
    port map (
            O => \N__46274\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\
        );

    \I__10896\ : InMux
    port map (
            O => \N__46271\,
            I => \N__46267\
        );

    \I__10895\ : InMux
    port map (
            O => \N__46270\,
            I => \N__46264\
        );

    \I__10894\ : LocalMux
    port map (
            O => \N__46267\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__10893\ : LocalMux
    port map (
            O => \N__46264\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__10892\ : InMux
    port map (
            O => \N__46259\,
            I => \N__46256\
        );

    \I__10891\ : LocalMux
    port map (
            O => \N__46256\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13\
        );

    \I__10890\ : InMux
    port map (
            O => \N__46253\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\
        );

    \I__10889\ : InMux
    port map (
            O => \N__46250\,
            I => \N__46246\
        );

    \I__10888\ : InMux
    port map (
            O => \N__46249\,
            I => \N__46243\
        );

    \I__10887\ : LocalMux
    port map (
            O => \N__46246\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__10886\ : LocalMux
    port map (
            O => \N__46243\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__10885\ : InMux
    port map (
            O => \N__46238\,
            I => \N__46235\
        );

    \I__10884\ : LocalMux
    port map (
            O => \N__46235\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14\
        );

    \I__10883\ : InMux
    port map (
            O => \N__46232\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\
        );

    \I__10882\ : InMux
    port map (
            O => \N__46229\,
            I => \N__46226\
        );

    \I__10881\ : LocalMux
    port map (
            O => \N__46226\,
            I => \N__46222\
        );

    \I__10880\ : InMux
    port map (
            O => \N__46225\,
            I => \N__46219\
        );

    \I__10879\ : Odrv4
    port map (
            O => \N__46222\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__10878\ : LocalMux
    port map (
            O => \N__46219\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__10877\ : InMux
    port map (
            O => \N__46214\,
            I => \N__46211\
        );

    \I__10876\ : LocalMux
    port map (
            O => \N__46211\,
            I => \N__46208\
        );

    \I__10875\ : Odrv4
    port map (
            O => \N__46208\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15\
        );

    \I__10874\ : InMux
    port map (
            O => \N__46205\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\
        );

    \I__10873\ : InMux
    port map (
            O => \N__46202\,
            I => \N__46198\
        );

    \I__10872\ : InMux
    port map (
            O => \N__46201\,
            I => \N__46195\
        );

    \I__10871\ : LocalMux
    port map (
            O => \N__46198\,
            I => \N__46192\
        );

    \I__10870\ : LocalMux
    port map (
            O => \N__46195\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__10869\ : Odrv4
    port map (
            O => \N__46192\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__10868\ : InMux
    port map (
            O => \N__46187\,
            I => \N__46184\
        );

    \I__10867\ : LocalMux
    port map (
            O => \N__46184\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16\
        );

    \I__10866\ : InMux
    port map (
            O => \N__46181\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\
        );

    \I__10865\ : InMux
    port map (
            O => \N__46178\,
            I => \N__46174\
        );

    \I__10864\ : InMux
    port map (
            O => \N__46177\,
            I => \N__46171\
        );

    \I__10863\ : LocalMux
    port map (
            O => \N__46174\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__10862\ : LocalMux
    port map (
            O => \N__46171\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__10861\ : InMux
    port map (
            O => \N__46166\,
            I => \N__46163\
        );

    \I__10860\ : LocalMux
    port map (
            O => \N__46163\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17\
        );

    \I__10859\ : InMux
    port map (
            O => \N__46160\,
            I => \bfn_18_19_0_\
        );

    \I__10858\ : InMux
    port map (
            O => \N__46157\,
            I => \N__46153\
        );

    \I__10857\ : InMux
    port map (
            O => \N__46156\,
            I => \N__46150\
        );

    \I__10856\ : LocalMux
    port map (
            O => \N__46153\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__10855\ : LocalMux
    port map (
            O => \N__46150\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__10854\ : InMux
    port map (
            O => \N__46145\,
            I => \N__46142\
        );

    \I__10853\ : LocalMux
    port map (
            O => \N__46142\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18\
        );

    \I__10852\ : InMux
    port map (
            O => \N__46139\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\
        );

    \I__10851\ : InMux
    port map (
            O => \N__46136\,
            I => \N__46132\
        );

    \I__10850\ : InMux
    port map (
            O => \N__46135\,
            I => \N__46129\
        );

    \I__10849\ : LocalMux
    port map (
            O => \N__46132\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__10848\ : LocalMux
    port map (
            O => \N__46129\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__10847\ : InMux
    port map (
            O => \N__46124\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17\
        );

    \I__10846\ : InMux
    port map (
            O => \N__46121\,
            I => \N__46118\
        );

    \I__10845\ : LocalMux
    port map (
            O => \N__46118\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19\
        );

    \I__10844\ : CascadeMux
    port map (
            O => \N__46115\,
            I => \N__46112\
        );

    \I__10843\ : InMux
    port map (
            O => \N__46112\,
            I => \N__46108\
        );

    \I__10842\ : InMux
    port map (
            O => \N__46111\,
            I => \N__46105\
        );

    \I__10841\ : LocalMux
    port map (
            O => \N__46108\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__10840\ : LocalMux
    port map (
            O => \N__46105\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__10839\ : InMux
    port map (
            O => \N__46100\,
            I => \N__46097\
        );

    \I__10838\ : LocalMux
    port map (
            O => \N__46097\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4\
        );

    \I__10837\ : InMux
    port map (
            O => \N__46094\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\
        );

    \I__10836\ : InMux
    port map (
            O => \N__46091\,
            I => \N__46087\
        );

    \I__10835\ : InMux
    port map (
            O => \N__46090\,
            I => \N__46084\
        );

    \I__10834\ : LocalMux
    port map (
            O => \N__46087\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__10833\ : LocalMux
    port map (
            O => \N__46084\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__10832\ : InMux
    port map (
            O => \N__46079\,
            I => \N__46076\
        );

    \I__10831\ : LocalMux
    port map (
            O => \N__46076\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5\
        );

    \I__10830\ : InMux
    port map (
            O => \N__46073\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\
        );

    \I__10829\ : InMux
    port map (
            O => \N__46070\,
            I => \N__46066\
        );

    \I__10828\ : InMux
    port map (
            O => \N__46069\,
            I => \N__46063\
        );

    \I__10827\ : LocalMux
    port map (
            O => \N__46066\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__10826\ : LocalMux
    port map (
            O => \N__46063\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__10825\ : InMux
    port map (
            O => \N__46058\,
            I => \N__46055\
        );

    \I__10824\ : LocalMux
    port map (
            O => \N__46055\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6\
        );

    \I__10823\ : InMux
    port map (
            O => \N__46052\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\
        );

    \I__10822\ : InMux
    port map (
            O => \N__46049\,
            I => \N__46045\
        );

    \I__10821\ : InMux
    port map (
            O => \N__46048\,
            I => \N__46042\
        );

    \I__10820\ : LocalMux
    port map (
            O => \N__46045\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__10819\ : LocalMux
    port map (
            O => \N__46042\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__10818\ : InMux
    port map (
            O => \N__46037\,
            I => \N__46034\
        );

    \I__10817\ : LocalMux
    port map (
            O => \N__46034\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7\
        );

    \I__10816\ : InMux
    port map (
            O => \N__46031\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\
        );

    \I__10815\ : InMux
    port map (
            O => \N__46028\,
            I => \N__46024\
        );

    \I__10814\ : InMux
    port map (
            O => \N__46027\,
            I => \N__46021\
        );

    \I__10813\ : LocalMux
    port map (
            O => \N__46024\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__10812\ : LocalMux
    port map (
            O => \N__46021\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__10811\ : InMux
    port map (
            O => \N__46016\,
            I => \N__46013\
        );

    \I__10810\ : LocalMux
    port map (
            O => \N__46013\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8\
        );

    \I__10809\ : InMux
    port map (
            O => \N__46010\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\
        );

    \I__10808\ : InMux
    port map (
            O => \N__46007\,
            I => \bfn_18_18_0_\
        );

    \I__10807\ : InMux
    port map (
            O => \N__46004\,
            I => \N__46000\
        );

    \I__10806\ : InMux
    port map (
            O => \N__46003\,
            I => \N__45997\
        );

    \I__10805\ : LocalMux
    port map (
            O => \N__46000\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__10804\ : LocalMux
    port map (
            O => \N__45997\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__10803\ : InMux
    port map (
            O => \N__45992\,
            I => \N__45989\
        );

    \I__10802\ : LocalMux
    port map (
            O => \N__45989\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10\
        );

    \I__10801\ : InMux
    port map (
            O => \N__45986\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\
        );

    \I__10800\ : InMux
    port map (
            O => \N__45983\,
            I => \N__45979\
        );

    \I__10799\ : InMux
    port map (
            O => \N__45982\,
            I => \N__45976\
        );

    \I__10798\ : LocalMux
    port map (
            O => \N__45979\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__10797\ : LocalMux
    port map (
            O => \N__45976\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__10796\ : InMux
    port map (
            O => \N__45971\,
            I => \N__45968\
        );

    \I__10795\ : LocalMux
    port map (
            O => \N__45968\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11\
        );

    \I__10794\ : InMux
    port map (
            O => \N__45965\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\
        );

    \I__10793\ : InMux
    port map (
            O => \N__45962\,
            I => \N__45959\
        );

    \I__10792\ : LocalMux
    port map (
            O => \N__45959\,
            I => \N__45955\
        );

    \I__10791\ : CascadeMux
    port map (
            O => \N__45958\,
            I => \N__45951\
        );

    \I__10790\ : Span4Mux_h
    port map (
            O => \N__45955\,
            I => \N__45948\
        );

    \I__10789\ : InMux
    port map (
            O => \N__45954\,
            I => \N__45945\
        );

    \I__10788\ : InMux
    port map (
            O => \N__45951\,
            I => \N__45942\
        );

    \I__10787\ : Odrv4
    port map (
            O => \N__45948\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__10786\ : LocalMux
    port map (
            O => \N__45945\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__10785\ : LocalMux
    port map (
            O => \N__45942\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__10784\ : CascadeMux
    port map (
            O => \N__45935\,
            I => \N__45932\
        );

    \I__10783\ : InMux
    port map (
            O => \N__45932\,
            I => \N__45929\
        );

    \I__10782\ : LocalMux
    port map (
            O => \N__45929\,
            I => \N__45926\
        );

    \I__10781\ : Span4Mux_h
    port map (
            O => \N__45926\,
            I => \N__45923\
        );

    \I__10780\ : Odrv4
    port map (
            O => \N__45923\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__10779\ : InMux
    port map (
            O => \N__45920\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__10778\ : InMux
    port map (
            O => \N__45917\,
            I => \N__45914\
        );

    \I__10777\ : LocalMux
    port map (
            O => \N__45914\,
            I => \N__45910\
        );

    \I__10776\ : InMux
    port map (
            O => \N__45913\,
            I => \N__45907\
        );

    \I__10775\ : Span4Mux_h
    port map (
            O => \N__45910\,
            I => \N__45904\
        );

    \I__10774\ : LocalMux
    port map (
            O => \N__45907\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__10773\ : Odrv4
    port map (
            O => \N__45904\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__10772\ : CascadeMux
    port map (
            O => \N__45899\,
            I => \N__45895\
        );

    \I__10771\ : CascadeMux
    port map (
            O => \N__45898\,
            I => \N__45892\
        );

    \I__10770\ : InMux
    port map (
            O => \N__45895\,
            I => \N__45886\
        );

    \I__10769\ : InMux
    port map (
            O => \N__45892\,
            I => \N__45886\
        );

    \I__10768\ : InMux
    port map (
            O => \N__45891\,
            I => \N__45883\
        );

    \I__10767\ : LocalMux
    port map (
            O => \N__45886\,
            I => \N__45880\
        );

    \I__10766\ : LocalMux
    port map (
            O => \N__45883\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__10765\ : Odrv4
    port map (
            O => \N__45880\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__10764\ : InMux
    port map (
            O => \N__45875\,
            I => \N__45872\
        );

    \I__10763\ : LocalMux
    port map (
            O => \N__45872\,
            I => \N__45869\
        );

    \I__10762\ : Span4Mux_v
    port map (
            O => \N__45869\,
            I => \N__45866\
        );

    \I__10761\ : Odrv4
    port map (
            O => \N__45866\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__10760\ : InMux
    port map (
            O => \N__45863\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__10759\ : InMux
    port map (
            O => \N__45860\,
            I => \N__45856\
        );

    \I__10758\ : InMux
    port map (
            O => \N__45859\,
            I => \N__45853\
        );

    \I__10757\ : LocalMux
    port map (
            O => \N__45856\,
            I => \N__45850\
        );

    \I__10756\ : LocalMux
    port map (
            O => \N__45853\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__10755\ : Odrv4
    port map (
            O => \N__45850\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__10754\ : CascadeMux
    port map (
            O => \N__45845\,
            I => \N__45841\
        );

    \I__10753\ : CascadeMux
    port map (
            O => \N__45844\,
            I => \N__45838\
        );

    \I__10752\ : InMux
    port map (
            O => \N__45841\,
            I => \N__45832\
        );

    \I__10751\ : InMux
    port map (
            O => \N__45838\,
            I => \N__45832\
        );

    \I__10750\ : InMux
    port map (
            O => \N__45837\,
            I => \N__45829\
        );

    \I__10749\ : LocalMux
    port map (
            O => \N__45832\,
            I => \N__45826\
        );

    \I__10748\ : LocalMux
    port map (
            O => \N__45829\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__10747\ : Odrv4
    port map (
            O => \N__45826\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__10746\ : InMux
    port map (
            O => \N__45821\,
            I => \N__45818\
        );

    \I__10745\ : LocalMux
    port map (
            O => \N__45818\,
            I => \N__45815\
        );

    \I__10744\ : Span4Mux_v
    port map (
            O => \N__45815\,
            I => \N__45812\
        );

    \I__10743\ : Odrv4
    port map (
            O => \N__45812\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30\
        );

    \I__10742\ : InMux
    port map (
            O => \N__45809\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__10741\ : InMux
    port map (
            O => \N__45806\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__10740\ : CascadeMux
    port map (
            O => \N__45803\,
            I => \N__45798\
        );

    \I__10739\ : InMux
    port map (
            O => \N__45802\,
            I => \N__45791\
        );

    \I__10738\ : CascadeMux
    port map (
            O => \N__45801\,
            I => \N__45787\
        );

    \I__10737\ : InMux
    port map (
            O => \N__45798\,
            I => \N__45782\
        );

    \I__10736\ : InMux
    port map (
            O => \N__45797\,
            I => \N__45773\
        );

    \I__10735\ : InMux
    port map (
            O => \N__45796\,
            I => \N__45773\
        );

    \I__10734\ : InMux
    port map (
            O => \N__45795\,
            I => \N__45773\
        );

    \I__10733\ : InMux
    port map (
            O => \N__45794\,
            I => \N__45773\
        );

    \I__10732\ : LocalMux
    port map (
            O => \N__45791\,
            I => \N__45770\
        );

    \I__10731\ : InMux
    port map (
            O => \N__45790\,
            I => \N__45765\
        );

    \I__10730\ : InMux
    port map (
            O => \N__45787\,
            I => \N__45765\
        );

    \I__10729\ : CascadeMux
    port map (
            O => \N__45786\,
            I => \N__45762\
        );

    \I__10728\ : InMux
    port map (
            O => \N__45785\,
            I => \N__45757\
        );

    \I__10727\ : LocalMux
    port map (
            O => \N__45782\,
            I => \N__45748\
        );

    \I__10726\ : LocalMux
    port map (
            O => \N__45773\,
            I => \N__45748\
        );

    \I__10725\ : Span4Mux_h
    port map (
            O => \N__45770\,
            I => \N__45748\
        );

    \I__10724\ : LocalMux
    port map (
            O => \N__45765\,
            I => \N__45748\
        );

    \I__10723\ : InMux
    port map (
            O => \N__45762\,
            I => \N__45741\
        );

    \I__10722\ : InMux
    port map (
            O => \N__45761\,
            I => \N__45741\
        );

    \I__10721\ : InMux
    port map (
            O => \N__45760\,
            I => \N__45741\
        );

    \I__10720\ : LocalMux
    port map (
            O => \N__45757\,
            I => \N__45736\
        );

    \I__10719\ : Span4Mux_v
    port map (
            O => \N__45748\,
            I => \N__45736\
        );

    \I__10718\ : LocalMux
    port map (
            O => \N__45741\,
            I => \delay_measurement_inst.elapsed_time_tr_31\
        );

    \I__10717\ : Odrv4
    port map (
            O => \N__45736\,
            I => \delay_measurement_inst.elapsed_time_tr_31\
        );

    \I__10716\ : CEMux
    port map (
            O => \N__45731\,
            I => \N__45728\
        );

    \I__10715\ : LocalMux
    port map (
            O => \N__45728\,
            I => \N__45722\
        );

    \I__10714\ : CEMux
    port map (
            O => \N__45727\,
            I => \N__45719\
        );

    \I__10713\ : CEMux
    port map (
            O => \N__45726\,
            I => \N__45715\
        );

    \I__10712\ : CEMux
    port map (
            O => \N__45725\,
            I => \N__45712\
        );

    \I__10711\ : Span4Mux_v
    port map (
            O => \N__45722\,
            I => \N__45707\
        );

    \I__10710\ : LocalMux
    port map (
            O => \N__45719\,
            I => \N__45707\
        );

    \I__10709\ : CEMux
    port map (
            O => \N__45718\,
            I => \N__45704\
        );

    \I__10708\ : LocalMux
    port map (
            O => \N__45715\,
            I => \N__45698\
        );

    \I__10707\ : LocalMux
    port map (
            O => \N__45712\,
            I => \N__45698\
        );

    \I__10706\ : Span4Mux_v
    port map (
            O => \N__45707\,
            I => \N__45693\
        );

    \I__10705\ : LocalMux
    port map (
            O => \N__45704\,
            I => \N__45693\
        );

    \I__10704\ : CEMux
    port map (
            O => \N__45703\,
            I => \N__45690\
        );

    \I__10703\ : Span4Mux_v
    port map (
            O => \N__45698\,
            I => \N__45687\
        );

    \I__10702\ : Span4Mux_h
    port map (
            O => \N__45693\,
            I => \N__45684\
        );

    \I__10701\ : LocalMux
    port map (
            O => \N__45690\,
            I => \N__45681\
        );

    \I__10700\ : Odrv4
    port map (
            O => \N__45687\,
            I => \delay_measurement_inst.delay_tr_timer.N_323_i\
        );

    \I__10699\ : Odrv4
    port map (
            O => \N__45684\,
            I => \delay_measurement_inst.delay_tr_timer.N_323_i\
        );

    \I__10698\ : Odrv12
    port map (
            O => \N__45681\,
            I => \delay_measurement_inst.delay_tr_timer.N_323_i\
        );

    \I__10697\ : InMux
    port map (
            O => \N__45674\,
            I => \N__45671\
        );

    \I__10696\ : LocalMux
    port map (
            O => \N__45671\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0\
        );

    \I__10695\ : CascadeMux
    port map (
            O => \N__45668\,
            I => \N__45665\
        );

    \I__10694\ : InMux
    port map (
            O => \N__45665\,
            I => \N__45661\
        );

    \I__10693\ : InMux
    port map (
            O => \N__45664\,
            I => \N__45657\
        );

    \I__10692\ : LocalMux
    port map (
            O => \N__45661\,
            I => \N__45654\
        );

    \I__10691\ : InMux
    port map (
            O => \N__45660\,
            I => \N__45651\
        );

    \I__10690\ : LocalMux
    port map (
            O => \N__45657\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__10689\ : Odrv4
    port map (
            O => \N__45654\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__10688\ : LocalMux
    port map (
            O => \N__45651\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__10687\ : InMux
    port map (
            O => \N__45644\,
            I => \N__45640\
        );

    \I__10686\ : InMux
    port map (
            O => \N__45643\,
            I => \N__45637\
        );

    \I__10685\ : LocalMux
    port map (
            O => \N__45640\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__10684\ : LocalMux
    port map (
            O => \N__45637\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__10683\ : InMux
    port map (
            O => \N__45632\,
            I => \N__45629\
        );

    \I__10682\ : LocalMux
    port map (
            O => \N__45629\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2\
        );

    \I__10681\ : InMux
    port map (
            O => \N__45626\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\
        );

    \I__10680\ : InMux
    port map (
            O => \N__45623\,
            I => \N__45620\
        );

    \I__10679\ : LocalMux
    port map (
            O => \N__45620\,
            I => \N__45617\
        );

    \I__10678\ : Odrv4
    port map (
            O => \N__45617\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0\
        );

    \I__10677\ : CascadeMux
    port map (
            O => \N__45614\,
            I => \N__45611\
        );

    \I__10676\ : InMux
    port map (
            O => \N__45611\,
            I => \N__45607\
        );

    \I__10675\ : InMux
    port map (
            O => \N__45610\,
            I => \N__45604\
        );

    \I__10674\ : LocalMux
    port map (
            O => \N__45607\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__10673\ : LocalMux
    port map (
            O => \N__45604\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__10672\ : InMux
    port map (
            O => \N__45599\,
            I => \N__45596\
        );

    \I__10671\ : LocalMux
    port map (
            O => \N__45596\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3\
        );

    \I__10670\ : InMux
    port map (
            O => \N__45593\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\
        );

    \I__10669\ : CascadeMux
    port map (
            O => \N__45590\,
            I => \N__45587\
        );

    \I__10668\ : InMux
    port map (
            O => \N__45587\,
            I => \N__45584\
        );

    \I__10667\ : LocalMux
    port map (
            O => \N__45584\,
            I => \N__45580\
        );

    \I__10666\ : InMux
    port map (
            O => \N__45583\,
            I => \N__45576\
        );

    \I__10665\ : Span4Mux_h
    port map (
            O => \N__45580\,
            I => \N__45573\
        );

    \I__10664\ : InMux
    port map (
            O => \N__45579\,
            I => \N__45570\
        );

    \I__10663\ : LocalMux
    port map (
            O => \N__45576\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__10662\ : Odrv4
    port map (
            O => \N__45573\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__10661\ : LocalMux
    port map (
            O => \N__45570\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__10660\ : InMux
    port map (
            O => \N__45563\,
            I => \N__45560\
        );

    \I__10659\ : LocalMux
    port map (
            O => \N__45560\,
            I => \N__45557\
        );

    \I__10658\ : Span4Mux_v
    port map (
            O => \N__45557\,
            I => \N__45554\
        );

    \I__10657\ : Odrv4
    port map (
            O => \N__45554\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__10656\ : InMux
    port map (
            O => \N__45551\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__10655\ : CascadeMux
    port map (
            O => \N__45548\,
            I => \N__45544\
        );

    \I__10654\ : InMux
    port map (
            O => \N__45547\,
            I => \N__45541\
        );

    \I__10653\ : InMux
    port map (
            O => \N__45544\,
            I => \N__45538\
        );

    \I__10652\ : LocalMux
    port map (
            O => \N__45541\,
            I => \N__45534\
        );

    \I__10651\ : LocalMux
    port map (
            O => \N__45538\,
            I => \N__45531\
        );

    \I__10650\ : InMux
    port map (
            O => \N__45537\,
            I => \N__45528\
        );

    \I__10649\ : Span4Mux_v
    port map (
            O => \N__45534\,
            I => \N__45525\
        );

    \I__10648\ : Span4Mux_v
    port map (
            O => \N__45531\,
            I => \N__45522\
        );

    \I__10647\ : LocalMux
    port map (
            O => \N__45528\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__10646\ : Odrv4
    port map (
            O => \N__45525\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__10645\ : Odrv4
    port map (
            O => \N__45522\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__10644\ : InMux
    port map (
            O => \N__45515\,
            I => \N__45512\
        );

    \I__10643\ : LocalMux
    port map (
            O => \N__45512\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__10642\ : InMux
    port map (
            O => \N__45509\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__10641\ : InMux
    port map (
            O => \N__45506\,
            I => \N__45499\
        );

    \I__10640\ : InMux
    port map (
            O => \N__45505\,
            I => \N__45499\
        );

    \I__10639\ : InMux
    port map (
            O => \N__45504\,
            I => \N__45496\
        );

    \I__10638\ : LocalMux
    port map (
            O => \N__45499\,
            I => \N__45493\
        );

    \I__10637\ : LocalMux
    port map (
            O => \N__45496\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__10636\ : Odrv4
    port map (
            O => \N__45493\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__10635\ : InMux
    port map (
            O => \N__45488\,
            I => \N__45485\
        );

    \I__10634\ : LocalMux
    port map (
            O => \N__45485\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__10633\ : InMux
    port map (
            O => \N__45482\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__10632\ : CascadeMux
    port map (
            O => \N__45479\,
            I => \N__45475\
        );

    \I__10631\ : CascadeMux
    port map (
            O => \N__45478\,
            I => \N__45472\
        );

    \I__10630\ : InMux
    port map (
            O => \N__45475\,
            I => \N__45466\
        );

    \I__10629\ : InMux
    port map (
            O => \N__45472\,
            I => \N__45466\
        );

    \I__10628\ : InMux
    port map (
            O => \N__45471\,
            I => \N__45463\
        );

    \I__10627\ : LocalMux
    port map (
            O => \N__45466\,
            I => \N__45460\
        );

    \I__10626\ : LocalMux
    port map (
            O => \N__45463\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__10625\ : Odrv4
    port map (
            O => \N__45460\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__10624\ : InMux
    port map (
            O => \N__45455\,
            I => \N__45452\
        );

    \I__10623\ : LocalMux
    port map (
            O => \N__45452\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__10622\ : InMux
    port map (
            O => \N__45449\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__10621\ : CascadeMux
    port map (
            O => \N__45446\,
            I => \N__45442\
        );

    \I__10620\ : CascadeMux
    port map (
            O => \N__45445\,
            I => \N__45439\
        );

    \I__10619\ : InMux
    port map (
            O => \N__45442\,
            I => \N__45433\
        );

    \I__10618\ : InMux
    port map (
            O => \N__45439\,
            I => \N__45433\
        );

    \I__10617\ : InMux
    port map (
            O => \N__45438\,
            I => \N__45430\
        );

    \I__10616\ : LocalMux
    port map (
            O => \N__45433\,
            I => \N__45427\
        );

    \I__10615\ : LocalMux
    port map (
            O => \N__45430\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__10614\ : Odrv4
    port map (
            O => \N__45427\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__10613\ : CascadeMux
    port map (
            O => \N__45422\,
            I => \N__45419\
        );

    \I__10612\ : InMux
    port map (
            O => \N__45419\,
            I => \N__45416\
        );

    \I__10611\ : LocalMux
    port map (
            O => \N__45416\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__10610\ : InMux
    port map (
            O => \N__45413\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__10609\ : InMux
    port map (
            O => \N__45410\,
            I => \N__45403\
        );

    \I__10608\ : InMux
    port map (
            O => \N__45409\,
            I => \N__45403\
        );

    \I__10607\ : InMux
    port map (
            O => \N__45408\,
            I => \N__45400\
        );

    \I__10606\ : LocalMux
    port map (
            O => \N__45403\,
            I => \N__45397\
        );

    \I__10605\ : LocalMux
    port map (
            O => \N__45400\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__10604\ : Odrv4
    port map (
            O => \N__45397\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__10603\ : InMux
    port map (
            O => \N__45392\,
            I => \N__45389\
        );

    \I__10602\ : LocalMux
    port map (
            O => \N__45389\,
            I => \N__45386\
        );

    \I__10601\ : Span4Mux_h
    port map (
            O => \N__45386\,
            I => \N__45383\
        );

    \I__10600\ : Odrv4
    port map (
            O => \N__45383\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__10599\ : InMux
    port map (
            O => \N__45380\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__10598\ : InMux
    port map (
            O => \N__45377\,
            I => \N__45371\
        );

    \I__10597\ : InMux
    port map (
            O => \N__45376\,
            I => \N__45371\
        );

    \I__10596\ : LocalMux
    port map (
            O => \N__45371\,
            I => \N__45367\
        );

    \I__10595\ : InMux
    port map (
            O => \N__45370\,
            I => \N__45364\
        );

    \I__10594\ : Span4Mux_v
    port map (
            O => \N__45367\,
            I => \N__45361\
        );

    \I__10593\ : LocalMux
    port map (
            O => \N__45364\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__10592\ : Odrv4
    port map (
            O => \N__45361\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__10591\ : InMux
    port map (
            O => \N__45356\,
            I => \N__45353\
        );

    \I__10590\ : LocalMux
    port map (
            O => \N__45353\,
            I => \N__45350\
        );

    \I__10589\ : Span4Mux_h
    port map (
            O => \N__45350\,
            I => \N__45347\
        );

    \I__10588\ : Odrv4
    port map (
            O => \N__45347\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__10587\ : InMux
    port map (
            O => \N__45344\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__10586\ : InMux
    port map (
            O => \N__45341\,
            I => \N__45337\
        );

    \I__10585\ : CascadeMux
    port map (
            O => \N__45340\,
            I => \N__45333\
        );

    \I__10584\ : LocalMux
    port map (
            O => \N__45337\,
            I => \N__45330\
        );

    \I__10583\ : InMux
    port map (
            O => \N__45336\,
            I => \N__45327\
        );

    \I__10582\ : InMux
    port map (
            O => \N__45333\,
            I => \N__45324\
        );

    \I__10581\ : Odrv4
    port map (
            O => \N__45330\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__10580\ : LocalMux
    port map (
            O => \N__45327\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__10579\ : LocalMux
    port map (
            O => \N__45324\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__10578\ : InMux
    port map (
            O => \N__45317\,
            I => \N__45314\
        );

    \I__10577\ : LocalMux
    port map (
            O => \N__45314\,
            I => \N__45311\
        );

    \I__10576\ : Span4Mux_h
    port map (
            O => \N__45311\,
            I => \N__45308\
        );

    \I__10575\ : Odrv4
    port map (
            O => \N__45308\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__10574\ : InMux
    port map (
            O => \N__45305\,
            I => \bfn_18_16_0_\
        );

    \I__10573\ : InMux
    port map (
            O => \N__45302\,
            I => \N__45299\
        );

    \I__10572\ : LocalMux
    port map (
            O => \N__45299\,
            I => \N__45294\
        );

    \I__10571\ : InMux
    port map (
            O => \N__45298\,
            I => \N__45291\
        );

    \I__10570\ : InMux
    port map (
            O => \N__45297\,
            I => \N__45288\
        );

    \I__10569\ : Odrv4
    port map (
            O => \N__45294\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__10568\ : LocalMux
    port map (
            O => \N__45291\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__10567\ : LocalMux
    port map (
            O => \N__45288\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__10566\ : InMux
    port map (
            O => \N__45281\,
            I => \N__45278\
        );

    \I__10565\ : LocalMux
    port map (
            O => \N__45278\,
            I => \N__45274\
        );

    \I__10564\ : InMux
    port map (
            O => \N__45277\,
            I => \N__45271\
        );

    \I__10563\ : Span4Mux_v
    port map (
            O => \N__45274\,
            I => \N__45266\
        );

    \I__10562\ : LocalMux
    port map (
            O => \N__45271\,
            I => \N__45266\
        );

    \I__10561\ : Odrv4
    port map (
            O => \N__45266\,
            I => \delay_measurement_inst.elapsed_time_tr_12\
        );

    \I__10560\ : InMux
    port map (
            O => \N__45263\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__10559\ : CascadeMux
    port map (
            O => \N__45260\,
            I => \N__45256\
        );

    \I__10558\ : CascadeMux
    port map (
            O => \N__45259\,
            I => \N__45253\
        );

    \I__10557\ : InMux
    port map (
            O => \N__45256\,
            I => \N__45247\
        );

    \I__10556\ : InMux
    port map (
            O => \N__45253\,
            I => \N__45247\
        );

    \I__10555\ : InMux
    port map (
            O => \N__45252\,
            I => \N__45244\
        );

    \I__10554\ : LocalMux
    port map (
            O => \N__45247\,
            I => \N__45241\
        );

    \I__10553\ : LocalMux
    port map (
            O => \N__45244\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__10552\ : Odrv4
    port map (
            O => \N__45241\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__10551\ : InMux
    port map (
            O => \N__45236\,
            I => \N__45232\
        );

    \I__10550\ : CascadeMux
    port map (
            O => \N__45235\,
            I => \N__45229\
        );

    \I__10549\ : LocalMux
    port map (
            O => \N__45232\,
            I => \N__45226\
        );

    \I__10548\ : InMux
    port map (
            O => \N__45229\,
            I => \N__45223\
        );

    \I__10547\ : Span4Mux_h
    port map (
            O => \N__45226\,
            I => \N__45220\
        );

    \I__10546\ : LocalMux
    port map (
            O => \N__45223\,
            I => \N__45217\
        );

    \I__10545\ : Odrv4
    port map (
            O => \N__45220\,
            I => \delay_measurement_inst.elapsed_time_tr_13\
        );

    \I__10544\ : Odrv4
    port map (
            O => \N__45217\,
            I => \delay_measurement_inst.elapsed_time_tr_13\
        );

    \I__10543\ : InMux
    port map (
            O => \N__45212\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__10542\ : CascadeMux
    port map (
            O => \N__45209\,
            I => \N__45205\
        );

    \I__10541\ : CascadeMux
    port map (
            O => \N__45208\,
            I => \N__45202\
        );

    \I__10540\ : InMux
    port map (
            O => \N__45205\,
            I => \N__45196\
        );

    \I__10539\ : InMux
    port map (
            O => \N__45202\,
            I => \N__45196\
        );

    \I__10538\ : InMux
    port map (
            O => \N__45201\,
            I => \N__45193\
        );

    \I__10537\ : LocalMux
    port map (
            O => \N__45196\,
            I => \N__45190\
        );

    \I__10536\ : LocalMux
    port map (
            O => \N__45193\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__10535\ : Odrv4
    port map (
            O => \N__45190\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__10534\ : InMux
    port map (
            O => \N__45185\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__10533\ : InMux
    port map (
            O => \N__45182\,
            I => \N__45176\
        );

    \I__10532\ : InMux
    port map (
            O => \N__45181\,
            I => \N__45176\
        );

    \I__10531\ : LocalMux
    port map (
            O => \N__45176\,
            I => \N__45172\
        );

    \I__10530\ : InMux
    port map (
            O => \N__45175\,
            I => \N__45169\
        );

    \I__10529\ : Span4Mux_h
    port map (
            O => \N__45172\,
            I => \N__45166\
        );

    \I__10528\ : LocalMux
    port map (
            O => \N__45169\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__10527\ : Odrv4
    port map (
            O => \N__45166\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__10526\ : InMux
    port map (
            O => \N__45161\,
            I => \N__45156\
        );

    \I__10525\ : CascadeMux
    port map (
            O => \N__45160\,
            I => \N__45150\
        );

    \I__10524\ : InMux
    port map (
            O => \N__45159\,
            I => \N__45147\
        );

    \I__10523\ : LocalMux
    port map (
            O => \N__45156\,
            I => \N__45144\
        );

    \I__10522\ : InMux
    port map (
            O => \N__45155\,
            I => \N__45139\
        );

    \I__10521\ : InMux
    port map (
            O => \N__45154\,
            I => \N__45139\
        );

    \I__10520\ : InMux
    port map (
            O => \N__45153\,
            I => \N__45134\
        );

    \I__10519\ : InMux
    port map (
            O => \N__45150\,
            I => \N__45134\
        );

    \I__10518\ : LocalMux
    port map (
            O => \N__45147\,
            I => \N__45131\
        );

    \I__10517\ : Span4Mux_v
    port map (
            O => \N__45144\,
            I => \N__45128\
        );

    \I__10516\ : LocalMux
    port map (
            O => \N__45139\,
            I => \N__45125\
        );

    \I__10515\ : LocalMux
    port map (
            O => \N__45134\,
            I => \N__45122\
        );

    \I__10514\ : Span4Mux_v
    port map (
            O => \N__45131\,
            I => \N__45117\
        );

    \I__10513\ : Span4Mux_h
    port map (
            O => \N__45128\,
            I => \N__45117\
        );

    \I__10512\ : Span4Mux_h
    port map (
            O => \N__45125\,
            I => \N__45114\
        );

    \I__10511\ : Span4Mux_h
    port map (
            O => \N__45122\,
            I => \N__45111\
        );

    \I__10510\ : Odrv4
    port map (
            O => \N__45117\,
            I => \delay_measurement_inst.elapsed_time_tr_15\
        );

    \I__10509\ : Odrv4
    port map (
            O => \N__45114\,
            I => \delay_measurement_inst.elapsed_time_tr_15\
        );

    \I__10508\ : Odrv4
    port map (
            O => \N__45111\,
            I => \delay_measurement_inst.elapsed_time_tr_15\
        );

    \I__10507\ : InMux
    port map (
            O => \N__45104\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__10506\ : InMux
    port map (
            O => \N__45101\,
            I => \N__45095\
        );

    \I__10505\ : InMux
    port map (
            O => \N__45100\,
            I => \N__45095\
        );

    \I__10504\ : LocalMux
    port map (
            O => \N__45095\,
            I => \N__45091\
        );

    \I__10503\ : InMux
    port map (
            O => \N__45094\,
            I => \N__45088\
        );

    \I__10502\ : Span4Mux_h
    port map (
            O => \N__45091\,
            I => \N__45085\
        );

    \I__10501\ : LocalMux
    port map (
            O => \N__45088\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__10500\ : Odrv4
    port map (
            O => \N__45085\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__10499\ : InMux
    port map (
            O => \N__45080\,
            I => \N__45077\
        );

    \I__10498\ : LocalMux
    port map (
            O => \N__45077\,
            I => \N__45072\
        );

    \I__10497\ : InMux
    port map (
            O => \N__45076\,
            I => \N__45067\
        );

    \I__10496\ : InMux
    port map (
            O => \N__45075\,
            I => \N__45067\
        );

    \I__10495\ : Odrv4
    port map (
            O => \N__45072\,
            I => \delay_measurement_inst.elapsed_time_tr_16\
        );

    \I__10494\ : LocalMux
    port map (
            O => \N__45067\,
            I => \delay_measurement_inst.elapsed_time_tr_16\
        );

    \I__10493\ : InMux
    port map (
            O => \N__45062\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__10492\ : CascadeMux
    port map (
            O => \N__45059\,
            I => \N__45056\
        );

    \I__10491\ : InMux
    port map (
            O => \N__45056\,
            I => \N__45052\
        );

    \I__10490\ : InMux
    port map (
            O => \N__45055\,
            I => \N__45048\
        );

    \I__10489\ : LocalMux
    port map (
            O => \N__45052\,
            I => \N__45045\
        );

    \I__10488\ : InMux
    port map (
            O => \N__45051\,
            I => \N__45042\
        );

    \I__10487\ : LocalMux
    port map (
            O => \N__45048\,
            I => \N__45039\
        );

    \I__10486\ : Span4Mux_h
    port map (
            O => \N__45045\,
            I => \N__45036\
        );

    \I__10485\ : LocalMux
    port map (
            O => \N__45042\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__10484\ : Odrv4
    port map (
            O => \N__45039\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__10483\ : Odrv4
    port map (
            O => \N__45036\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__10482\ : InMux
    port map (
            O => \N__45029\,
            I => \N__45026\
        );

    \I__10481\ : LocalMux
    port map (
            O => \N__45026\,
            I => \N__45021\
        );

    \I__10480\ : InMux
    port map (
            O => \N__45025\,
            I => \N__45018\
        );

    \I__10479\ : InMux
    port map (
            O => \N__45024\,
            I => \N__45015\
        );

    \I__10478\ : Odrv4
    port map (
            O => \N__45021\,
            I => \delay_measurement_inst.elapsed_time_tr_17\
        );

    \I__10477\ : LocalMux
    port map (
            O => \N__45018\,
            I => \delay_measurement_inst.elapsed_time_tr_17\
        );

    \I__10476\ : LocalMux
    port map (
            O => \N__45015\,
            I => \delay_measurement_inst.elapsed_time_tr_17\
        );

    \I__10475\ : InMux
    port map (
            O => \N__45008\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__10474\ : CascadeMux
    port map (
            O => \N__45005\,
            I => \N__45001\
        );

    \I__10473\ : CascadeMux
    port map (
            O => \N__45004\,
            I => \N__44998\
        );

    \I__10472\ : InMux
    port map (
            O => \N__45001\,
            I => \N__44993\
        );

    \I__10471\ : InMux
    port map (
            O => \N__44998\,
            I => \N__44993\
        );

    \I__10470\ : LocalMux
    port map (
            O => \N__44993\,
            I => \N__44989\
        );

    \I__10469\ : InMux
    port map (
            O => \N__44992\,
            I => \N__44986\
        );

    \I__10468\ : Span4Mux_v
    port map (
            O => \N__44989\,
            I => \N__44983\
        );

    \I__10467\ : LocalMux
    port map (
            O => \N__44986\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__10466\ : Odrv4
    port map (
            O => \N__44983\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__10465\ : InMux
    port map (
            O => \N__44978\,
            I => \N__44975\
        );

    \I__10464\ : LocalMux
    port map (
            O => \N__44975\,
            I => \N__44970\
        );

    \I__10463\ : InMux
    port map (
            O => \N__44974\,
            I => \N__44965\
        );

    \I__10462\ : InMux
    port map (
            O => \N__44973\,
            I => \N__44965\
        );

    \I__10461\ : Odrv4
    port map (
            O => \N__44970\,
            I => \delay_measurement_inst.elapsed_time_tr_18\
        );

    \I__10460\ : LocalMux
    port map (
            O => \N__44965\,
            I => \delay_measurement_inst.elapsed_time_tr_18\
        );

    \I__10459\ : InMux
    port map (
            O => \N__44960\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__10458\ : InMux
    port map (
            O => \N__44957\,
            I => \N__44954\
        );

    \I__10457\ : LocalMux
    port map (
            O => \N__44954\,
            I => \N__44950\
        );

    \I__10456\ : CascadeMux
    port map (
            O => \N__44953\,
            I => \N__44946\
        );

    \I__10455\ : Span4Mux_h
    port map (
            O => \N__44950\,
            I => \N__44943\
        );

    \I__10454\ : InMux
    port map (
            O => \N__44949\,
            I => \N__44940\
        );

    \I__10453\ : InMux
    port map (
            O => \N__44946\,
            I => \N__44937\
        );

    \I__10452\ : Odrv4
    port map (
            O => \N__44943\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__10451\ : LocalMux
    port map (
            O => \N__44940\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__10450\ : LocalMux
    port map (
            O => \N__44937\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__10449\ : InMux
    port map (
            O => \N__44930\,
            I => \N__44927\
        );

    \I__10448\ : LocalMux
    port map (
            O => \N__44927\,
            I => \N__44922\
        );

    \I__10447\ : CascadeMux
    port map (
            O => \N__44926\,
            I => \N__44919\
        );

    \I__10446\ : CascadeMux
    port map (
            O => \N__44925\,
            I => \N__44916\
        );

    \I__10445\ : Span4Mux_h
    port map (
            O => \N__44922\,
            I => \N__44913\
        );

    \I__10444\ : InMux
    port map (
            O => \N__44919\,
            I => \N__44910\
        );

    \I__10443\ : InMux
    port map (
            O => \N__44916\,
            I => \N__44907\
        );

    \I__10442\ : Odrv4
    port map (
            O => \N__44913\,
            I => \delay_measurement_inst.elapsed_time_tr_19\
        );

    \I__10441\ : LocalMux
    port map (
            O => \N__44910\,
            I => \delay_measurement_inst.elapsed_time_tr_19\
        );

    \I__10440\ : LocalMux
    port map (
            O => \N__44907\,
            I => \delay_measurement_inst.elapsed_time_tr_19\
        );

    \I__10439\ : InMux
    port map (
            O => \N__44900\,
            I => \bfn_18_15_0_\
        );

    \I__10438\ : InMux
    port map (
            O => \N__44897\,
            I => \N__44894\
        );

    \I__10437\ : LocalMux
    port map (
            O => \N__44894\,
            I => \N__44890\
        );

    \I__10436\ : InMux
    port map (
            O => \N__44893\,
            I => \N__44886\
        );

    \I__10435\ : Span4Mux_v
    port map (
            O => \N__44890\,
            I => \N__44883\
        );

    \I__10434\ : InMux
    port map (
            O => \N__44889\,
            I => \N__44880\
        );

    \I__10433\ : LocalMux
    port map (
            O => \N__44886\,
            I => \N__44877\
        );

    \I__10432\ : Odrv4
    port map (
            O => \N__44883\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__10431\ : LocalMux
    port map (
            O => \N__44880\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__10430\ : Odrv4
    port map (
            O => \N__44877\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__10429\ : InMux
    port map (
            O => \N__44870\,
            I => \N__44867\
        );

    \I__10428\ : LocalMux
    port map (
            O => \N__44867\,
            I => \N__44862\
        );

    \I__10427\ : InMux
    port map (
            O => \N__44866\,
            I => \N__44859\
        );

    \I__10426\ : InMux
    port map (
            O => \N__44865\,
            I => \N__44856\
        );

    \I__10425\ : Span4Mux_v
    port map (
            O => \N__44862\,
            I => \N__44851\
        );

    \I__10424\ : LocalMux
    port map (
            O => \N__44859\,
            I => \N__44851\
        );

    \I__10423\ : LocalMux
    port map (
            O => \N__44856\,
            I => \delay_measurement_inst.elapsed_time_tr_4\
        );

    \I__10422\ : Odrv4
    port map (
            O => \N__44851\,
            I => \delay_measurement_inst.elapsed_time_tr_4\
        );

    \I__10421\ : InMux
    port map (
            O => \N__44846\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__10420\ : CascadeMux
    port map (
            O => \N__44843\,
            I => \N__44839\
        );

    \I__10419\ : CascadeMux
    port map (
            O => \N__44842\,
            I => \N__44836\
        );

    \I__10418\ : InMux
    port map (
            O => \N__44839\,
            I => \N__44830\
        );

    \I__10417\ : InMux
    port map (
            O => \N__44836\,
            I => \N__44830\
        );

    \I__10416\ : InMux
    port map (
            O => \N__44835\,
            I => \N__44827\
        );

    \I__10415\ : LocalMux
    port map (
            O => \N__44830\,
            I => \N__44824\
        );

    \I__10414\ : LocalMux
    port map (
            O => \N__44827\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__10413\ : Odrv4
    port map (
            O => \N__44824\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__10412\ : CascadeMux
    port map (
            O => \N__44819\,
            I => \N__44816\
        );

    \I__10411\ : InMux
    port map (
            O => \N__44816\,
            I => \N__44813\
        );

    \I__10410\ : LocalMux
    port map (
            O => \N__44813\,
            I => \N__44808\
        );

    \I__10409\ : InMux
    port map (
            O => \N__44812\,
            I => \N__44803\
        );

    \I__10408\ : InMux
    port map (
            O => \N__44811\,
            I => \N__44803\
        );

    \I__10407\ : Span4Mux_h
    port map (
            O => \N__44808\,
            I => \N__44800\
        );

    \I__10406\ : LocalMux
    port map (
            O => \N__44803\,
            I => \N__44797\
        );

    \I__10405\ : Odrv4
    port map (
            O => \N__44800\,
            I => \delay_measurement_inst.elapsed_time_tr_5\
        );

    \I__10404\ : Odrv12
    port map (
            O => \N__44797\,
            I => \delay_measurement_inst.elapsed_time_tr_5\
        );

    \I__10403\ : InMux
    port map (
            O => \N__44792\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__10402\ : CascadeMux
    port map (
            O => \N__44789\,
            I => \N__44785\
        );

    \I__10401\ : CascadeMux
    port map (
            O => \N__44788\,
            I => \N__44782\
        );

    \I__10400\ : InMux
    port map (
            O => \N__44785\,
            I => \N__44776\
        );

    \I__10399\ : InMux
    port map (
            O => \N__44782\,
            I => \N__44776\
        );

    \I__10398\ : InMux
    port map (
            O => \N__44781\,
            I => \N__44773\
        );

    \I__10397\ : LocalMux
    port map (
            O => \N__44776\,
            I => \N__44770\
        );

    \I__10396\ : LocalMux
    port map (
            O => \N__44773\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__10395\ : Odrv4
    port map (
            O => \N__44770\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__10394\ : InMux
    port map (
            O => \N__44765\,
            I => \N__44762\
        );

    \I__10393\ : LocalMux
    port map (
            O => \N__44762\,
            I => \N__44757\
        );

    \I__10392\ : InMux
    port map (
            O => \N__44761\,
            I => \N__44752\
        );

    \I__10391\ : InMux
    port map (
            O => \N__44760\,
            I => \N__44752\
        );

    \I__10390\ : Span4Mux_h
    port map (
            O => \N__44757\,
            I => \N__44749\
        );

    \I__10389\ : LocalMux
    port map (
            O => \N__44752\,
            I => \N__44746\
        );

    \I__10388\ : Odrv4
    port map (
            O => \N__44749\,
            I => \delay_measurement_inst.elapsed_time_tr_6\
        );

    \I__10387\ : Odrv4
    port map (
            O => \N__44746\,
            I => \delay_measurement_inst.elapsed_time_tr_6\
        );

    \I__10386\ : InMux
    port map (
            O => \N__44741\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__10385\ : InMux
    port map (
            O => \N__44738\,
            I => \N__44732\
        );

    \I__10384\ : InMux
    port map (
            O => \N__44737\,
            I => \N__44732\
        );

    \I__10383\ : LocalMux
    port map (
            O => \N__44732\,
            I => \N__44728\
        );

    \I__10382\ : InMux
    port map (
            O => \N__44731\,
            I => \N__44725\
        );

    \I__10381\ : Span4Mux_h
    port map (
            O => \N__44728\,
            I => \N__44722\
        );

    \I__10380\ : LocalMux
    port map (
            O => \N__44725\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__10379\ : Odrv4
    port map (
            O => \N__44722\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__10378\ : InMux
    port map (
            O => \N__44717\,
            I => \N__44712\
        );

    \I__10377\ : InMux
    port map (
            O => \N__44716\,
            I => \N__44709\
        );

    \I__10376\ : InMux
    port map (
            O => \N__44715\,
            I => \N__44706\
        );

    \I__10375\ : LocalMux
    port map (
            O => \N__44712\,
            I => \N__44701\
        );

    \I__10374\ : LocalMux
    port map (
            O => \N__44709\,
            I => \N__44701\
        );

    \I__10373\ : LocalMux
    port map (
            O => \N__44706\,
            I => \N__44698\
        );

    \I__10372\ : Span4Mux_h
    port map (
            O => \N__44701\,
            I => \N__44695\
        );

    \I__10371\ : Span4Mux_h
    port map (
            O => \N__44698\,
            I => \N__44692\
        );

    \I__10370\ : Odrv4
    port map (
            O => \N__44695\,
            I => \delay_measurement_inst.elapsed_time_tr_7\
        );

    \I__10369\ : Odrv4
    port map (
            O => \N__44692\,
            I => \delay_measurement_inst.elapsed_time_tr_7\
        );

    \I__10368\ : InMux
    port map (
            O => \N__44687\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__10367\ : InMux
    port map (
            O => \N__44684\,
            I => \N__44678\
        );

    \I__10366\ : InMux
    port map (
            O => \N__44683\,
            I => \N__44678\
        );

    \I__10365\ : LocalMux
    port map (
            O => \N__44678\,
            I => \N__44674\
        );

    \I__10364\ : InMux
    port map (
            O => \N__44677\,
            I => \N__44671\
        );

    \I__10363\ : Span4Mux_h
    port map (
            O => \N__44674\,
            I => \N__44668\
        );

    \I__10362\ : LocalMux
    port map (
            O => \N__44671\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__10361\ : Odrv4
    port map (
            O => \N__44668\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__10360\ : InMux
    port map (
            O => \N__44663\,
            I => \N__44659\
        );

    \I__10359\ : InMux
    port map (
            O => \N__44662\,
            I => \N__44656\
        );

    \I__10358\ : LocalMux
    port map (
            O => \N__44659\,
            I => \N__44652\
        );

    \I__10357\ : LocalMux
    port map (
            O => \N__44656\,
            I => \N__44649\
        );

    \I__10356\ : InMux
    port map (
            O => \N__44655\,
            I => \N__44646\
        );

    \I__10355\ : Span4Mux_v
    port map (
            O => \N__44652\,
            I => \N__44639\
        );

    \I__10354\ : Span4Mux_v
    port map (
            O => \N__44649\,
            I => \N__44639\
        );

    \I__10353\ : LocalMux
    port map (
            O => \N__44646\,
            I => \N__44639\
        );

    \I__10352\ : Odrv4
    port map (
            O => \N__44639\,
            I => \delay_measurement_inst.elapsed_time_tr_8\
        );

    \I__10351\ : InMux
    port map (
            O => \N__44636\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__10350\ : CascadeMux
    port map (
            O => \N__44633\,
            I => \N__44630\
        );

    \I__10349\ : InMux
    port map (
            O => \N__44630\,
            I => \N__44626\
        );

    \I__10348\ : InMux
    port map (
            O => \N__44629\,
            I => \N__44622\
        );

    \I__10347\ : LocalMux
    port map (
            O => \N__44626\,
            I => \N__44619\
        );

    \I__10346\ : InMux
    port map (
            O => \N__44625\,
            I => \N__44616\
        );

    \I__10345\ : LocalMux
    port map (
            O => \N__44622\,
            I => \N__44613\
        );

    \I__10344\ : Span4Mux_h
    port map (
            O => \N__44619\,
            I => \N__44610\
        );

    \I__10343\ : LocalMux
    port map (
            O => \N__44616\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__10342\ : Odrv4
    port map (
            O => \N__44613\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__10341\ : Odrv4
    port map (
            O => \N__44610\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__10340\ : InMux
    port map (
            O => \N__44603\,
            I => \N__44598\
        );

    \I__10339\ : InMux
    port map (
            O => \N__44602\,
            I => \N__44595\
        );

    \I__10338\ : CascadeMux
    port map (
            O => \N__44601\,
            I => \N__44591\
        );

    \I__10337\ : LocalMux
    port map (
            O => \N__44598\,
            I => \N__44586\
        );

    \I__10336\ : LocalMux
    port map (
            O => \N__44595\,
            I => \N__44586\
        );

    \I__10335\ : InMux
    port map (
            O => \N__44594\,
            I => \N__44581\
        );

    \I__10334\ : InMux
    port map (
            O => \N__44591\,
            I => \N__44581\
        );

    \I__10333\ : Span12Mux_v
    port map (
            O => \N__44586\,
            I => \N__44576\
        );

    \I__10332\ : LocalMux
    port map (
            O => \N__44581\,
            I => \N__44576\
        );

    \I__10331\ : Odrv12
    port map (
            O => \N__44576\,
            I => \delay_measurement_inst.elapsed_time_tr_9\
        );

    \I__10330\ : InMux
    port map (
            O => \N__44573\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__10329\ : CascadeMux
    port map (
            O => \N__44570\,
            I => \N__44566\
        );

    \I__10328\ : CascadeMux
    port map (
            O => \N__44569\,
            I => \N__44563\
        );

    \I__10327\ : InMux
    port map (
            O => \N__44566\,
            I => \N__44558\
        );

    \I__10326\ : InMux
    port map (
            O => \N__44563\,
            I => \N__44558\
        );

    \I__10325\ : LocalMux
    port map (
            O => \N__44558\,
            I => \N__44554\
        );

    \I__10324\ : InMux
    port map (
            O => \N__44557\,
            I => \N__44551\
        );

    \I__10323\ : Span4Mux_v
    port map (
            O => \N__44554\,
            I => \N__44548\
        );

    \I__10322\ : LocalMux
    port map (
            O => \N__44551\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__10321\ : Odrv4
    port map (
            O => \N__44548\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__10320\ : InMux
    port map (
            O => \N__44543\,
            I => \N__44539\
        );

    \I__10319\ : InMux
    port map (
            O => \N__44542\,
            I => \N__44536\
        );

    \I__10318\ : LocalMux
    port map (
            O => \N__44539\,
            I => \N__44533\
        );

    \I__10317\ : LocalMux
    port map (
            O => \N__44536\,
            I => \N__44530\
        );

    \I__10316\ : Span4Mux_h
    port map (
            O => \N__44533\,
            I => \N__44527\
        );

    \I__10315\ : Span4Mux_h
    port map (
            O => \N__44530\,
            I => \N__44524\
        );

    \I__10314\ : Odrv4
    port map (
            O => \N__44527\,
            I => \delay_measurement_inst.elapsed_time_tr_10\
        );

    \I__10313\ : Odrv4
    port map (
            O => \N__44524\,
            I => \delay_measurement_inst.elapsed_time_tr_10\
        );

    \I__10312\ : InMux
    port map (
            O => \N__44519\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__10311\ : InMux
    port map (
            O => \N__44516\,
            I => \N__44512\
        );

    \I__10310\ : CascadeMux
    port map (
            O => \N__44515\,
            I => \N__44508\
        );

    \I__10309\ : LocalMux
    port map (
            O => \N__44512\,
            I => \N__44505\
        );

    \I__10308\ : InMux
    port map (
            O => \N__44511\,
            I => \N__44502\
        );

    \I__10307\ : InMux
    port map (
            O => \N__44508\,
            I => \N__44499\
        );

    \I__10306\ : Odrv4
    port map (
            O => \N__44505\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__10305\ : LocalMux
    port map (
            O => \N__44502\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__10304\ : LocalMux
    port map (
            O => \N__44499\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__10303\ : InMux
    port map (
            O => \N__44492\,
            I => \N__44489\
        );

    \I__10302\ : LocalMux
    port map (
            O => \N__44489\,
            I => \N__44485\
        );

    \I__10301\ : InMux
    port map (
            O => \N__44488\,
            I => \N__44482\
        );

    \I__10300\ : Span4Mux_v
    port map (
            O => \N__44485\,
            I => \N__44477\
        );

    \I__10299\ : LocalMux
    port map (
            O => \N__44482\,
            I => \N__44477\
        );

    \I__10298\ : Odrv4
    port map (
            O => \N__44477\,
            I => \delay_measurement_inst.elapsed_time_tr_11\
        );

    \I__10297\ : InMux
    port map (
            O => \N__44474\,
            I => \bfn_18_14_0_\
        );

    \I__10296\ : CascadeMux
    port map (
            O => \N__44471\,
            I => \N__44468\
        );

    \I__10295\ : InMux
    port map (
            O => \N__44468\,
            I => \N__44465\
        );

    \I__10294\ : LocalMux
    port map (
            O => \N__44465\,
            I => \N__44462\
        );

    \I__10293\ : Span4Mux_v
    port map (
            O => \N__44462\,
            I => \N__44459\
        );

    \I__10292\ : Span4Mux_h
    port map (
            O => \N__44459\,
            I => \N__44456\
        );

    \I__10291\ : Odrv4
    port map (
            O => \N__44456\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_16\
        );

    \I__10290\ : CEMux
    port map (
            O => \N__44453\,
            I => \N__44450\
        );

    \I__10289\ : LocalMux
    port map (
            O => \N__44450\,
            I => \N__44446\
        );

    \I__10288\ : CEMux
    port map (
            O => \N__44449\,
            I => \N__44441\
        );

    \I__10287\ : Span4Mux_v
    port map (
            O => \N__44446\,
            I => \N__44438\
        );

    \I__10286\ : CEMux
    port map (
            O => \N__44445\,
            I => \N__44435\
        );

    \I__10285\ : CEMux
    port map (
            O => \N__44444\,
            I => \N__44432\
        );

    \I__10284\ : LocalMux
    port map (
            O => \N__44441\,
            I => \N__44429\
        );

    \I__10283\ : Span4Mux_h
    port map (
            O => \N__44438\,
            I => \N__44424\
        );

    \I__10282\ : LocalMux
    port map (
            O => \N__44435\,
            I => \N__44424\
        );

    \I__10281\ : LocalMux
    port map (
            O => \N__44432\,
            I => \N__44421\
        );

    \I__10280\ : Span4Mux_v
    port map (
            O => \N__44429\,
            I => \N__44418\
        );

    \I__10279\ : Span4Mux_v
    port map (
            O => \N__44424\,
            I => \N__44414\
        );

    \I__10278\ : Span4Mux_h
    port map (
            O => \N__44421\,
            I => \N__44411\
        );

    \I__10277\ : Span4Mux_h
    port map (
            O => \N__44418\,
            I => \N__44408\
        );

    \I__10276\ : CEMux
    port map (
            O => \N__44417\,
            I => \N__44405\
        );

    \I__10275\ : Span4Mux_v
    port map (
            O => \N__44414\,
            I => \N__44402\
        );

    \I__10274\ : Span4Mux_v
    port map (
            O => \N__44411\,
            I => \N__44399\
        );

    \I__10273\ : Span4Mux_v
    port map (
            O => \N__44408\,
            I => \N__44394\
        );

    \I__10272\ : LocalMux
    port map (
            O => \N__44405\,
            I => \N__44394\
        );

    \I__10271\ : Odrv4
    port map (
            O => \N__44402\,
            I => \phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__10270\ : Odrv4
    port map (
            O => \N__44399\,
            I => \phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__10269\ : Odrv4
    port map (
            O => \N__44394\,
            I => \phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__10268\ : InMux
    port map (
            O => \N__44387\,
            I => \N__44379\
        );

    \I__10267\ : InMux
    port map (
            O => \N__44386\,
            I => \N__44379\
        );

    \I__10266\ : InMux
    port map (
            O => \N__44385\,
            I => \N__44376\
        );

    \I__10265\ : InMux
    port map (
            O => \N__44384\,
            I => \N__44373\
        );

    \I__10264\ : LocalMux
    port map (
            O => \N__44379\,
            I => \N__44370\
        );

    \I__10263\ : LocalMux
    port map (
            O => \N__44376\,
            I => \N__44365\
        );

    \I__10262\ : LocalMux
    port map (
            O => \N__44373\,
            I => \N__44365\
        );

    \I__10261\ : Span4Mux_v
    port map (
            O => \N__44370\,
            I => \N__44362\
        );

    \I__10260\ : Odrv12
    port map (
            O => \N__44365\,
            I => measured_delay_tr_16
        );

    \I__10259\ : Odrv4
    port map (
            O => \N__44362\,
            I => measured_delay_tr_16
        );

    \I__10258\ : CascadeMux
    port map (
            O => \N__44357\,
            I => \N__44354\
        );

    \I__10257\ : InMux
    port map (
            O => \N__44354\,
            I => \N__44351\
        );

    \I__10256\ : LocalMux
    port map (
            O => \N__44351\,
            I => \N__44348\
        );

    \I__10255\ : Span4Mux_h
    port map (
            O => \N__44348\,
            I => \N__44345\
        );

    \I__10254\ : Odrv4
    port map (
            O => \N__44345\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\
        );

    \I__10253\ : InMux
    port map (
            O => \N__44342\,
            I => \N__44338\
        );

    \I__10252\ : InMux
    port map (
            O => \N__44341\,
            I => \N__44335\
        );

    \I__10251\ : LocalMux
    port map (
            O => \N__44338\,
            I => measured_delay_hc_29
        );

    \I__10250\ : LocalMux
    port map (
            O => \N__44335\,
            I => measured_delay_hc_29
        );

    \I__10249\ : InMux
    port map (
            O => \N__44330\,
            I => \N__44326\
        );

    \I__10248\ : InMux
    port map (
            O => \N__44329\,
            I => \N__44323\
        );

    \I__10247\ : LocalMux
    port map (
            O => \N__44326\,
            I => measured_delay_hc_28
        );

    \I__10246\ : LocalMux
    port map (
            O => \N__44323\,
            I => measured_delay_hc_28
        );

    \I__10245\ : CascadeMux
    port map (
            O => \N__44318\,
            I => \N__44314\
        );

    \I__10244\ : InMux
    port map (
            O => \N__44317\,
            I => \N__44311\
        );

    \I__10243\ : InMux
    port map (
            O => \N__44314\,
            I => \N__44308\
        );

    \I__10242\ : LocalMux
    port map (
            O => \N__44311\,
            I => measured_delay_hc_30
        );

    \I__10241\ : LocalMux
    port map (
            O => \N__44308\,
            I => measured_delay_hc_30
        );

    \I__10240\ : InMux
    port map (
            O => \N__44303\,
            I => \N__44299\
        );

    \I__10239\ : InMux
    port map (
            O => \N__44302\,
            I => \N__44296\
        );

    \I__10238\ : LocalMux
    port map (
            O => \N__44299\,
            I => measured_delay_hc_27
        );

    \I__10237\ : LocalMux
    port map (
            O => \N__44296\,
            I => measured_delay_hc_27
        );

    \I__10236\ : InMux
    port map (
            O => \N__44291\,
            I => \N__44288\
        );

    \I__10235\ : LocalMux
    port map (
            O => \N__44288\,
            I => \N__44285\
        );

    \I__10234\ : Odrv4
    port map (
            O => \N__44285\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_4\
        );

    \I__10233\ : InMux
    port map (
            O => \N__44282\,
            I => \N__44278\
        );

    \I__10232\ : InMux
    port map (
            O => \N__44281\,
            I => \N__44275\
        );

    \I__10231\ : LocalMux
    port map (
            O => \N__44278\,
            I => \N__44270\
        );

    \I__10230\ : LocalMux
    port map (
            O => \N__44275\,
            I => \N__44267\
        );

    \I__10229\ : InMux
    port map (
            O => \N__44274\,
            I => \N__44264\
        );

    \I__10228\ : CascadeMux
    port map (
            O => \N__44273\,
            I => \N__44261\
        );

    \I__10227\ : Span4Mux_h
    port map (
            O => \N__44270\,
            I => \N__44257\
        );

    \I__10226\ : Span4Mux_v
    port map (
            O => \N__44267\,
            I => \N__44254\
        );

    \I__10225\ : LocalMux
    port map (
            O => \N__44264\,
            I => \N__44251\
        );

    \I__10224\ : InMux
    port map (
            O => \N__44261\,
            I => \N__44248\
        );

    \I__10223\ : CascadeMux
    port map (
            O => \N__44260\,
            I => \N__44245\
        );

    \I__10222\ : Span4Mux_h
    port map (
            O => \N__44257\,
            I => \N__44236\
        );

    \I__10221\ : Span4Mux_h
    port map (
            O => \N__44254\,
            I => \N__44236\
        );

    \I__10220\ : Span4Mux_v
    port map (
            O => \N__44251\,
            I => \N__44236\
        );

    \I__10219\ : LocalMux
    port map (
            O => \N__44248\,
            I => \N__44236\
        );

    \I__10218\ : InMux
    port map (
            O => \N__44245\,
            I => \N__44233\
        );

    \I__10217\ : Span4Mux_v
    port map (
            O => \N__44236\,
            I => \N__44230\
        );

    \I__10216\ : LocalMux
    port map (
            O => \N__44233\,
            I => measured_delay_hc_13
        );

    \I__10215\ : Odrv4
    port map (
            O => \N__44230\,
            I => measured_delay_hc_13
        );

    \I__10214\ : CascadeMux
    port map (
            O => \N__44225\,
            I => \N__44222\
        );

    \I__10213\ : InMux
    port map (
            O => \N__44222\,
            I => \N__44219\
        );

    \I__10212\ : LocalMux
    port map (
            O => \N__44219\,
            I => \N__44216\
        );

    \I__10211\ : Span4Mux_v
    port map (
            O => \N__44216\,
            I => \N__44213\
        );

    \I__10210\ : Span4Mux_v
    port map (
            O => \N__44213\,
            I => \N__44210\
        );

    \I__10209\ : Odrv4
    port map (
            O => \N__44210\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_13\
        );

    \I__10208\ : CascadeMux
    port map (
            O => \N__44207\,
            I => \N__44201\
        );

    \I__10207\ : InMux
    port map (
            O => \N__44206\,
            I => \N__44189\
        );

    \I__10206\ : InMux
    port map (
            O => \N__44205\,
            I => \N__44189\
        );

    \I__10205\ : InMux
    port map (
            O => \N__44204\,
            I => \N__44189\
        );

    \I__10204\ : InMux
    port map (
            O => \N__44201\,
            I => \N__44189\
        );

    \I__10203\ : CascadeMux
    port map (
            O => \N__44200\,
            I => \N__44174\
        );

    \I__10202\ : CascadeMux
    port map (
            O => \N__44199\,
            I => \N__44170\
        );

    \I__10201\ : CascadeMux
    port map (
            O => \N__44198\,
            I => \N__44161\
        );

    \I__10200\ : LocalMux
    port map (
            O => \N__44189\,
            I => \N__44158\
        );

    \I__10199\ : CascadeMux
    port map (
            O => \N__44188\,
            I => \N__44151\
        );

    \I__10198\ : CascadeMux
    port map (
            O => \N__44187\,
            I => \N__44148\
        );

    \I__10197\ : CascadeMux
    port map (
            O => \N__44186\,
            I => \N__44145\
        );

    \I__10196\ : CascadeMux
    port map (
            O => \N__44185\,
            I => \N__44141\
        );

    \I__10195\ : InMux
    port map (
            O => \N__44184\,
            I => \N__44126\
        );

    \I__10194\ : InMux
    port map (
            O => \N__44183\,
            I => \N__44126\
        );

    \I__10193\ : InMux
    port map (
            O => \N__44182\,
            I => \N__44126\
        );

    \I__10192\ : InMux
    port map (
            O => \N__44181\,
            I => \N__44126\
        );

    \I__10191\ : InMux
    port map (
            O => \N__44180\,
            I => \N__44126\
        );

    \I__10190\ : InMux
    port map (
            O => \N__44179\,
            I => \N__44126\
        );

    \I__10189\ : InMux
    port map (
            O => \N__44178\,
            I => \N__44109\
        );

    \I__10188\ : InMux
    port map (
            O => \N__44177\,
            I => \N__44109\
        );

    \I__10187\ : InMux
    port map (
            O => \N__44174\,
            I => \N__44109\
        );

    \I__10186\ : InMux
    port map (
            O => \N__44173\,
            I => \N__44109\
        );

    \I__10185\ : InMux
    port map (
            O => \N__44170\,
            I => \N__44109\
        );

    \I__10184\ : InMux
    port map (
            O => \N__44169\,
            I => \N__44109\
        );

    \I__10183\ : InMux
    port map (
            O => \N__44168\,
            I => \N__44109\
        );

    \I__10182\ : InMux
    port map (
            O => \N__44167\,
            I => \N__44109\
        );

    \I__10181\ : InMux
    port map (
            O => \N__44166\,
            I => \N__44100\
        );

    \I__10180\ : InMux
    port map (
            O => \N__44165\,
            I => \N__44100\
        );

    \I__10179\ : InMux
    port map (
            O => \N__44164\,
            I => \N__44100\
        );

    \I__10178\ : InMux
    port map (
            O => \N__44161\,
            I => \N__44100\
        );

    \I__10177\ : Span4Mux_v
    port map (
            O => \N__44158\,
            I => \N__44097\
        );

    \I__10176\ : InMux
    port map (
            O => \N__44157\,
            I => \N__44094\
        );

    \I__10175\ : InMux
    port map (
            O => \N__44156\,
            I => \N__44091\
        );

    \I__10174\ : CascadeMux
    port map (
            O => \N__44155\,
            I => \N__44088\
        );

    \I__10173\ : InMux
    port map (
            O => \N__44154\,
            I => \N__44081\
        );

    \I__10172\ : InMux
    port map (
            O => \N__44151\,
            I => \N__44066\
        );

    \I__10171\ : InMux
    port map (
            O => \N__44148\,
            I => \N__44066\
        );

    \I__10170\ : InMux
    port map (
            O => \N__44145\,
            I => \N__44066\
        );

    \I__10169\ : InMux
    port map (
            O => \N__44144\,
            I => \N__44066\
        );

    \I__10168\ : InMux
    port map (
            O => \N__44141\,
            I => \N__44066\
        );

    \I__10167\ : InMux
    port map (
            O => \N__44140\,
            I => \N__44066\
        );

    \I__10166\ : InMux
    port map (
            O => \N__44139\,
            I => \N__44066\
        );

    \I__10165\ : LocalMux
    port map (
            O => \N__44126\,
            I => \N__44063\
        );

    \I__10164\ : LocalMux
    port map (
            O => \N__44109\,
            I => \N__44055\
        );

    \I__10163\ : LocalMux
    port map (
            O => \N__44100\,
            I => \N__44055\
        );

    \I__10162\ : Span4Mux_h
    port map (
            O => \N__44097\,
            I => \N__44052\
        );

    \I__10161\ : LocalMux
    port map (
            O => \N__44094\,
            I => \N__44049\
        );

    \I__10160\ : LocalMux
    port map (
            O => \N__44091\,
            I => \N__44046\
        );

    \I__10159\ : InMux
    port map (
            O => \N__44088\,
            I => \N__44039\
        );

    \I__10158\ : InMux
    port map (
            O => \N__44087\,
            I => \N__44039\
        );

    \I__10157\ : InMux
    port map (
            O => \N__44086\,
            I => \N__44039\
        );

    \I__10156\ : InMux
    port map (
            O => \N__44085\,
            I => \N__44034\
        );

    \I__10155\ : InMux
    port map (
            O => \N__44084\,
            I => \N__44034\
        );

    \I__10154\ : LocalMux
    port map (
            O => \N__44081\,
            I => \N__44031\
        );

    \I__10153\ : LocalMux
    port map (
            O => \N__44066\,
            I => \N__44028\
        );

    \I__10152\ : Span4Mux_h
    port map (
            O => \N__44063\,
            I => \N__44025\
        );

    \I__10151\ : InMux
    port map (
            O => \N__44062\,
            I => \N__44018\
        );

    \I__10150\ : InMux
    port map (
            O => \N__44061\,
            I => \N__44018\
        );

    \I__10149\ : InMux
    port map (
            O => \N__44060\,
            I => \N__44018\
        );

    \I__10148\ : Span4Mux_v
    port map (
            O => \N__44055\,
            I => \N__44014\
        );

    \I__10147\ : Span4Mux_h
    port map (
            O => \N__44052\,
            I => \N__44009\
        );

    \I__10146\ : Span4Mux_h
    port map (
            O => \N__44049\,
            I => \N__44009\
        );

    \I__10145\ : Span4Mux_h
    port map (
            O => \N__44046\,
            I => \N__44006\
        );

    \I__10144\ : LocalMux
    port map (
            O => \N__44039\,
            I => \N__44001\
        );

    \I__10143\ : LocalMux
    port map (
            O => \N__44034\,
            I => \N__44001\
        );

    \I__10142\ : Span4Mux_h
    port map (
            O => \N__44031\,
            I => \N__43998\
        );

    \I__10141\ : Span4Mux_v
    port map (
            O => \N__44028\,
            I => \N__43995\
        );

    \I__10140\ : Span4Mux_v
    port map (
            O => \N__44025\,
            I => \N__43990\
        );

    \I__10139\ : LocalMux
    port map (
            O => \N__44018\,
            I => \N__43990\
        );

    \I__10138\ : InMux
    port map (
            O => \N__44017\,
            I => \N__43987\
        );

    \I__10137\ : Span4Mux_v
    port map (
            O => \N__44014\,
            I => \N__43984\
        );

    \I__10136\ : Span4Mux_v
    port map (
            O => \N__44009\,
            I => \N__43979\
        );

    \I__10135\ : Span4Mux_v
    port map (
            O => \N__44006\,
            I => \N__43979\
        );

    \I__10134\ : Span12Mux_h
    port map (
            O => \N__44001\,
            I => \N__43976\
        );

    \I__10133\ : Span4Mux_h
    port map (
            O => \N__43998\,
            I => \N__43969\
        );

    \I__10132\ : Span4Mux_h
    port map (
            O => \N__43995\,
            I => \N__43969\
        );

    \I__10131\ : Span4Mux_v
    port map (
            O => \N__43990\,
            I => \N__43969\
        );

    \I__10130\ : LocalMux
    port map (
            O => \N__43987\,
            I => measured_delay_hc_31
        );

    \I__10129\ : Odrv4
    port map (
            O => \N__43984\,
            I => measured_delay_hc_31
        );

    \I__10128\ : Odrv4
    port map (
            O => \N__43979\,
            I => measured_delay_hc_31
        );

    \I__10127\ : Odrv12
    port map (
            O => \N__43976\,
            I => measured_delay_hc_31
        );

    \I__10126\ : Odrv4
    port map (
            O => \N__43969\,
            I => measured_delay_hc_31
        );

    \I__10125\ : CascadeMux
    port map (
            O => \N__43958\,
            I => \N__43951\
        );

    \I__10124\ : InMux
    port map (
            O => \N__43957\,
            I => \N__43948\
        );

    \I__10123\ : InMux
    port map (
            O => \N__43956\,
            I => \N__43945\
        );

    \I__10122\ : InMux
    port map (
            O => \N__43955\,
            I => \N__43942\
        );

    \I__10121\ : InMux
    port map (
            O => \N__43954\,
            I => \N__43939\
        );

    \I__10120\ : InMux
    port map (
            O => \N__43951\,
            I => \N__43936\
        );

    \I__10119\ : LocalMux
    port map (
            O => \N__43948\,
            I => \N__43933\
        );

    \I__10118\ : LocalMux
    port map (
            O => \N__43945\,
            I => \N__43930\
        );

    \I__10117\ : LocalMux
    port map (
            O => \N__43942\,
            I => \N__43927\
        );

    \I__10116\ : LocalMux
    port map (
            O => \N__43939\,
            I => \N__43924\
        );

    \I__10115\ : LocalMux
    port map (
            O => \N__43936\,
            I => measured_delay_hc_5
        );

    \I__10114\ : Odrv12
    port map (
            O => \N__43933\,
            I => measured_delay_hc_5
        );

    \I__10113\ : Odrv12
    port map (
            O => \N__43930\,
            I => measured_delay_hc_5
        );

    \I__10112\ : Odrv4
    port map (
            O => \N__43927\,
            I => measured_delay_hc_5
        );

    \I__10111\ : Odrv4
    port map (
            O => \N__43924\,
            I => measured_delay_hc_5
        );

    \I__10110\ : InMux
    port map (
            O => \N__43913\,
            I => \N__43901\
        );

    \I__10109\ : InMux
    port map (
            O => \N__43912\,
            I => \N__43901\
        );

    \I__10108\ : InMux
    port map (
            O => \N__43911\,
            I => \N__43901\
        );

    \I__10107\ : InMux
    port map (
            O => \N__43910\,
            I => \N__43901\
        );

    \I__10106\ : LocalMux
    port map (
            O => \N__43901\,
            I => \N__43889\
        );

    \I__10105\ : InMux
    port map (
            O => \N__43900\,
            I => \N__43880\
        );

    \I__10104\ : InMux
    port map (
            O => \N__43899\,
            I => \N__43880\
        );

    \I__10103\ : InMux
    port map (
            O => \N__43898\,
            I => \N__43880\
        );

    \I__10102\ : InMux
    port map (
            O => \N__43897\,
            I => \N__43875\
        );

    \I__10101\ : InMux
    port map (
            O => \N__43896\,
            I => \N__43864\
        );

    \I__10100\ : InMux
    port map (
            O => \N__43895\,
            I => \N__43864\
        );

    \I__10099\ : InMux
    port map (
            O => \N__43894\,
            I => \N__43864\
        );

    \I__10098\ : InMux
    port map (
            O => \N__43893\,
            I => \N__43864\
        );

    \I__10097\ : InMux
    port map (
            O => \N__43892\,
            I => \N__43864\
        );

    \I__10096\ : Span4Mux_h
    port map (
            O => \N__43889\,
            I => \N__43841\
        );

    \I__10095\ : InMux
    port map (
            O => \N__43888\,
            I => \N__43836\
        );

    \I__10094\ : InMux
    port map (
            O => \N__43887\,
            I => \N__43836\
        );

    \I__10093\ : LocalMux
    port map (
            O => \N__43880\,
            I => \N__43833\
        );

    \I__10092\ : InMux
    port map (
            O => \N__43879\,
            I => \N__43828\
        );

    \I__10091\ : InMux
    port map (
            O => \N__43878\,
            I => \N__43828\
        );

    \I__10090\ : LocalMux
    port map (
            O => \N__43875\,
            I => \N__43824\
        );

    \I__10089\ : LocalMux
    port map (
            O => \N__43864\,
            I => \N__43821\
        );

    \I__10088\ : InMux
    port map (
            O => \N__43863\,
            I => \N__43804\
        );

    \I__10087\ : InMux
    port map (
            O => \N__43862\,
            I => \N__43804\
        );

    \I__10086\ : InMux
    port map (
            O => \N__43861\,
            I => \N__43804\
        );

    \I__10085\ : InMux
    port map (
            O => \N__43860\,
            I => \N__43804\
        );

    \I__10084\ : InMux
    port map (
            O => \N__43859\,
            I => \N__43804\
        );

    \I__10083\ : InMux
    port map (
            O => \N__43858\,
            I => \N__43804\
        );

    \I__10082\ : InMux
    port map (
            O => \N__43857\,
            I => \N__43804\
        );

    \I__10081\ : InMux
    port map (
            O => \N__43856\,
            I => \N__43804\
        );

    \I__10080\ : InMux
    port map (
            O => \N__43855\,
            I => \N__43795\
        );

    \I__10079\ : InMux
    port map (
            O => \N__43854\,
            I => \N__43795\
        );

    \I__10078\ : InMux
    port map (
            O => \N__43853\,
            I => \N__43795\
        );

    \I__10077\ : InMux
    port map (
            O => \N__43852\,
            I => \N__43795\
        );

    \I__10076\ : InMux
    port map (
            O => \N__43851\,
            I => \N__43792\
        );

    \I__10075\ : InMux
    port map (
            O => \N__43850\,
            I => \N__43777\
        );

    \I__10074\ : InMux
    port map (
            O => \N__43849\,
            I => \N__43777\
        );

    \I__10073\ : InMux
    port map (
            O => \N__43848\,
            I => \N__43777\
        );

    \I__10072\ : InMux
    port map (
            O => \N__43847\,
            I => \N__43777\
        );

    \I__10071\ : InMux
    port map (
            O => \N__43846\,
            I => \N__43777\
        );

    \I__10070\ : InMux
    port map (
            O => \N__43845\,
            I => \N__43777\
        );

    \I__10069\ : InMux
    port map (
            O => \N__43844\,
            I => \N__43777\
        );

    \I__10068\ : Span4Mux_h
    port map (
            O => \N__43841\,
            I => \N__43772\
        );

    \I__10067\ : LocalMux
    port map (
            O => \N__43836\,
            I => \N__43772\
        );

    \I__10066\ : Sp12to4
    port map (
            O => \N__43833\,
            I => \N__43767\
        );

    \I__10065\ : LocalMux
    port map (
            O => \N__43828\,
            I => \N__43767\
        );

    \I__10064\ : InMux
    port map (
            O => \N__43827\,
            I => \N__43764\
        );

    \I__10063\ : Span4Mux_h
    port map (
            O => \N__43824\,
            I => \N__43761\
        );

    \I__10062\ : Span12Mux_s11_h
    port map (
            O => \N__43821\,
            I => \N__43754\
        );

    \I__10061\ : LocalMux
    port map (
            O => \N__43804\,
            I => \N__43754\
        );

    \I__10060\ : LocalMux
    port map (
            O => \N__43795\,
            I => \N__43754\
        );

    \I__10059\ : LocalMux
    port map (
            O => \N__43792\,
            I => \N__43749\
        );

    \I__10058\ : LocalMux
    port map (
            O => \N__43777\,
            I => \N__43749\
        );

    \I__10057\ : Span4Mux_h
    port map (
            O => \N__43772\,
            I => \N__43746\
        );

    \I__10056\ : Span12Mux_v
    port map (
            O => \N__43767\,
            I => \N__43741\
        );

    \I__10055\ : LocalMux
    port map (
            O => \N__43764\,
            I => \N__43741\
        );

    \I__10054\ : Odrv4
    port map (
            O => \N__43761\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt31_0\
        );

    \I__10053\ : Odrv12
    port map (
            O => \N__43754\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt31_0\
        );

    \I__10052\ : Odrv12
    port map (
            O => \N__43749\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt31_0\
        );

    \I__10051\ : Odrv4
    port map (
            O => \N__43746\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt31_0\
        );

    \I__10050\ : Odrv12
    port map (
            O => \N__43741\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt31_0\
        );

    \I__10049\ : CascadeMux
    port map (
            O => \N__43730\,
            I => \N__43727\
        );

    \I__10048\ : InMux
    port map (
            O => \N__43727\,
            I => \N__43724\
        );

    \I__10047\ : LocalMux
    port map (
            O => \N__43724\,
            I => \N__43721\
        );

    \I__10046\ : Span4Mux_v
    port map (
            O => \N__43721\,
            I => \N__43718\
        );

    \I__10045\ : Span4Mux_h
    port map (
            O => \N__43718\,
            I => \N__43715\
        );

    \I__10044\ : Odrv4
    port map (
            O => \N__43715\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_5\
        );

    \I__10043\ : CEMux
    port map (
            O => \N__43712\,
            I => \N__43708\
        );

    \I__10042\ : CEMux
    port map (
            O => \N__43711\,
            I => \N__43704\
        );

    \I__10041\ : LocalMux
    port map (
            O => \N__43708\,
            I => \N__43701\
        );

    \I__10040\ : CEMux
    port map (
            O => \N__43707\,
            I => \N__43697\
        );

    \I__10039\ : LocalMux
    port map (
            O => \N__43704\,
            I => \N__43694\
        );

    \I__10038\ : Span4Mux_v
    port map (
            O => \N__43701\,
            I => \N__43691\
        );

    \I__10037\ : CEMux
    port map (
            O => \N__43700\,
            I => \N__43688\
        );

    \I__10036\ : LocalMux
    port map (
            O => \N__43697\,
            I => \N__43684\
        );

    \I__10035\ : Span4Mux_v
    port map (
            O => \N__43694\,
            I => \N__43681\
        );

    \I__10034\ : Span4Mux_h
    port map (
            O => \N__43691\,
            I => \N__43676\
        );

    \I__10033\ : LocalMux
    port map (
            O => \N__43688\,
            I => \N__43676\
        );

    \I__10032\ : CEMux
    port map (
            O => \N__43687\,
            I => \N__43673\
        );

    \I__10031\ : Span4Mux_h
    port map (
            O => \N__43684\,
            I => \N__43670\
        );

    \I__10030\ : Span4Mux_h
    port map (
            O => \N__43681\,
            I => \N__43667\
        );

    \I__10029\ : Span4Mux_v
    port map (
            O => \N__43676\,
            I => \N__43662\
        );

    \I__10028\ : LocalMux
    port map (
            O => \N__43673\,
            I => \N__43662\
        );

    \I__10027\ : Span4Mux_h
    port map (
            O => \N__43670\,
            I => \N__43659\
        );

    \I__10026\ : Span4Mux_v
    port map (
            O => \N__43667\,
            I => \N__43654\
        );

    \I__10025\ : Span4Mux_h
    port map (
            O => \N__43662\,
            I => \N__43654\
        );

    \I__10024\ : Odrv4
    port map (
            O => \N__43659\,
            I => \phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__10023\ : Odrv4
    port map (
            O => \N__43654\,
            I => \phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__10022\ : CascadeMux
    port map (
            O => \N__43649\,
            I => \N__43642\
        );

    \I__10021\ : CascadeMux
    port map (
            O => \N__43648\,
            I => \N__43639\
        );

    \I__10020\ : InMux
    port map (
            O => \N__43647\,
            I => \N__43635\
        );

    \I__10019\ : InMux
    port map (
            O => \N__43646\,
            I => \N__43632\
        );

    \I__10018\ : InMux
    port map (
            O => \N__43645\,
            I => \N__43623\
        );

    \I__10017\ : InMux
    port map (
            O => \N__43642\,
            I => \N__43623\
        );

    \I__10016\ : InMux
    port map (
            O => \N__43639\,
            I => \N__43623\
        );

    \I__10015\ : InMux
    port map (
            O => \N__43638\,
            I => \N__43623\
        );

    \I__10014\ : LocalMux
    port map (
            O => \N__43635\,
            I => \N__43620\
        );

    \I__10013\ : LocalMux
    port map (
            O => \N__43632\,
            I => \N__43612\
        );

    \I__10012\ : LocalMux
    port map (
            O => \N__43623\,
            I => \N__43612\
        );

    \I__10011\ : Span4Mux_h
    port map (
            O => \N__43620\,
            I => \N__43612\
        );

    \I__10010\ : InMux
    port map (
            O => \N__43619\,
            I => \N__43609\
        );

    \I__10009\ : Odrv4
    port map (
            O => \N__43612\,
            I => \delay_measurement_inst.N_410\
        );

    \I__10008\ : LocalMux
    port map (
            O => \N__43609\,
            I => \delay_measurement_inst.N_410\
        );

    \I__10007\ : CascadeMux
    port map (
            O => \N__43604\,
            I => \N__43598\
        );

    \I__10006\ : CascadeMux
    port map (
            O => \N__43603\,
            I => \N__43595\
        );

    \I__10005\ : CascadeMux
    port map (
            O => \N__43602\,
            I => \N__43588\
        );

    \I__10004\ : CascadeMux
    port map (
            O => \N__43601\,
            I => \N__43585\
        );

    \I__10003\ : InMux
    port map (
            O => \N__43598\,
            I => \N__43582\
        );

    \I__10002\ : InMux
    port map (
            O => \N__43595\,
            I => \N__43577\
        );

    \I__10001\ : InMux
    port map (
            O => \N__43594\,
            I => \N__43577\
        );

    \I__10000\ : InMux
    port map (
            O => \N__43593\,
            I => \N__43566\
        );

    \I__9999\ : InMux
    port map (
            O => \N__43592\,
            I => \N__43566\
        );

    \I__9998\ : InMux
    port map (
            O => \N__43591\,
            I => \N__43566\
        );

    \I__9997\ : InMux
    port map (
            O => \N__43588\,
            I => \N__43566\
        );

    \I__9996\ : InMux
    port map (
            O => \N__43585\,
            I => \N__43566\
        );

    \I__9995\ : LocalMux
    port map (
            O => \N__43582\,
            I => \N__43563\
        );

    \I__9994\ : LocalMux
    port map (
            O => \N__43577\,
            I => \N__43560\
        );

    \I__9993\ : LocalMux
    port map (
            O => \N__43566\,
            I => \N__43553\
        );

    \I__9992\ : Span4Mux_h
    port map (
            O => \N__43563\,
            I => \N__43553\
        );

    \I__9991\ : Span4Mux_h
    port map (
            O => \N__43560\,
            I => \N__43553\
        );

    \I__9990\ : Odrv4
    port map (
            O => \N__43553\,
            I => \delay_measurement_inst.N_358\
        );

    \I__9989\ : InMux
    port map (
            O => \N__43550\,
            I => \N__43547\
        );

    \I__9988\ : LocalMux
    port map (
            O => \N__43547\,
            I => \N__43538\
        );

    \I__9987\ : InMux
    port map (
            O => \N__43546\,
            I => \N__43527\
        );

    \I__9986\ : InMux
    port map (
            O => \N__43545\,
            I => \N__43527\
        );

    \I__9985\ : InMux
    port map (
            O => \N__43544\,
            I => \N__43527\
        );

    \I__9984\ : InMux
    port map (
            O => \N__43543\,
            I => \N__43527\
        );

    \I__9983\ : InMux
    port map (
            O => \N__43542\,
            I => \N__43527\
        );

    \I__9982\ : InMux
    port map (
            O => \N__43541\,
            I => \N__43524\
        );

    \I__9981\ : Span4Mux_v
    port map (
            O => \N__43538\,
            I => \N__43520\
        );

    \I__9980\ : LocalMux
    port map (
            O => \N__43527\,
            I => \N__43517\
        );

    \I__9979\ : LocalMux
    port map (
            O => \N__43524\,
            I => \N__43514\
        );

    \I__9978\ : InMux
    port map (
            O => \N__43523\,
            I => \N__43511\
        );

    \I__9977\ : Odrv4
    port map (
            O => \N__43520\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15\
        );

    \I__9976\ : Odrv12
    port map (
            O => \N__43517\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15\
        );

    \I__9975\ : Odrv4
    port map (
            O => \N__43514\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15\
        );

    \I__9974\ : LocalMux
    port map (
            O => \N__43511\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15\
        );

    \I__9973\ : InMux
    port map (
            O => \N__43502\,
            I => \N__43498\
        );

    \I__9972\ : CascadeMux
    port map (
            O => \N__43501\,
            I => \N__43494\
        );

    \I__9971\ : LocalMux
    port map (
            O => \N__43498\,
            I => \N__43491\
        );

    \I__9970\ : InMux
    port map (
            O => \N__43497\,
            I => \N__43488\
        );

    \I__9969\ : InMux
    port map (
            O => \N__43494\,
            I => \N__43485\
        );

    \I__9968\ : Span4Mux_v
    port map (
            O => \N__43491\,
            I => \N__43480\
        );

    \I__9967\ : LocalMux
    port map (
            O => \N__43488\,
            I => \N__43480\
        );

    \I__9966\ : LocalMux
    port map (
            O => \N__43485\,
            I => \N__43477\
        );

    \I__9965\ : Span4Mux_v
    port map (
            O => \N__43480\,
            I => \N__43474\
        );

    \I__9964\ : Span12Mux_h
    port map (
            O => \N__43477\,
            I => \N__43471\
        );

    \I__9963\ : Span4Mux_v
    port map (
            O => \N__43474\,
            I => \N__43468\
        );

    \I__9962\ : Odrv12
    port map (
            O => \N__43471\,
            I => measured_delay_tr_4
        );

    \I__9961\ : Odrv4
    port map (
            O => \N__43468\,
            I => measured_delay_tr_4
        );

    \I__9960\ : CEMux
    port map (
            O => \N__43463\,
            I => \N__43458\
        );

    \I__9959\ : CEMux
    port map (
            O => \N__43462\,
            I => \N__43455\
        );

    \I__9958\ : CEMux
    port map (
            O => \N__43461\,
            I => \N__43452\
        );

    \I__9957\ : LocalMux
    port map (
            O => \N__43458\,
            I => \N__43448\
        );

    \I__9956\ : LocalMux
    port map (
            O => \N__43455\,
            I => \N__43445\
        );

    \I__9955\ : LocalMux
    port map (
            O => \N__43452\,
            I => \N__43442\
        );

    \I__9954\ : CEMux
    port map (
            O => \N__43451\,
            I => \N__43439\
        );

    \I__9953\ : Span4Mux_v
    port map (
            O => \N__43448\,
            I => \N__43434\
        );

    \I__9952\ : Span4Mux_h
    port map (
            O => \N__43445\,
            I => \N__43434\
        );

    \I__9951\ : Span4Mux_v
    port map (
            O => \N__43442\,
            I => \N__43429\
        );

    \I__9950\ : LocalMux
    port map (
            O => \N__43439\,
            I => \N__43429\
        );

    \I__9949\ : Odrv4
    port map (
            O => \N__43434\,
            I => \delay_measurement_inst.N_265_i_0\
        );

    \I__9948\ : Odrv4
    port map (
            O => \N__43429\,
            I => \delay_measurement_inst.N_265_i_0\
        );

    \I__9947\ : InMux
    port map (
            O => \N__43424\,
            I => \N__43420\
        );

    \I__9946\ : InMux
    port map (
            O => \N__43423\,
            I => \N__43416\
        );

    \I__9945\ : LocalMux
    port map (
            O => \N__43420\,
            I => \N__43413\
        );

    \I__9944\ : InMux
    port map (
            O => \N__43419\,
            I => \N__43410\
        );

    \I__9943\ : LocalMux
    port map (
            O => \N__43416\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__9942\ : Odrv4
    port map (
            O => \N__43413\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__9941\ : LocalMux
    port map (
            O => \N__43410\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__9940\ : CascadeMux
    port map (
            O => \N__43403\,
            I => \N__43398\
        );

    \I__9939\ : CascadeMux
    port map (
            O => \N__43402\,
            I => \N__43395\
        );

    \I__9938\ : InMux
    port map (
            O => \N__43401\,
            I => \N__43392\
        );

    \I__9937\ : InMux
    port map (
            O => \N__43398\,
            I => \N__43389\
        );

    \I__9936\ : InMux
    port map (
            O => \N__43395\,
            I => \N__43386\
        );

    \I__9935\ : LocalMux
    port map (
            O => \N__43392\,
            I => \N__43383\
        );

    \I__9934\ : LocalMux
    port map (
            O => \N__43389\,
            I => \N__43380\
        );

    \I__9933\ : LocalMux
    port map (
            O => \N__43386\,
            I => \N__43377\
        );

    \I__9932\ : Span4Mux_v
    port map (
            O => \N__43383\,
            I => \N__43370\
        );

    \I__9931\ : Span4Mux_h
    port map (
            O => \N__43380\,
            I => \N__43370\
        );

    \I__9930\ : Span4Mux_v
    port map (
            O => \N__43377\,
            I => \N__43370\
        );

    \I__9929\ : Odrv4
    port map (
            O => \N__43370\,
            I => \delay_measurement_inst.elapsed_time_tr_3\
        );

    \I__9928\ : InMux
    port map (
            O => \N__43367\,
            I => \N__43363\
        );

    \I__9927\ : InMux
    port map (
            O => \N__43366\,
            I => \N__43359\
        );

    \I__9926\ : LocalMux
    port map (
            O => \N__43363\,
            I => \N__43356\
        );

    \I__9925\ : InMux
    port map (
            O => \N__43362\,
            I => \N__43353\
        );

    \I__9924\ : LocalMux
    port map (
            O => \N__43359\,
            I => \phase_controller_inst1.stoper_tr.time_passed11\
        );

    \I__9923\ : Odrv4
    port map (
            O => \N__43356\,
            I => \phase_controller_inst1.stoper_tr.time_passed11\
        );

    \I__9922\ : LocalMux
    port map (
            O => \N__43353\,
            I => \phase_controller_inst1.stoper_tr.time_passed11\
        );

    \I__9921\ : InMux
    port map (
            O => \N__43346\,
            I => \N__43338\
        );

    \I__9920\ : InMux
    port map (
            O => \N__43345\,
            I => \N__43338\
        );

    \I__9919\ : CascadeMux
    port map (
            O => \N__43344\,
            I => \N__43335\
        );

    \I__9918\ : InMux
    port map (
            O => \N__43343\,
            I => \N__43330\
        );

    \I__9917\ : LocalMux
    port map (
            O => \N__43338\,
            I => \N__43327\
        );

    \I__9916\ : InMux
    port map (
            O => \N__43335\,
            I => \N__43320\
        );

    \I__9915\ : InMux
    port map (
            O => \N__43334\,
            I => \N__43320\
        );

    \I__9914\ : InMux
    port map (
            O => \N__43333\,
            I => \N__43320\
        );

    \I__9913\ : LocalMux
    port map (
            O => \N__43330\,
            I => \N__43317\
        );

    \I__9912\ : Span4Mux_h
    port map (
            O => \N__43327\,
            I => \N__43314\
        );

    \I__9911\ : LocalMux
    port map (
            O => \N__43320\,
            I => \N__43311\
        );

    \I__9910\ : Odrv4
    port map (
            O => \N__43317\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__9909\ : Odrv4
    port map (
            O => \N__43314\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__9908\ : Odrv12
    port map (
            O => \N__43311\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__9907\ : CascadeMux
    port map (
            O => \N__43304\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\
        );

    \I__9906\ : CascadeMux
    port map (
            O => \N__43301\,
            I => \phase_controller_inst1.stoper_tr.time_passed11_cascade_\
        );

    \I__9905\ : InMux
    port map (
            O => \N__43298\,
            I => \N__43293\
        );

    \I__9904\ : InMux
    port map (
            O => \N__43297\,
            I => \N__43290\
        );

    \I__9903\ : CascadeMux
    port map (
            O => \N__43296\,
            I => \N__43286\
        );

    \I__9902\ : LocalMux
    port map (
            O => \N__43293\,
            I => \N__43283\
        );

    \I__9901\ : LocalMux
    port map (
            O => \N__43290\,
            I => \N__43280\
        );

    \I__9900\ : InMux
    port map (
            O => \N__43289\,
            I => \N__43275\
        );

    \I__9899\ : InMux
    port map (
            O => \N__43286\,
            I => \N__43275\
        );

    \I__9898\ : Span4Mux_h
    port map (
            O => \N__43283\,
            I => \N__43272\
        );

    \I__9897\ : Span4Mux_v
    port map (
            O => \N__43280\,
            I => \N__43267\
        );

    \I__9896\ : LocalMux
    port map (
            O => \N__43275\,
            I => \N__43267\
        );

    \I__9895\ : Span4Mux_v
    port map (
            O => \N__43272\,
            I => \N__43264\
        );

    \I__9894\ : Span4Mux_v
    port map (
            O => \N__43267\,
            I => \N__43261\
        );

    \I__9893\ : Odrv4
    port map (
            O => \N__43264\,
            I => measured_delay_tr_17
        );

    \I__9892\ : Odrv4
    port map (
            O => \N__43261\,
            I => measured_delay_tr_17
        );

    \I__9891\ : InMux
    port map (
            O => \N__43256\,
            I => \N__43246\
        );

    \I__9890\ : InMux
    port map (
            O => \N__43255\,
            I => \N__43246\
        );

    \I__9889\ : InMux
    port map (
            O => \N__43254\,
            I => \N__43246\
        );

    \I__9888\ : InMux
    port map (
            O => \N__43253\,
            I => \N__43243\
        );

    \I__9887\ : LocalMux
    port map (
            O => \N__43246\,
            I => \N__43236\
        );

    \I__9886\ : LocalMux
    port map (
            O => \N__43243\,
            I => \N__43233\
        );

    \I__9885\ : InMux
    port map (
            O => \N__43242\,
            I => \N__43230\
        );

    \I__9884\ : InMux
    port map (
            O => \N__43241\,
            I => \N__43225\
        );

    \I__9883\ : InMux
    port map (
            O => \N__43240\,
            I => \N__43225\
        );

    \I__9882\ : InMux
    port map (
            O => \N__43239\,
            I => \N__43222\
        );

    \I__9881\ : Odrv4
    port map (
            O => \N__43236\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20\
        );

    \I__9880\ : Odrv4
    port map (
            O => \N__43233\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20\
        );

    \I__9879\ : LocalMux
    port map (
            O => \N__43230\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20\
        );

    \I__9878\ : LocalMux
    port map (
            O => \N__43225\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20\
        );

    \I__9877\ : LocalMux
    port map (
            O => \N__43222\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20\
        );

    \I__9876\ : InMux
    port map (
            O => \N__43211\,
            I => \N__43207\
        );

    \I__9875\ : InMux
    port map (
            O => \N__43210\,
            I => \N__43202\
        );

    \I__9874\ : LocalMux
    port map (
            O => \N__43207\,
            I => \N__43199\
        );

    \I__9873\ : InMux
    port map (
            O => \N__43206\,
            I => \N__43194\
        );

    \I__9872\ : InMux
    port map (
            O => \N__43205\,
            I => \N__43194\
        );

    \I__9871\ : LocalMux
    port map (
            O => \N__43202\,
            I => \N__43191\
        );

    \I__9870\ : Span4Mux_v
    port map (
            O => \N__43199\,
            I => \N__43186\
        );

    \I__9869\ : LocalMux
    port map (
            O => \N__43194\,
            I => \N__43186\
        );

    \I__9868\ : Span4Mux_v
    port map (
            O => \N__43191\,
            I => \N__43183\
        );

    \I__9867\ : Span4Mux_v
    port map (
            O => \N__43186\,
            I => \N__43180\
        );

    \I__9866\ : Odrv4
    port map (
            O => \N__43183\,
            I => measured_delay_tr_18
        );

    \I__9865\ : Odrv4
    port map (
            O => \N__43180\,
            I => measured_delay_tr_18
        );

    \I__9864\ : InMux
    port map (
            O => \N__43175\,
            I => \N__43172\
        );

    \I__9863\ : LocalMux
    port map (
            O => \N__43172\,
            I => \N__43169\
        );

    \I__9862\ : Span4Mux_v
    port map (
            O => \N__43169\,
            I => \N__43166\
        );

    \I__9861\ : Span4Mux_h
    port map (
            O => \N__43166\,
            I => \N__43163\
        );

    \I__9860\ : Odrv4
    port map (
            O => \N__43163\,
            I => \phase_controller_inst1.N_83\
        );

    \I__9859\ : InMux
    port map (
            O => \N__43160\,
            I => \N__43157\
        );

    \I__9858\ : LocalMux
    port map (
            O => \N__43157\,
            I => \N__43154\
        );

    \I__9857\ : Span12Mux_h
    port map (
            O => \N__43154\,
            I => \N__43147\
        );

    \I__9856\ : InMux
    port map (
            O => \N__43153\,
            I => \N__43144\
        );

    \I__9855\ : InMux
    port map (
            O => \N__43152\,
            I => \N__43141\
        );

    \I__9854\ : InMux
    port map (
            O => \N__43151\,
            I => \N__43136\
        );

    \I__9853\ : InMux
    port map (
            O => \N__43150\,
            I => \N__43136\
        );

    \I__9852\ : Odrv12
    port map (
            O => \N__43147\,
            I => \phase_controller_inst1.stateZ0Z_4\
        );

    \I__9851\ : LocalMux
    port map (
            O => \N__43144\,
            I => \phase_controller_inst1.stateZ0Z_4\
        );

    \I__9850\ : LocalMux
    port map (
            O => \N__43141\,
            I => \phase_controller_inst1.stateZ0Z_4\
        );

    \I__9849\ : LocalMux
    port map (
            O => \N__43136\,
            I => \phase_controller_inst1.stateZ0Z_4\
        );

    \I__9848\ : CascadeMux
    port map (
            O => \N__43127\,
            I => \phase_controller_inst1.N_83_cascade_\
        );

    \I__9847\ : InMux
    port map (
            O => \N__43124\,
            I => \N__43121\
        );

    \I__9846\ : LocalMux
    port map (
            O => \N__43121\,
            I => \N__43118\
        );

    \I__9845\ : Span4Mux_v
    port map (
            O => \N__43118\,
            I => \N__43114\
        );

    \I__9844\ : InMux
    port map (
            O => \N__43117\,
            I => \N__43111\
        );

    \I__9843\ : Span4Mux_h
    port map (
            O => \N__43114\,
            I => \N__43106\
        );

    \I__9842\ : LocalMux
    port map (
            O => \N__43111\,
            I => \N__43106\
        );

    \I__9841\ : Odrv4
    port map (
            O => \N__43106\,
            I => \phase_controller_inst1.T01_0_sqmuxa\
        );

    \I__9840\ : CascadeMux
    port map (
            O => \N__43103\,
            I => \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa_cascade_\
        );

    \I__9839\ : InMux
    port map (
            O => \N__43100\,
            I => \N__43097\
        );

    \I__9838\ : LocalMux
    port map (
            O => \N__43097\,
            I => \N__43093\
        );

    \I__9837\ : InMux
    port map (
            O => \N__43096\,
            I => \N__43090\
        );

    \I__9836\ : Span4Mux_v
    port map (
            O => \N__43093\,
            I => \N__43087\
        );

    \I__9835\ : LocalMux
    port map (
            O => \N__43090\,
            I => \N__43084\
        );

    \I__9834\ : Span4Mux_v
    port map (
            O => \N__43087\,
            I => \N__43081\
        );

    \I__9833\ : Span4Mux_v
    port map (
            O => \N__43084\,
            I => \N__43078\
        );

    \I__9832\ : Span4Mux_v
    port map (
            O => \N__43081\,
            I => \N__43071\
        );

    \I__9831\ : Span4Mux_h
    port map (
            O => \N__43078\,
            I => \N__43071\
        );

    \I__9830\ : InMux
    port map (
            O => \N__43077\,
            I => \N__43068\
        );

    \I__9829\ : InMux
    port map (
            O => \N__43076\,
            I => \N__43065\
        );

    \I__9828\ : Span4Mux_v
    port map (
            O => \N__43071\,
            I => \N__43060\
        );

    \I__9827\ : LocalMux
    port map (
            O => \N__43068\,
            I => \N__43060\
        );

    \I__9826\ : LocalMux
    port map (
            O => \N__43065\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__9825\ : Odrv4
    port map (
            O => \N__43060\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__9824\ : CascadeMux
    port map (
            O => \N__43055\,
            I => \N__43051\
        );

    \I__9823\ : InMux
    port map (
            O => \N__43054\,
            I => \N__43043\
        );

    \I__9822\ : InMux
    port map (
            O => \N__43051\,
            I => \N__43043\
        );

    \I__9821\ : InMux
    port map (
            O => \N__43050\,
            I => \N__43043\
        );

    \I__9820\ : LocalMux
    port map (
            O => \N__43043\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__9819\ : InMux
    port map (
            O => \N__43040\,
            I => \N__43037\
        );

    \I__9818\ : LocalMux
    port map (
            O => \N__43037\,
            I => \N__43034\
        );

    \I__9817\ : Span4Mux_h
    port map (
            O => \N__43034\,
            I => \N__43030\
        );

    \I__9816\ : InMux
    port map (
            O => \N__43033\,
            I => \N__43027\
        );

    \I__9815\ : Span4Mux_h
    port map (
            O => \N__43030\,
            I => \N__43024\
        );

    \I__9814\ : LocalMux
    port map (
            O => \N__43027\,
            I => \N__43020\
        );

    \I__9813\ : Span4Mux_v
    port map (
            O => \N__43024\,
            I => \N__43017\
        );

    \I__9812\ : InMux
    port map (
            O => \N__43023\,
            I => \N__43014\
        );

    \I__9811\ : Span4Mux_h
    port map (
            O => \N__43020\,
            I => \N__43011\
        );

    \I__9810\ : Odrv4
    port map (
            O => \N__43017\,
            I => \il_min_comp1_D2\
        );

    \I__9809\ : LocalMux
    port map (
            O => \N__43014\,
            I => \il_min_comp1_D2\
        );

    \I__9808\ : Odrv4
    port map (
            O => \N__43011\,
            I => \il_min_comp1_D2\
        );

    \I__9807\ : InMux
    port map (
            O => \N__43004\,
            I => \N__42998\
        );

    \I__9806\ : InMux
    port map (
            O => \N__43003\,
            I => \N__42998\
        );

    \I__9805\ : LocalMux
    port map (
            O => \N__42998\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__9804\ : InMux
    port map (
            O => \N__42995\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_24\
        );

    \I__9803\ : InMux
    port map (
            O => \N__42992\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_25\
        );

    \I__9802\ : InMux
    port map (
            O => \N__42989\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_26\
        );

    \I__9801\ : InMux
    port map (
            O => \N__42986\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_27\
        );

    \I__9800\ : InMux
    port map (
            O => \N__42983\,
            I => \N__42971\
        );

    \I__9799\ : InMux
    port map (
            O => \N__42982\,
            I => \N__42971\
        );

    \I__9798\ : InMux
    port map (
            O => \N__42981\,
            I => \N__42971\
        );

    \I__9797\ : InMux
    port map (
            O => \N__42980\,
            I => \N__42971\
        );

    \I__9796\ : LocalMux
    port map (
            O => \N__42971\,
            I => \N__42942\
        );

    \I__9795\ : InMux
    port map (
            O => \N__42970\,
            I => \N__42937\
        );

    \I__9794\ : InMux
    port map (
            O => \N__42969\,
            I => \N__42937\
        );

    \I__9793\ : InMux
    port map (
            O => \N__42968\,
            I => \N__42928\
        );

    \I__9792\ : InMux
    port map (
            O => \N__42967\,
            I => \N__42928\
        );

    \I__9791\ : InMux
    port map (
            O => \N__42966\,
            I => \N__42928\
        );

    \I__9790\ : InMux
    port map (
            O => \N__42965\,
            I => \N__42928\
        );

    \I__9789\ : InMux
    port map (
            O => \N__42964\,
            I => \N__42919\
        );

    \I__9788\ : InMux
    port map (
            O => \N__42963\,
            I => \N__42919\
        );

    \I__9787\ : InMux
    port map (
            O => \N__42962\,
            I => \N__42919\
        );

    \I__9786\ : InMux
    port map (
            O => \N__42961\,
            I => \N__42919\
        );

    \I__9785\ : InMux
    port map (
            O => \N__42960\,
            I => \N__42910\
        );

    \I__9784\ : InMux
    port map (
            O => \N__42959\,
            I => \N__42910\
        );

    \I__9783\ : InMux
    port map (
            O => \N__42958\,
            I => \N__42910\
        );

    \I__9782\ : InMux
    port map (
            O => \N__42957\,
            I => \N__42910\
        );

    \I__9781\ : InMux
    port map (
            O => \N__42956\,
            I => \N__42901\
        );

    \I__9780\ : InMux
    port map (
            O => \N__42955\,
            I => \N__42901\
        );

    \I__9779\ : InMux
    port map (
            O => \N__42954\,
            I => \N__42901\
        );

    \I__9778\ : InMux
    port map (
            O => \N__42953\,
            I => \N__42901\
        );

    \I__9777\ : InMux
    port map (
            O => \N__42952\,
            I => \N__42892\
        );

    \I__9776\ : InMux
    port map (
            O => \N__42951\,
            I => \N__42892\
        );

    \I__9775\ : InMux
    port map (
            O => \N__42950\,
            I => \N__42892\
        );

    \I__9774\ : InMux
    port map (
            O => \N__42949\,
            I => \N__42892\
        );

    \I__9773\ : InMux
    port map (
            O => \N__42948\,
            I => \N__42883\
        );

    \I__9772\ : InMux
    port map (
            O => \N__42947\,
            I => \N__42883\
        );

    \I__9771\ : InMux
    port map (
            O => \N__42946\,
            I => \N__42883\
        );

    \I__9770\ : InMux
    port map (
            O => \N__42945\,
            I => \N__42883\
        );

    \I__9769\ : Span4Mux_h
    port map (
            O => \N__42942\,
            I => \N__42878\
        );

    \I__9768\ : LocalMux
    port map (
            O => \N__42937\,
            I => \N__42878\
        );

    \I__9767\ : LocalMux
    port map (
            O => \N__42928\,
            I => \N__42873\
        );

    \I__9766\ : LocalMux
    port map (
            O => \N__42919\,
            I => \N__42873\
        );

    \I__9765\ : LocalMux
    port map (
            O => \N__42910\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__9764\ : LocalMux
    port map (
            O => \N__42901\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__9763\ : LocalMux
    port map (
            O => \N__42892\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__9762\ : LocalMux
    port map (
            O => \N__42883\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__9761\ : Odrv4
    port map (
            O => \N__42878\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__9760\ : Odrv4
    port map (
            O => \N__42873\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__9759\ : InMux
    port map (
            O => \N__42860\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_28\
        );

    \I__9758\ : CEMux
    port map (
            O => \N__42857\,
            I => \N__42853\
        );

    \I__9757\ : CEMux
    port map (
            O => \N__42856\,
            I => \N__42850\
        );

    \I__9756\ : LocalMux
    port map (
            O => \N__42853\,
            I => \N__42846\
        );

    \I__9755\ : LocalMux
    port map (
            O => \N__42850\,
            I => \N__42843\
        );

    \I__9754\ : CEMux
    port map (
            O => \N__42849\,
            I => \N__42840\
        );

    \I__9753\ : Span4Mux_v
    port map (
            O => \N__42846\,
            I => \N__42832\
        );

    \I__9752\ : Span4Mux_v
    port map (
            O => \N__42843\,
            I => \N__42832\
        );

    \I__9751\ : LocalMux
    port map (
            O => \N__42840\,
            I => \N__42832\
        );

    \I__9750\ : CEMux
    port map (
            O => \N__42839\,
            I => \N__42829\
        );

    \I__9749\ : Span4Mux_v
    port map (
            O => \N__42832\,
            I => \N__42826\
        );

    \I__9748\ : LocalMux
    port map (
            O => \N__42829\,
            I => \N__42823\
        );

    \I__9747\ : Span4Mux_h
    port map (
            O => \N__42826\,
            I => \N__42818\
        );

    \I__9746\ : Span4Mux_v
    port map (
            O => \N__42823\,
            I => \N__42818\
        );

    \I__9745\ : Span4Mux_v
    port map (
            O => \N__42818\,
            I => \N__42815\
        );

    \I__9744\ : Odrv4
    port map (
            O => \N__42815\,
            I => \delay_measurement_inst.delay_tr_timer.N_324_i\
        );

    \I__9743\ : InMux
    port map (
            O => \N__42812\,
            I => \N__42809\
        );

    \I__9742\ : LocalMux
    port map (
            O => \N__42809\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_7_19\
        );

    \I__9741\ : InMux
    port map (
            O => \N__42806\,
            I => \N__42803\
        );

    \I__9740\ : LocalMux
    port map (
            O => \N__42803\,
            I => \N__42800\
        );

    \I__9739\ : Odrv4
    port map (
            O => \N__42800\,
            I => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_4\
        );

    \I__9738\ : InMux
    port map (
            O => \N__42797\,
            I => \N__42793\
        );

    \I__9737\ : InMux
    port map (
            O => \N__42796\,
            I => \N__42790\
        );

    \I__9736\ : LocalMux
    port map (
            O => \N__42793\,
            I => \N__42786\
        );

    \I__9735\ : LocalMux
    port map (
            O => \N__42790\,
            I => \N__42783\
        );

    \I__9734\ : InMux
    port map (
            O => \N__42789\,
            I => \N__42780\
        );

    \I__9733\ : Span4Mux_v
    port map (
            O => \N__42786\,
            I => \N__42775\
        );

    \I__9732\ : Span4Mux_v
    port map (
            O => \N__42783\,
            I => \N__42775\
        );

    \I__9731\ : LocalMux
    port map (
            O => \N__42780\,
            I => \delay_measurement_inst.elapsed_time_tr_2\
        );

    \I__9730\ : Odrv4
    port map (
            O => \N__42775\,
            I => \delay_measurement_inst.elapsed_time_tr_2\
        );

    \I__9729\ : InMux
    port map (
            O => \N__42770\,
            I => \N__42765\
        );

    \I__9728\ : CascadeMux
    port map (
            O => \N__42769\,
            I => \N__42761\
        );

    \I__9727\ : InMux
    port map (
            O => \N__42768\,
            I => \N__42758\
        );

    \I__9726\ : LocalMux
    port map (
            O => \N__42765\,
            I => \N__42755\
        );

    \I__9725\ : InMux
    port map (
            O => \N__42764\,
            I => \N__42752\
        );

    \I__9724\ : InMux
    port map (
            O => \N__42761\,
            I => \N__42749\
        );

    \I__9723\ : LocalMux
    port map (
            O => \N__42758\,
            I => \N__42744\
        );

    \I__9722\ : Span4Mux_h
    port map (
            O => \N__42755\,
            I => \N__42744\
        );

    \I__9721\ : LocalMux
    port map (
            O => \N__42752\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16\
        );

    \I__9720\ : LocalMux
    port map (
            O => \N__42749\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16\
        );

    \I__9719\ : Odrv4
    port map (
            O => \N__42744\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16\
        );

    \I__9718\ : InMux
    port map (
            O => \N__42737\,
            I => \bfn_17_13_0_\
        );

    \I__9717\ : InMux
    port map (
            O => \N__42734\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_16\
        );

    \I__9716\ : InMux
    port map (
            O => \N__42731\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_17\
        );

    \I__9715\ : InMux
    port map (
            O => \N__42728\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_18\
        );

    \I__9714\ : InMux
    port map (
            O => \N__42725\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_19\
        );

    \I__9713\ : InMux
    port map (
            O => \N__42722\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_20\
        );

    \I__9712\ : InMux
    port map (
            O => \N__42719\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_21\
        );

    \I__9711\ : InMux
    port map (
            O => \N__42716\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_22\
        );

    \I__9710\ : InMux
    port map (
            O => \N__42713\,
            I => \bfn_17_14_0_\
        );

    \I__9709\ : InMux
    port map (
            O => \N__42710\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_6\
        );

    \I__9708\ : InMux
    port map (
            O => \N__42707\,
            I => \bfn_17_12_0_\
        );

    \I__9707\ : InMux
    port map (
            O => \N__42704\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_8\
        );

    \I__9706\ : InMux
    port map (
            O => \N__42701\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_9\
        );

    \I__9705\ : InMux
    port map (
            O => \N__42698\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_10\
        );

    \I__9704\ : InMux
    port map (
            O => \N__42695\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_11\
        );

    \I__9703\ : InMux
    port map (
            O => \N__42692\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_12\
        );

    \I__9702\ : InMux
    port map (
            O => \N__42689\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_13\
        );

    \I__9701\ : InMux
    port map (
            O => \N__42686\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_14\
        );

    \I__9700\ : CascadeMux
    port map (
            O => \N__42683\,
            I => \N__42679\
        );

    \I__9699\ : CascadeMux
    port map (
            O => \N__42682\,
            I => \N__42676\
        );

    \I__9698\ : InMux
    port map (
            O => \N__42679\,
            I => \N__42671\
        );

    \I__9697\ : InMux
    port map (
            O => \N__42676\,
            I => \N__42671\
        );

    \I__9696\ : LocalMux
    port map (
            O => \N__42671\,
            I => \N__42668\
        );

    \I__9695\ : Span4Mux_v
    port map (
            O => \N__42668\,
            I => \N__42664\
        );

    \I__9694\ : InMux
    port map (
            O => \N__42667\,
            I => \N__42661\
        );

    \I__9693\ : Span4Mux_h
    port map (
            O => \N__42664\,
            I => \N__42658\
        );

    \I__9692\ : LocalMux
    port map (
            O => \N__42661\,
            I => measured_delay_hc_22
        );

    \I__9691\ : Odrv4
    port map (
            O => \N__42658\,
            I => measured_delay_hc_22
        );

    \I__9690\ : CascadeMux
    port map (
            O => \N__42653\,
            I => \N__42641\
        );

    \I__9689\ : CascadeMux
    port map (
            O => \N__42652\,
            I => \N__42637\
        );

    \I__9688\ : CascadeMux
    port map (
            O => \N__42651\,
            I => \N__42633\
        );

    \I__9687\ : InMux
    port map (
            O => \N__42650\,
            I => \N__42615\
        );

    \I__9686\ : InMux
    port map (
            O => \N__42649\,
            I => \N__42615\
        );

    \I__9685\ : InMux
    port map (
            O => \N__42648\,
            I => \N__42612\
        );

    \I__9684\ : InMux
    port map (
            O => \N__42647\,
            I => \N__42605\
        );

    \I__9683\ : InMux
    port map (
            O => \N__42646\,
            I => \N__42605\
        );

    \I__9682\ : InMux
    port map (
            O => \N__42645\,
            I => \N__42605\
        );

    \I__9681\ : InMux
    port map (
            O => \N__42644\,
            I => \N__42594\
        );

    \I__9680\ : InMux
    port map (
            O => \N__42641\,
            I => \N__42594\
        );

    \I__9679\ : InMux
    port map (
            O => \N__42640\,
            I => \N__42594\
        );

    \I__9678\ : InMux
    port map (
            O => \N__42637\,
            I => \N__42594\
        );

    \I__9677\ : InMux
    port map (
            O => \N__42636\,
            I => \N__42594\
        );

    \I__9676\ : InMux
    port map (
            O => \N__42633\,
            I => \N__42583\
        );

    \I__9675\ : InMux
    port map (
            O => \N__42632\,
            I => \N__42583\
        );

    \I__9674\ : InMux
    port map (
            O => \N__42631\,
            I => \N__42583\
        );

    \I__9673\ : InMux
    port map (
            O => \N__42630\,
            I => \N__42583\
        );

    \I__9672\ : InMux
    port map (
            O => \N__42629\,
            I => \N__42583\
        );

    \I__9671\ : InMux
    port map (
            O => \N__42628\,
            I => \N__42574\
        );

    \I__9670\ : InMux
    port map (
            O => \N__42627\,
            I => \N__42574\
        );

    \I__9669\ : InMux
    port map (
            O => \N__42626\,
            I => \N__42574\
        );

    \I__9668\ : InMux
    port map (
            O => \N__42625\,
            I => \N__42574\
        );

    \I__9667\ : InMux
    port map (
            O => \N__42624\,
            I => \N__42571\
        );

    \I__9666\ : InMux
    port map (
            O => \N__42623\,
            I => \N__42564\
        );

    \I__9665\ : InMux
    port map (
            O => \N__42622\,
            I => \N__42564\
        );

    \I__9664\ : InMux
    port map (
            O => \N__42621\,
            I => \N__42564\
        );

    \I__9663\ : InMux
    port map (
            O => \N__42620\,
            I => \N__42561\
        );

    \I__9662\ : LocalMux
    port map (
            O => \N__42615\,
            I => \N__42555\
        );

    \I__9661\ : LocalMux
    port map (
            O => \N__42612\,
            I => \N__42552\
        );

    \I__9660\ : LocalMux
    port map (
            O => \N__42605\,
            I => \N__42544\
        );

    \I__9659\ : LocalMux
    port map (
            O => \N__42594\,
            I => \N__42544\
        );

    \I__9658\ : LocalMux
    port map (
            O => \N__42583\,
            I => \N__42544\
        );

    \I__9657\ : LocalMux
    port map (
            O => \N__42574\,
            I => \N__42535\
        );

    \I__9656\ : LocalMux
    port map (
            O => \N__42571\,
            I => \N__42535\
        );

    \I__9655\ : LocalMux
    port map (
            O => \N__42564\,
            I => \N__42535\
        );

    \I__9654\ : LocalMux
    port map (
            O => \N__42561\,
            I => \N__42535\
        );

    \I__9653\ : InMux
    port map (
            O => \N__42560\,
            I => \N__42528\
        );

    \I__9652\ : InMux
    port map (
            O => \N__42559\,
            I => \N__42528\
        );

    \I__9651\ : InMux
    port map (
            O => \N__42558\,
            I => \N__42528\
        );

    \I__9650\ : Span4Mux_v
    port map (
            O => \N__42555\,
            I => \N__42522\
        );

    \I__9649\ : Span4Mux_h
    port map (
            O => \N__42552\,
            I => \N__42519\
        );

    \I__9648\ : InMux
    port map (
            O => \N__42551\,
            I => \N__42516\
        );

    \I__9647\ : Span4Mux_v
    port map (
            O => \N__42544\,
            I => \N__42509\
        );

    \I__9646\ : Span4Mux_v
    port map (
            O => \N__42535\,
            I => \N__42509\
        );

    \I__9645\ : LocalMux
    port map (
            O => \N__42528\,
            I => \N__42509\
        );

    \I__9644\ : InMux
    port map (
            O => \N__42527\,
            I => \N__42502\
        );

    \I__9643\ : InMux
    port map (
            O => \N__42526\,
            I => \N__42502\
        );

    \I__9642\ : InMux
    port map (
            O => \N__42525\,
            I => \N__42502\
        );

    \I__9641\ : Odrv4
    port map (
            O => \N__42522\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__9640\ : Odrv4
    port map (
            O => \N__42519\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__9639\ : LocalMux
    port map (
            O => \N__42516\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__9638\ : Odrv4
    port map (
            O => \N__42509\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__9637\ : LocalMux
    port map (
            O => \N__42502\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__9636\ : CascadeMux
    port map (
            O => \N__42491\,
            I => \N__42488\
        );

    \I__9635\ : InMux
    port map (
            O => \N__42488\,
            I => \N__42485\
        );

    \I__9634\ : LocalMux
    port map (
            O => \N__42485\,
            I => \N__42482\
        );

    \I__9633\ : Span4Mux_h
    port map (
            O => \N__42482\,
            I => \N__42477\
        );

    \I__9632\ : InMux
    port map (
            O => \N__42481\,
            I => \N__42472\
        );

    \I__9631\ : InMux
    port map (
            O => \N__42480\,
            I => \N__42472\
        );

    \I__9630\ : Odrv4
    port map (
            O => \N__42477\,
            I => \delay_measurement_inst.elapsed_time_hc_17\
        );

    \I__9629\ : LocalMux
    port map (
            O => \N__42472\,
            I => \delay_measurement_inst.elapsed_time_hc_17\
        );

    \I__9628\ : InMux
    port map (
            O => \N__42467\,
            I => \N__42454\
        );

    \I__9627\ : InMux
    port map (
            O => \N__42466\,
            I => \N__42454\
        );

    \I__9626\ : InMux
    port map (
            O => \N__42465\,
            I => \N__42454\
        );

    \I__9625\ : InMux
    port map (
            O => \N__42464\,
            I => \N__42447\
        );

    \I__9624\ : InMux
    port map (
            O => \N__42463\,
            I => \N__42447\
        );

    \I__9623\ : InMux
    port map (
            O => \N__42462\,
            I => \N__42447\
        );

    \I__9622\ : InMux
    port map (
            O => \N__42461\,
            I => \N__42435\
        );

    \I__9621\ : LocalMux
    port map (
            O => \N__42454\,
            I => \N__42432\
        );

    \I__9620\ : LocalMux
    port map (
            O => \N__42447\,
            I => \N__42429\
        );

    \I__9619\ : InMux
    port map (
            O => \N__42446\,
            I => \N__42422\
        );

    \I__9618\ : InMux
    port map (
            O => \N__42445\,
            I => \N__42422\
        );

    \I__9617\ : InMux
    port map (
            O => \N__42444\,
            I => \N__42422\
        );

    \I__9616\ : InMux
    port map (
            O => \N__42443\,
            I => \N__42412\
        );

    \I__9615\ : InMux
    port map (
            O => \N__42442\,
            I => \N__42412\
        );

    \I__9614\ : InMux
    port map (
            O => \N__42441\,
            I => \N__42403\
        );

    \I__9613\ : InMux
    port map (
            O => \N__42440\,
            I => \N__42403\
        );

    \I__9612\ : InMux
    port map (
            O => \N__42439\,
            I => \N__42403\
        );

    \I__9611\ : InMux
    port map (
            O => \N__42438\,
            I => \N__42403\
        );

    \I__9610\ : LocalMux
    port map (
            O => \N__42435\,
            I => \N__42400\
        );

    \I__9609\ : Span4Mux_v
    port map (
            O => \N__42432\,
            I => \N__42393\
        );

    \I__9608\ : Span4Mux_v
    port map (
            O => \N__42429\,
            I => \N__42393\
        );

    \I__9607\ : LocalMux
    port map (
            O => \N__42422\,
            I => \N__42393\
        );

    \I__9606\ : InMux
    port map (
            O => \N__42421\,
            I => \N__42384\
        );

    \I__9605\ : InMux
    port map (
            O => \N__42420\,
            I => \N__42384\
        );

    \I__9604\ : InMux
    port map (
            O => \N__42419\,
            I => \N__42384\
        );

    \I__9603\ : InMux
    port map (
            O => \N__42418\,
            I => \N__42384\
        );

    \I__9602\ : InMux
    port map (
            O => \N__42417\,
            I => \N__42381\
        );

    \I__9601\ : LocalMux
    port map (
            O => \N__42412\,
            I => \N__42375\
        );

    \I__9600\ : LocalMux
    port map (
            O => \N__42403\,
            I => \N__42372\
        );

    \I__9599\ : Span4Mux_v
    port map (
            O => \N__42400\,
            I => \N__42363\
        );

    \I__9598\ : Span4Mux_h
    port map (
            O => \N__42393\,
            I => \N__42363\
        );

    \I__9597\ : LocalMux
    port map (
            O => \N__42384\,
            I => \N__42363\
        );

    \I__9596\ : LocalMux
    port map (
            O => \N__42381\,
            I => \N__42363\
        );

    \I__9595\ : InMux
    port map (
            O => \N__42380\,
            I => \N__42356\
        );

    \I__9594\ : InMux
    port map (
            O => \N__42379\,
            I => \N__42356\
        );

    \I__9593\ : InMux
    port map (
            O => \N__42378\,
            I => \N__42356\
        );

    \I__9592\ : Odrv4
    port map (
            O => \N__42375\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__9591\ : Odrv12
    port map (
            O => \N__42372\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__9590\ : Odrv4
    port map (
            O => \N__42363\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__9589\ : LocalMux
    port map (
            O => \N__42356\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__9588\ : InMux
    port map (
            O => \N__42347\,
            I => \N__42343\
        );

    \I__9587\ : InMux
    port map (
            O => \N__42346\,
            I => \N__42340\
        );

    \I__9586\ : LocalMux
    port map (
            O => \N__42343\,
            I => \N__42336\
        );

    \I__9585\ : LocalMux
    port map (
            O => \N__42340\,
            I => \N__42333\
        );

    \I__9584\ : InMux
    port map (
            O => \N__42339\,
            I => \N__42330\
        );

    \I__9583\ : Span4Mux_v
    port map (
            O => \N__42336\,
            I => \N__42326\
        );

    \I__9582\ : Span4Mux_h
    port map (
            O => \N__42333\,
            I => \N__42323\
        );

    \I__9581\ : LocalMux
    port map (
            O => \N__42330\,
            I => \N__42320\
        );

    \I__9580\ : InMux
    port map (
            O => \N__42329\,
            I => \N__42316\
        );

    \I__9579\ : Span4Mux_v
    port map (
            O => \N__42326\,
            I => \N__42311\
        );

    \I__9578\ : Span4Mux_h
    port map (
            O => \N__42323\,
            I => \N__42311\
        );

    \I__9577\ : Span4Mux_v
    port map (
            O => \N__42320\,
            I => \N__42308\
        );

    \I__9576\ : InMux
    port map (
            O => \N__42319\,
            I => \N__42305\
        );

    \I__9575\ : LocalMux
    port map (
            O => \N__42316\,
            I => measured_delay_hc_17
        );

    \I__9574\ : Odrv4
    port map (
            O => \N__42311\,
            I => measured_delay_hc_17
        );

    \I__9573\ : Odrv4
    port map (
            O => \N__42308\,
            I => measured_delay_hc_17
        );

    \I__9572\ : LocalMux
    port map (
            O => \N__42305\,
            I => measured_delay_hc_17
        );

    \I__9571\ : InMux
    port map (
            O => \N__42296\,
            I => \bfn_17_11_0_\
        );

    \I__9570\ : InMux
    port map (
            O => \N__42293\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_0\
        );

    \I__9569\ : InMux
    port map (
            O => \N__42290\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_1\
        );

    \I__9568\ : InMux
    port map (
            O => \N__42287\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_2\
        );

    \I__9567\ : InMux
    port map (
            O => \N__42284\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_3\
        );

    \I__9566\ : InMux
    port map (
            O => \N__42281\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_4\
        );

    \I__9565\ : InMux
    port map (
            O => \N__42278\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_5\
        );

    \I__9564\ : CascadeMux
    port map (
            O => \N__42275\,
            I => \N__42271\
        );

    \I__9563\ : InMux
    port map (
            O => \N__42274\,
            I => \N__42268\
        );

    \I__9562\ : InMux
    port map (
            O => \N__42271\,
            I => \N__42265\
        );

    \I__9561\ : LocalMux
    port map (
            O => \N__42268\,
            I => measured_delay_hc_24
        );

    \I__9560\ : LocalMux
    port map (
            O => \N__42265\,
            I => measured_delay_hc_24
        );

    \I__9559\ : CascadeMux
    port map (
            O => \N__42260\,
            I => \N__42256\
        );

    \I__9558\ : CascadeMux
    port map (
            O => \N__42259\,
            I => \N__42253\
        );

    \I__9557\ : InMux
    port map (
            O => \N__42256\,
            I => \N__42250\
        );

    \I__9556\ : InMux
    port map (
            O => \N__42253\,
            I => \N__42247\
        );

    \I__9555\ : LocalMux
    port map (
            O => \N__42250\,
            I => \N__42244\
        );

    \I__9554\ : LocalMux
    port map (
            O => \N__42247\,
            I => \N__42240\
        );

    \I__9553\ : Span4Mux_v
    port map (
            O => \N__42244\,
            I => \N__42237\
        );

    \I__9552\ : InMux
    port map (
            O => \N__42243\,
            I => \N__42234\
        );

    \I__9551\ : Span4Mux_v
    port map (
            O => \N__42240\,
            I => \N__42230\
        );

    \I__9550\ : Span4Mux_h
    port map (
            O => \N__42237\,
            I => \N__42225\
        );

    \I__9549\ : LocalMux
    port map (
            O => \N__42234\,
            I => \N__42225\
        );

    \I__9548\ : InMux
    port map (
            O => \N__42233\,
            I => \N__42222\
        );

    \I__9547\ : Span4Mux_v
    port map (
            O => \N__42230\,
            I => \N__42219\
        );

    \I__9546\ : Span4Mux_h
    port map (
            O => \N__42225\,
            I => \N__42216\
        );

    \I__9545\ : LocalMux
    port map (
            O => \N__42222\,
            I => measured_delay_hc_0
        );

    \I__9544\ : Odrv4
    port map (
            O => \N__42219\,
            I => measured_delay_hc_0
        );

    \I__9543\ : Odrv4
    port map (
            O => \N__42216\,
            I => measured_delay_hc_0
        );

    \I__9542\ : InMux
    port map (
            O => \N__42209\,
            I => \N__42206\
        );

    \I__9541\ : LocalMux
    port map (
            O => \N__42206\,
            I => \N__42201\
        );

    \I__9540\ : InMux
    port map (
            O => \N__42205\,
            I => \N__42196\
        );

    \I__9539\ : InMux
    port map (
            O => \N__42204\,
            I => \N__42196\
        );

    \I__9538\ : Odrv4
    port map (
            O => \N__42201\,
            I => \delay_measurement_inst.elapsed_time_hc_18\
        );

    \I__9537\ : LocalMux
    port map (
            O => \N__42196\,
            I => \delay_measurement_inst.elapsed_time_hc_18\
        );

    \I__9536\ : InMux
    port map (
            O => \N__42191\,
            I => \N__42187\
        );

    \I__9535\ : InMux
    port map (
            O => \N__42190\,
            I => \N__42184\
        );

    \I__9534\ : LocalMux
    port map (
            O => \N__42187\,
            I => \N__42178\
        );

    \I__9533\ : LocalMux
    port map (
            O => \N__42184\,
            I => \N__42175\
        );

    \I__9532\ : InMux
    port map (
            O => \N__42183\,
            I => \N__42172\
        );

    \I__9531\ : CascadeMux
    port map (
            O => \N__42182\,
            I => \N__42169\
        );

    \I__9530\ : CascadeMux
    port map (
            O => \N__42181\,
            I => \N__42166\
        );

    \I__9529\ : Span4Mux_v
    port map (
            O => \N__42178\,
            I => \N__42163\
        );

    \I__9528\ : Span4Mux_v
    port map (
            O => \N__42175\,
            I => \N__42160\
        );

    \I__9527\ : LocalMux
    port map (
            O => \N__42172\,
            I => \N__42157\
        );

    \I__9526\ : InMux
    port map (
            O => \N__42169\,
            I => \N__42154\
        );

    \I__9525\ : InMux
    port map (
            O => \N__42166\,
            I => \N__42151\
        );

    \I__9524\ : Span4Mux_h
    port map (
            O => \N__42163\,
            I => \N__42148\
        );

    \I__9523\ : Span4Mux_v
    port map (
            O => \N__42160\,
            I => \N__42141\
        );

    \I__9522\ : Span4Mux_h
    port map (
            O => \N__42157\,
            I => \N__42141\
        );

    \I__9521\ : LocalMux
    port map (
            O => \N__42154\,
            I => \N__42141\
        );

    \I__9520\ : LocalMux
    port map (
            O => \N__42151\,
            I => measured_delay_hc_18
        );

    \I__9519\ : Odrv4
    port map (
            O => \N__42148\,
            I => measured_delay_hc_18
        );

    \I__9518\ : Odrv4
    port map (
            O => \N__42141\,
            I => measured_delay_hc_18
        );

    \I__9517\ : CascadeMux
    port map (
            O => \N__42134\,
            I => \N__42131\
        );

    \I__9516\ : InMux
    port map (
            O => \N__42131\,
            I => \N__42126\
        );

    \I__9515\ : InMux
    port map (
            O => \N__42130\,
            I => \N__42123\
        );

    \I__9514\ : CascadeMux
    port map (
            O => \N__42129\,
            I => \N__42120\
        );

    \I__9513\ : LocalMux
    port map (
            O => \N__42126\,
            I => \N__42117\
        );

    \I__9512\ : LocalMux
    port map (
            O => \N__42123\,
            I => \N__42114\
        );

    \I__9511\ : InMux
    port map (
            O => \N__42120\,
            I => \N__42111\
        );

    \I__9510\ : Odrv4
    port map (
            O => \N__42117\,
            I => \delay_measurement_inst.elapsed_time_hc_19\
        );

    \I__9509\ : Odrv4
    port map (
            O => \N__42114\,
            I => \delay_measurement_inst.elapsed_time_hc_19\
        );

    \I__9508\ : LocalMux
    port map (
            O => \N__42111\,
            I => \delay_measurement_inst.elapsed_time_hc_19\
        );

    \I__9507\ : InMux
    port map (
            O => \N__42104\,
            I => \N__42094\
        );

    \I__9506\ : InMux
    port map (
            O => \N__42103\,
            I => \N__42094\
        );

    \I__9505\ : InMux
    port map (
            O => \N__42102\,
            I => \N__42089\
        );

    \I__9504\ : InMux
    port map (
            O => \N__42101\,
            I => \N__42082\
        );

    \I__9503\ : InMux
    port map (
            O => \N__42100\,
            I => \N__42082\
        );

    \I__9502\ : InMux
    port map (
            O => \N__42099\,
            I => \N__42082\
        );

    \I__9501\ : LocalMux
    port map (
            O => \N__42094\,
            I => \N__42079\
        );

    \I__9500\ : InMux
    port map (
            O => \N__42093\,
            I => \N__42076\
        );

    \I__9499\ : InMux
    port map (
            O => \N__42092\,
            I => \N__42073\
        );

    \I__9498\ : LocalMux
    port map (
            O => \N__42089\,
            I => \N__42070\
        );

    \I__9497\ : LocalMux
    port map (
            O => \N__42082\,
            I => \N__42067\
        );

    \I__9496\ : Span4Mux_v
    port map (
            O => \N__42079\,
            I => \N__42062\
        );

    \I__9495\ : LocalMux
    port map (
            O => \N__42076\,
            I => \N__42062\
        );

    \I__9494\ : LocalMux
    port map (
            O => \N__42073\,
            I => \delay_measurement_inst.delay_hc_reg3lto31_0_0\
        );

    \I__9493\ : Odrv4
    port map (
            O => \N__42070\,
            I => \delay_measurement_inst.delay_hc_reg3lto31_0_0\
        );

    \I__9492\ : Odrv4
    port map (
            O => \N__42067\,
            I => \delay_measurement_inst.delay_hc_reg3lto31_0_0\
        );

    \I__9491\ : Odrv4
    port map (
            O => \N__42062\,
            I => \delay_measurement_inst.delay_hc_reg3lto31_0_0\
        );

    \I__9490\ : CascadeMux
    port map (
            O => \N__42053\,
            I => \N__42050\
        );

    \I__9489\ : InMux
    port map (
            O => \N__42050\,
            I => \N__42045\
        );

    \I__9488\ : InMux
    port map (
            O => \N__42049\,
            I => \N__42042\
        );

    \I__9487\ : InMux
    port map (
            O => \N__42048\,
            I => \N__42039\
        );

    \I__9486\ : LocalMux
    port map (
            O => \N__42045\,
            I => \N__42036\
        );

    \I__9485\ : LocalMux
    port map (
            O => \N__42042\,
            I => \N__42033\
        );

    \I__9484\ : LocalMux
    port map (
            O => \N__42039\,
            I => \N__42028\
        );

    \I__9483\ : Span4Mux_v
    port map (
            O => \N__42036\,
            I => \N__42028\
        );

    \I__9482\ : Span4Mux_v
    port map (
            O => \N__42033\,
            I => \N__42025\
        );

    \I__9481\ : Odrv4
    port map (
            O => \N__42028\,
            I => measured_delay_hc_19
        );

    \I__9480\ : Odrv4
    port map (
            O => \N__42025\,
            I => measured_delay_hc_19
        );

    \I__9479\ : InMux
    port map (
            O => \N__42020\,
            I => \N__42014\
        );

    \I__9478\ : InMux
    port map (
            O => \N__42019\,
            I => \N__42014\
        );

    \I__9477\ : LocalMux
    port map (
            O => \N__42014\,
            I => \N__42010\
        );

    \I__9476\ : InMux
    port map (
            O => \N__42013\,
            I => \N__42007\
        );

    \I__9475\ : Span4Mux_h
    port map (
            O => \N__42010\,
            I => \N__42004\
        );

    \I__9474\ : LocalMux
    port map (
            O => \N__42007\,
            I => measured_delay_hc_21
        );

    \I__9473\ : Odrv4
    port map (
            O => \N__42004\,
            I => measured_delay_hc_21
        );

    \I__9472\ : InMux
    port map (
            O => \N__41999\,
            I => \N__41995\
        );

    \I__9471\ : InMux
    port map (
            O => \N__41998\,
            I => \N__41992\
        );

    \I__9470\ : LocalMux
    port map (
            O => \N__41995\,
            I => \N__41988\
        );

    \I__9469\ : LocalMux
    port map (
            O => \N__41992\,
            I => \N__41985\
        );

    \I__9468\ : CascadeMux
    port map (
            O => \N__41991\,
            I => \N__41982\
        );

    \I__9467\ : Span4Mux_v
    port map (
            O => \N__41988\,
            I => \N__41979\
        );

    \I__9466\ : Span4Mux_v
    port map (
            O => \N__41985\,
            I => \N__41976\
        );

    \I__9465\ : InMux
    port map (
            O => \N__41982\,
            I => \N__41973\
        );

    \I__9464\ : Odrv4
    port map (
            O => \N__41979\,
            I => measured_delay_tr_13
        );

    \I__9463\ : Odrv4
    port map (
            O => \N__41976\,
            I => measured_delay_tr_13
        );

    \I__9462\ : LocalMux
    port map (
            O => \N__41973\,
            I => measured_delay_tr_13
        );

    \I__9461\ : CascadeMux
    port map (
            O => \N__41966\,
            I => \N__41963\
        );

    \I__9460\ : InMux
    port map (
            O => \N__41963\,
            I => \N__41960\
        );

    \I__9459\ : LocalMux
    port map (
            O => \N__41960\,
            I => \N__41957\
        );

    \I__9458\ : Odrv12
    port map (
            O => \N__41957\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\
        );

    \I__9457\ : InMux
    port map (
            O => \N__41954\,
            I => \N__41951\
        );

    \I__9456\ : LocalMux
    port map (
            O => \N__41951\,
            I => \N__41948\
        );

    \I__9455\ : Odrv12
    port map (
            O => \N__41948\,
            I => delay_hc_input_c
        );

    \I__9454\ : InMux
    port map (
            O => \N__41945\,
            I => \N__41942\
        );

    \I__9453\ : LocalMux
    port map (
            O => \N__41942\,
            I => delay_hc_d1
        );

    \I__9452\ : InMux
    port map (
            O => \N__41939\,
            I => \N__41936\
        );

    \I__9451\ : LocalMux
    port map (
            O => \N__41936\,
            I => \N__41933\
        );

    \I__9450\ : Span4Mux_v
    port map (
            O => \N__41933\,
            I => \N__41927\
        );

    \I__9449\ : InMux
    port map (
            O => \N__41932\,
            I => \N__41922\
        );

    \I__9448\ : InMux
    port map (
            O => \N__41931\,
            I => \N__41922\
        );

    \I__9447\ : InMux
    port map (
            O => \N__41930\,
            I => \N__41919\
        );

    \I__9446\ : Span4Mux_h
    port map (
            O => \N__41927\,
            I => \N__41916\
        );

    \I__9445\ : LocalMux
    port map (
            O => \N__41922\,
            I => \N__41913\
        );

    \I__9444\ : LocalMux
    port map (
            O => \N__41919\,
            I => \N__41910\
        );

    \I__9443\ : Span4Mux_v
    port map (
            O => \N__41916\,
            I => \N__41907\
        );

    \I__9442\ : Span12Mux_v
    port map (
            O => \N__41913\,
            I => \N__41904\
        );

    \I__9441\ : Span4Mux_v
    port map (
            O => \N__41910\,
            I => \N__41901\
        );

    \I__9440\ : Odrv4
    port map (
            O => \N__41907\,
            I => delay_hc_d2
        );

    \I__9439\ : Odrv12
    port map (
            O => \N__41904\,
            I => delay_hc_d2
        );

    \I__9438\ : Odrv4
    port map (
            O => \N__41901\,
            I => delay_hc_d2
        );

    \I__9437\ : InMux
    port map (
            O => \N__41894\,
            I => \N__41891\
        );

    \I__9436\ : LocalMux
    port map (
            O => \N__41891\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_3\
        );

    \I__9435\ : InMux
    port map (
            O => \N__41888\,
            I => \N__41883\
        );

    \I__9434\ : InMux
    port map (
            O => \N__41887\,
            I => \N__41880\
        );

    \I__9433\ : InMux
    port map (
            O => \N__41886\,
            I => \N__41877\
        );

    \I__9432\ : LocalMux
    port map (
            O => \N__41883\,
            I => \N__41873\
        );

    \I__9431\ : LocalMux
    port map (
            O => \N__41880\,
            I => \N__41870\
        );

    \I__9430\ : LocalMux
    port map (
            O => \N__41877\,
            I => \N__41867\
        );

    \I__9429\ : InMux
    port map (
            O => \N__41876\,
            I => \N__41864\
        );

    \I__9428\ : Span4Mux_v
    port map (
            O => \N__41873\,
            I => \N__41861\
        );

    \I__9427\ : Sp12to4
    port map (
            O => \N__41870\,
            I => \N__41856\
        );

    \I__9426\ : Sp12to4
    port map (
            O => \N__41867\,
            I => \N__41856\
        );

    \I__9425\ : LocalMux
    port map (
            O => \N__41864\,
            I => \N__41853\
        );

    \I__9424\ : Sp12to4
    port map (
            O => \N__41861\,
            I => \N__41850\
        );

    \I__9423\ : Span12Mux_v
    port map (
            O => \N__41856\,
            I => \N__41847\
        );

    \I__9422\ : Span4Mux_v
    port map (
            O => \N__41853\,
            I => \N__41844\
        );

    \I__9421\ : Odrv12
    port map (
            O => \N__41850\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_2\
        );

    \I__9420\ : Odrv12
    port map (
            O => \N__41847\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_2\
        );

    \I__9419\ : Odrv4
    port map (
            O => \N__41844\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_2\
        );

    \I__9418\ : InMux
    port map (
            O => \N__41837\,
            I => \N__41833\
        );

    \I__9417\ : InMux
    port map (
            O => \N__41836\,
            I => \N__41830\
        );

    \I__9416\ : LocalMux
    port map (
            O => \N__41833\,
            I => measured_delay_hc_25
        );

    \I__9415\ : LocalMux
    port map (
            O => \N__41830\,
            I => measured_delay_hc_25
        );

    \I__9414\ : InMux
    port map (
            O => \N__41825\,
            I => \N__41821\
        );

    \I__9413\ : InMux
    port map (
            O => \N__41824\,
            I => \N__41818\
        );

    \I__9412\ : LocalMux
    port map (
            O => \N__41821\,
            I => measured_delay_hc_26
        );

    \I__9411\ : LocalMux
    port map (
            O => \N__41818\,
            I => measured_delay_hc_26
        );

    \I__9410\ : CascadeMux
    port map (
            O => \N__41813\,
            I => \N__41810\
        );

    \I__9409\ : InMux
    port map (
            O => \N__41810\,
            I => \N__41804\
        );

    \I__9408\ : InMux
    port map (
            O => \N__41809\,
            I => \N__41804\
        );

    \I__9407\ : LocalMux
    port map (
            O => \N__41804\,
            I => measured_delay_hc_23
        );

    \I__9406\ : InMux
    port map (
            O => \N__41801\,
            I => \N__41798\
        );

    \I__9405\ : LocalMux
    port map (
            O => \N__41798\,
            I => \N__41794\
        );

    \I__9404\ : CascadeMux
    port map (
            O => \N__41797\,
            I => \N__41789\
        );

    \I__9403\ : Span4Mux_v
    port map (
            O => \N__41794\,
            I => \N__41786\
        );

    \I__9402\ : InMux
    port map (
            O => \N__41793\,
            I => \N__41783\
        );

    \I__9401\ : InMux
    port map (
            O => \N__41792\,
            I => \N__41780\
        );

    \I__9400\ : InMux
    port map (
            O => \N__41789\,
            I => \N__41777\
        );

    \I__9399\ : Odrv4
    port map (
            O => \N__41786\,
            I => \delay_measurement_inst.elapsed_time_hc_8\
        );

    \I__9398\ : LocalMux
    port map (
            O => \N__41783\,
            I => \delay_measurement_inst.elapsed_time_hc_8\
        );

    \I__9397\ : LocalMux
    port map (
            O => \N__41780\,
            I => \delay_measurement_inst.elapsed_time_hc_8\
        );

    \I__9396\ : LocalMux
    port map (
            O => \N__41777\,
            I => \delay_measurement_inst.elapsed_time_hc_8\
        );

    \I__9395\ : InMux
    port map (
            O => \N__41768\,
            I => \N__41764\
        );

    \I__9394\ : InMux
    port map (
            O => \N__41767\,
            I => \N__41760\
        );

    \I__9393\ : LocalMux
    port map (
            O => \N__41764\,
            I => \N__41757\
        );

    \I__9392\ : CascadeMux
    port map (
            O => \N__41763\,
            I => \N__41753\
        );

    \I__9391\ : LocalMux
    port map (
            O => \N__41760\,
            I => \N__41750\
        );

    \I__9390\ : Span4Mux_v
    port map (
            O => \N__41757\,
            I => \N__41747\
        );

    \I__9389\ : InMux
    port map (
            O => \N__41756\,
            I => \N__41744\
        );

    \I__9388\ : InMux
    port map (
            O => \N__41753\,
            I => \N__41741\
        );

    \I__9387\ : Span4Mux_v
    port map (
            O => \N__41750\,
            I => \N__41737\
        );

    \I__9386\ : Span4Mux_h
    port map (
            O => \N__41747\,
            I => \N__41734\
        );

    \I__9385\ : LocalMux
    port map (
            O => \N__41744\,
            I => \N__41731\
        );

    \I__9384\ : LocalMux
    port map (
            O => \N__41741\,
            I => \N__41728\
        );

    \I__9383\ : InMux
    port map (
            O => \N__41740\,
            I => \N__41725\
        );

    \I__9382\ : Span4Mux_v
    port map (
            O => \N__41737\,
            I => \N__41722\
        );

    \I__9381\ : Span4Mux_h
    port map (
            O => \N__41734\,
            I => \N__41715\
        );

    \I__9380\ : Span4Mux_v
    port map (
            O => \N__41731\,
            I => \N__41715\
        );

    \I__9379\ : Span4Mux_v
    port map (
            O => \N__41728\,
            I => \N__41715\
        );

    \I__9378\ : LocalMux
    port map (
            O => \N__41725\,
            I => measured_delay_hc_8
        );

    \I__9377\ : Odrv4
    port map (
            O => \N__41722\,
            I => measured_delay_hc_8
        );

    \I__9376\ : Odrv4
    port map (
            O => \N__41715\,
            I => measured_delay_hc_8
        );

    \I__9375\ : CascadeMux
    port map (
            O => \N__41708\,
            I => \N__41705\
        );

    \I__9374\ : InMux
    port map (
            O => \N__41705\,
            I => \N__41702\
        );

    \I__9373\ : LocalMux
    port map (
            O => \N__41702\,
            I => \N__41699\
        );

    \I__9372\ : Span4Mux_v
    port map (
            O => \N__41699\,
            I => \N__41693\
        );

    \I__9371\ : InMux
    port map (
            O => \N__41698\,
            I => \N__41690\
        );

    \I__9370\ : InMux
    port map (
            O => \N__41697\,
            I => \N__41687\
        );

    \I__9369\ : InMux
    port map (
            O => \N__41696\,
            I => \N__41684\
        );

    \I__9368\ : Odrv4
    port map (
            O => \N__41693\,
            I => \delay_measurement_inst.elapsed_time_hc_7\
        );

    \I__9367\ : LocalMux
    port map (
            O => \N__41690\,
            I => \delay_measurement_inst.elapsed_time_hc_7\
        );

    \I__9366\ : LocalMux
    port map (
            O => \N__41687\,
            I => \delay_measurement_inst.elapsed_time_hc_7\
        );

    \I__9365\ : LocalMux
    port map (
            O => \N__41684\,
            I => \delay_measurement_inst.elapsed_time_hc_7\
        );

    \I__9364\ : InMux
    port map (
            O => \N__41675\,
            I => \N__41672\
        );

    \I__9363\ : LocalMux
    port map (
            O => \N__41672\,
            I => \N__41667\
        );

    \I__9362\ : InMux
    port map (
            O => \N__41671\,
            I => \N__41664\
        );

    \I__9361\ : InMux
    port map (
            O => \N__41670\,
            I => \N__41661\
        );

    \I__9360\ : Span4Mux_v
    port map (
            O => \N__41667\,
            I => \N__41655\
        );

    \I__9359\ : LocalMux
    port map (
            O => \N__41664\,
            I => \N__41655\
        );

    \I__9358\ : LocalMux
    port map (
            O => \N__41661\,
            I => \N__41652\
        );

    \I__9357\ : InMux
    port map (
            O => \N__41660\,
            I => \N__41649\
        );

    \I__9356\ : Span4Mux_v
    port map (
            O => \N__41655\,
            I => \N__41645\
        );

    \I__9355\ : Span4Mux_h
    port map (
            O => \N__41652\,
            I => \N__41640\
        );

    \I__9354\ : LocalMux
    port map (
            O => \N__41649\,
            I => \N__41640\
        );

    \I__9353\ : InMux
    port map (
            O => \N__41648\,
            I => \N__41637\
        );

    \I__9352\ : Span4Mux_h
    port map (
            O => \N__41645\,
            I => \N__41634\
        );

    \I__9351\ : Span4Mux_h
    port map (
            O => \N__41640\,
            I => \N__41631\
        );

    \I__9350\ : LocalMux
    port map (
            O => \N__41637\,
            I => measured_delay_hc_7
        );

    \I__9349\ : Odrv4
    port map (
            O => \N__41634\,
            I => measured_delay_hc_7
        );

    \I__9348\ : Odrv4
    port map (
            O => \N__41631\,
            I => measured_delay_hc_7
        );

    \I__9347\ : InMux
    port map (
            O => \N__41624\,
            I => \N__41621\
        );

    \I__9346\ : LocalMux
    port map (
            O => \N__41621\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_16\
        );

    \I__9345\ : CascadeMux
    port map (
            O => \N__41618\,
            I => \N__41615\
        );

    \I__9344\ : InMux
    port map (
            O => \N__41615\,
            I => \N__41612\
        );

    \I__9343\ : LocalMux
    port map (
            O => \N__41612\,
            I => \N__41609\
        );

    \I__9342\ : Odrv4
    port map (
            O => \N__41609\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\
        );

    \I__9341\ : InMux
    port map (
            O => \N__41606\,
            I => \N__41603\
        );

    \I__9340\ : LocalMux
    port map (
            O => \N__41603\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_17\
        );

    \I__9339\ : InMux
    port map (
            O => \N__41600\,
            I => \N__41597\
        );

    \I__9338\ : LocalMux
    port map (
            O => \N__41597\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_18\
        );

    \I__9337\ : InMux
    port map (
            O => \N__41594\,
            I => \N__41591\
        );

    \I__9336\ : LocalMux
    port map (
            O => \N__41591\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_19\
        );

    \I__9335\ : InMux
    port map (
            O => \N__41588\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__9334\ : CascadeMux
    port map (
            O => \N__41585\,
            I => \N__41582\
        );

    \I__9333\ : InMux
    port map (
            O => \N__41582\,
            I => \N__41579\
        );

    \I__9332\ : LocalMux
    port map (
            O => \N__41579\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\
        );

    \I__9331\ : InMux
    port map (
            O => \N__41576\,
            I => \N__41572\
        );

    \I__9330\ : CascadeMux
    port map (
            O => \N__41575\,
            I => \N__41569\
        );

    \I__9329\ : LocalMux
    port map (
            O => \N__41572\,
            I => \N__41564\
        );

    \I__9328\ : InMux
    port map (
            O => \N__41569\,
            I => \N__41559\
        );

    \I__9327\ : InMux
    port map (
            O => \N__41568\,
            I => \N__41559\
        );

    \I__9326\ : InMux
    port map (
            O => \N__41567\,
            I => \N__41556\
        );

    \I__9325\ : Span4Mux_v
    port map (
            O => \N__41564\,
            I => \N__41551\
        );

    \I__9324\ : LocalMux
    port map (
            O => \N__41559\,
            I => \N__41551\
        );

    \I__9323\ : LocalMux
    port map (
            O => \N__41556\,
            I => \N__41548\
        );

    \I__9322\ : Span4Mux_v
    port map (
            O => \N__41551\,
            I => \N__41545\
        );

    \I__9321\ : Odrv12
    port map (
            O => \N__41548\,
            I => measured_delay_tr_19
        );

    \I__9320\ : Odrv4
    port map (
            O => \N__41545\,
            I => measured_delay_tr_19
        );

    \I__9319\ : CascadeMux
    port map (
            O => \N__41540\,
            I => \N__41537\
        );

    \I__9318\ : InMux
    port map (
            O => \N__41537\,
            I => \N__41534\
        );

    \I__9317\ : LocalMux
    port map (
            O => \N__41534\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\
        );

    \I__9316\ : InMux
    port map (
            O => \N__41531\,
            I => \N__41528\
        );

    \I__9315\ : LocalMux
    port map (
            O => \N__41528\,
            I => \N__41524\
        );

    \I__9314\ : InMux
    port map (
            O => \N__41527\,
            I => \N__41521\
        );

    \I__9313\ : Span4Mux_h
    port map (
            O => \N__41524\,
            I => \N__41517\
        );

    \I__9312\ : LocalMux
    port map (
            O => \N__41521\,
            I => \N__41514\
        );

    \I__9311\ : InMux
    port map (
            O => \N__41520\,
            I => \N__41511\
        );

    \I__9310\ : Odrv4
    port map (
            O => \N__41517\,
            I => measured_delay_tr_11
        );

    \I__9309\ : Odrv12
    port map (
            O => \N__41514\,
            I => measured_delay_tr_11
        );

    \I__9308\ : LocalMux
    port map (
            O => \N__41511\,
            I => measured_delay_tr_11
        );

    \I__9307\ : CascadeMux
    port map (
            O => \N__41504\,
            I => \N__41501\
        );

    \I__9306\ : InMux
    port map (
            O => \N__41501\,
            I => \N__41498\
        );

    \I__9305\ : LocalMux
    port map (
            O => \N__41498\,
            I => \N__41495\
        );

    \I__9304\ : Odrv4
    port map (
            O => \N__41495\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\
        );

    \I__9303\ : CascadeMux
    port map (
            O => \N__41492\,
            I => \N__41486\
        );

    \I__9302\ : InMux
    port map (
            O => \N__41491\,
            I => \N__41476\
        );

    \I__9301\ : InMux
    port map (
            O => \N__41490\,
            I => \N__41473\
        );

    \I__9300\ : InMux
    port map (
            O => \N__41489\,
            I => \N__41470\
        );

    \I__9299\ : InMux
    port map (
            O => \N__41486\,
            I => \N__41457\
        );

    \I__9298\ : InMux
    port map (
            O => \N__41485\,
            I => \N__41457\
        );

    \I__9297\ : InMux
    port map (
            O => \N__41484\,
            I => \N__41457\
        );

    \I__9296\ : InMux
    port map (
            O => \N__41483\,
            I => \N__41457\
        );

    \I__9295\ : InMux
    port map (
            O => \N__41482\,
            I => \N__41457\
        );

    \I__9294\ : InMux
    port map (
            O => \N__41481\,
            I => \N__41457\
        );

    \I__9293\ : CascadeMux
    port map (
            O => \N__41480\,
            I => \N__41454\
        );

    \I__9292\ : CascadeMux
    port map (
            O => \N__41479\,
            I => \N__41448\
        );

    \I__9291\ : LocalMux
    port map (
            O => \N__41476\,
            I => \N__41444\
        );

    \I__9290\ : LocalMux
    port map (
            O => \N__41473\,
            I => \N__41441\
        );

    \I__9289\ : LocalMux
    port map (
            O => \N__41470\,
            I => \N__41438\
        );

    \I__9288\ : LocalMux
    port map (
            O => \N__41457\,
            I => \N__41434\
        );

    \I__9287\ : InMux
    port map (
            O => \N__41454\,
            I => \N__41425\
        );

    \I__9286\ : InMux
    port map (
            O => \N__41453\,
            I => \N__41425\
        );

    \I__9285\ : InMux
    port map (
            O => \N__41452\,
            I => \N__41425\
        );

    \I__9284\ : InMux
    port map (
            O => \N__41451\,
            I => \N__41425\
        );

    \I__9283\ : InMux
    port map (
            O => \N__41448\,
            I => \N__41420\
        );

    \I__9282\ : InMux
    port map (
            O => \N__41447\,
            I => \N__41420\
        );

    \I__9281\ : Span4Mux_v
    port map (
            O => \N__41444\,
            I => \N__41415\
        );

    \I__9280\ : Span4Mux_v
    port map (
            O => \N__41441\,
            I => \N__41415\
        );

    \I__9279\ : Span12Mux_h
    port map (
            O => \N__41438\,
            I => \N__41412\
        );

    \I__9278\ : InMux
    port map (
            O => \N__41437\,
            I => \N__41409\
        );

    \I__9277\ : Span4Mux_h
    port map (
            O => \N__41434\,
            I => \N__41406\
        );

    \I__9276\ : LocalMux
    port map (
            O => \N__41425\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15\
        );

    \I__9275\ : LocalMux
    port map (
            O => \N__41420\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15\
        );

    \I__9274\ : Odrv4
    port map (
            O => \N__41415\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15\
        );

    \I__9273\ : Odrv12
    port map (
            O => \N__41412\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15\
        );

    \I__9272\ : LocalMux
    port map (
            O => \N__41409\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15\
        );

    \I__9271\ : Odrv4
    port map (
            O => \N__41406\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15\
        );

    \I__9270\ : CascadeMux
    port map (
            O => \N__41393\,
            I => \N__41390\
        );

    \I__9269\ : InMux
    port map (
            O => \N__41390\,
            I => \N__41387\
        );

    \I__9268\ : LocalMux
    port map (
            O => \N__41387\,
            I => \N__41384\
        );

    \I__9267\ : Odrv4
    port map (
            O => \N__41384\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\
        );

    \I__9266\ : CascadeMux
    port map (
            O => \N__41381\,
            I => \N__41378\
        );

    \I__9265\ : InMux
    port map (
            O => \N__41378\,
            I => \N__41375\
        );

    \I__9264\ : LocalMux
    port map (
            O => \N__41375\,
            I => \N__41372\
        );

    \I__9263\ : Odrv4
    port map (
            O => \N__41372\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\
        );

    \I__9262\ : InMux
    port map (
            O => \N__41369\,
            I => \N__41366\
        );

    \I__9261\ : LocalMux
    port map (
            O => \N__41366\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\
        );

    \I__9260\ : InMux
    port map (
            O => \N__41363\,
            I => \N__41360\
        );

    \I__9259\ : LocalMux
    port map (
            O => \N__41360\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\
        );

    \I__9258\ : CascadeMux
    port map (
            O => \N__41357\,
            I => \N__41354\
        );

    \I__9257\ : InMux
    port map (
            O => \N__41354\,
            I => \N__41351\
        );

    \I__9256\ : LocalMux
    port map (
            O => \N__41351\,
            I => \N__41348\
        );

    \I__9255\ : Span4Mux_h
    port map (
            O => \N__41348\,
            I => \N__41345\
        );

    \I__9254\ : Span4Mux_v
    port map (
            O => \N__41345\,
            I => \N__41342\
        );

    \I__9253\ : Odrv4
    port map (
            O => \N__41342\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\
        );

    \I__9252\ : InMux
    port map (
            O => \N__41339\,
            I => \N__41336\
        );

    \I__9251\ : LocalMux
    port map (
            O => \N__41336\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\
        );

    \I__9250\ : InMux
    port map (
            O => \N__41333\,
            I => \N__41330\
        );

    \I__9249\ : LocalMux
    port map (
            O => \N__41330\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\
        );

    \I__9248\ : CascadeMux
    port map (
            O => \N__41327\,
            I => \N__41324\
        );

    \I__9247\ : InMux
    port map (
            O => \N__41324\,
            I => \N__41321\
        );

    \I__9246\ : LocalMux
    port map (
            O => \N__41321\,
            I => \N__41318\
        );

    \I__9245\ : Span4Mux_h
    port map (
            O => \N__41318\,
            I => \N__41315\
        );

    \I__9244\ : Span4Mux_v
    port map (
            O => \N__41315\,
            I => \N__41312\
        );

    \I__9243\ : Odrv4
    port map (
            O => \N__41312\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\
        );

    \I__9242\ : InMux
    port map (
            O => \N__41309\,
            I => \N__41306\
        );

    \I__9241\ : LocalMux
    port map (
            O => \N__41306\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\
        );

    \I__9240\ : InMux
    port map (
            O => \N__41303\,
            I => \N__41300\
        );

    \I__9239\ : LocalMux
    port map (
            O => \N__41300\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\
        );

    \I__9238\ : CascadeMux
    port map (
            O => \N__41297\,
            I => \N__41294\
        );

    \I__9237\ : InMux
    port map (
            O => \N__41294\,
            I => \N__41291\
        );

    \I__9236\ : LocalMux
    port map (
            O => \N__41291\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\
        );

    \I__9235\ : InMux
    port map (
            O => \N__41288\,
            I => \N__41285\
        );

    \I__9234\ : LocalMux
    port map (
            O => \N__41285\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\
        );

    \I__9233\ : InMux
    port map (
            O => \N__41282\,
            I => \N__41279\
        );

    \I__9232\ : LocalMux
    port map (
            O => \N__41279\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\
        );

    \I__9231\ : CascadeMux
    port map (
            O => \N__41276\,
            I => \N__41272\
        );

    \I__9230\ : CascadeMux
    port map (
            O => \N__41275\,
            I => \N__41269\
        );

    \I__9229\ : InMux
    port map (
            O => \N__41272\,
            I => \N__41266\
        );

    \I__9228\ : InMux
    port map (
            O => \N__41269\,
            I => \N__41263\
        );

    \I__9227\ : LocalMux
    port map (
            O => \N__41266\,
            I => \N__41260\
        );

    \I__9226\ : LocalMux
    port map (
            O => \N__41263\,
            I => \N__41257\
        );

    \I__9225\ : Span4Mux_v
    port map (
            O => \N__41260\,
            I => \N__41254\
        );

    \I__9224\ : Span4Mux_h
    port map (
            O => \N__41257\,
            I => \N__41249\
        );

    \I__9223\ : Span4Mux_h
    port map (
            O => \N__41254\,
            I => \N__41245\
        );

    \I__9222\ : InMux
    port map (
            O => \N__41253\,
            I => \N__41242\
        );

    \I__9221\ : CascadeMux
    port map (
            O => \N__41252\,
            I => \N__41239\
        );

    \I__9220\ : Span4Mux_v
    port map (
            O => \N__41249\,
            I => \N__41236\
        );

    \I__9219\ : InMux
    port map (
            O => \N__41248\,
            I => \N__41233\
        );

    \I__9218\ : Span4Mux_h
    port map (
            O => \N__41245\,
            I => \N__41228\
        );

    \I__9217\ : LocalMux
    port map (
            O => \N__41242\,
            I => \N__41228\
        );

    \I__9216\ : InMux
    port map (
            O => \N__41239\,
            I => \N__41225\
        );

    \I__9215\ : Span4Mux_v
    port map (
            O => \N__41236\,
            I => \N__41220\
        );

    \I__9214\ : LocalMux
    port map (
            O => \N__41233\,
            I => \N__41220\
        );

    \I__9213\ : Span4Mux_v
    port map (
            O => \N__41228\,
            I => \N__41217\
        );

    \I__9212\ : LocalMux
    port map (
            O => \N__41225\,
            I => measured_delay_hc_1
        );

    \I__9211\ : Odrv4
    port map (
            O => \N__41220\,
            I => measured_delay_hc_1
        );

    \I__9210\ : Odrv4
    port map (
            O => \N__41217\,
            I => measured_delay_hc_1
        );

    \I__9209\ : CascadeMux
    port map (
            O => \N__41210\,
            I => \N__41207\
        );

    \I__9208\ : InMux
    port map (
            O => \N__41207\,
            I => \N__41204\
        );

    \I__9207\ : LocalMux
    port map (
            O => \N__41204\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_1\
        );

    \I__9206\ : CascadeMux
    port map (
            O => \N__41201\,
            I => \N__41198\
        );

    \I__9205\ : InMux
    port map (
            O => \N__41198\,
            I => \N__41195\
        );

    \I__9204\ : LocalMux
    port map (
            O => \N__41195\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\
        );

    \I__9203\ : InMux
    port map (
            O => \N__41192\,
            I => \N__41189\
        );

    \I__9202\ : LocalMux
    port map (
            O => \N__41189\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\
        );

    \I__9201\ : InMux
    port map (
            O => \N__41186\,
            I => \N__41183\
        );

    \I__9200\ : LocalMux
    port map (
            O => \N__41183\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\
        );

    \I__9199\ : CascadeMux
    port map (
            O => \N__41180\,
            I => \N__41177\
        );

    \I__9198\ : InMux
    port map (
            O => \N__41177\,
            I => \N__41174\
        );

    \I__9197\ : LocalMux
    port map (
            O => \N__41174\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\
        );

    \I__9196\ : CascadeMux
    port map (
            O => \N__41171\,
            I => \N__41168\
        );

    \I__9195\ : InMux
    port map (
            O => \N__41168\,
            I => \N__41165\
        );

    \I__9194\ : LocalMux
    port map (
            O => \N__41165\,
            I => \N__41162\
        );

    \I__9193\ : Span4Mux_h
    port map (
            O => \N__41162\,
            I => \N__41159\
        );

    \I__9192\ : Odrv4
    port map (
            O => \N__41159\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\
        );

    \I__9191\ : InMux
    port map (
            O => \N__41156\,
            I => \N__41153\
        );

    \I__9190\ : LocalMux
    port map (
            O => \N__41153\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\
        );

    \I__9189\ : CascadeMux
    port map (
            O => \N__41150\,
            I => \N__41147\
        );

    \I__9188\ : InMux
    port map (
            O => \N__41147\,
            I => \N__41144\
        );

    \I__9187\ : LocalMux
    port map (
            O => \N__41144\,
            I => \N__41141\
        );

    \I__9186\ : Odrv4
    port map (
            O => \N__41141\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\
        );

    \I__9185\ : InMux
    port map (
            O => \N__41138\,
            I => \N__41135\
        );

    \I__9184\ : LocalMux
    port map (
            O => \N__41135\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\
        );

    \I__9183\ : CascadeMux
    port map (
            O => \N__41132\,
            I => \N__41129\
        );

    \I__9182\ : InMux
    port map (
            O => \N__41129\,
            I => \N__41126\
        );

    \I__9181\ : LocalMux
    port map (
            O => \N__41126\,
            I => \N__41123\
        );

    \I__9180\ : Span4Mux_h
    port map (
            O => \N__41123\,
            I => \N__41120\
        );

    \I__9179\ : Odrv4
    port map (
            O => \N__41120\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\
        );

    \I__9178\ : InMux
    port map (
            O => \N__41117\,
            I => \N__41114\
        );

    \I__9177\ : LocalMux
    port map (
            O => \N__41114\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\
        );

    \I__9176\ : CascadeMux
    port map (
            O => \N__41111\,
            I => \N__41108\
        );

    \I__9175\ : InMux
    port map (
            O => \N__41108\,
            I => \N__41105\
        );

    \I__9174\ : LocalMux
    port map (
            O => \N__41105\,
            I => \N__41102\
        );

    \I__9173\ : Span4Mux_h
    port map (
            O => \N__41102\,
            I => \N__41099\
        );

    \I__9172\ : Odrv4
    port map (
            O => \N__41099\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\
        );

    \I__9171\ : InMux
    port map (
            O => \N__41096\,
            I => \N__41093\
        );

    \I__9170\ : LocalMux
    port map (
            O => \N__41093\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\
        );

    \I__9169\ : CascadeMux
    port map (
            O => \N__41090\,
            I => \N__41087\
        );

    \I__9168\ : InMux
    port map (
            O => \N__41087\,
            I => \N__41084\
        );

    \I__9167\ : LocalMux
    port map (
            O => \N__41084\,
            I => \N__41081\
        );

    \I__9166\ : Span4Mux_v
    port map (
            O => \N__41081\,
            I => \N__41078\
        );

    \I__9165\ : Odrv4
    port map (
            O => \N__41078\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\
        );

    \I__9164\ : InMux
    port map (
            O => \N__41075\,
            I => \N__41072\
        );

    \I__9163\ : LocalMux
    port map (
            O => \N__41072\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\
        );

    \I__9162\ : CascadeMux
    port map (
            O => \N__41069\,
            I => \N__41055\
        );

    \I__9161\ : InMux
    port map (
            O => \N__41068\,
            I => \N__41046\
        );

    \I__9160\ : InMux
    port map (
            O => \N__41067\,
            I => \N__41046\
        );

    \I__9159\ : InMux
    port map (
            O => \N__41066\,
            I => \N__41046\
        );

    \I__9158\ : InMux
    port map (
            O => \N__41065\,
            I => \N__41037\
        );

    \I__9157\ : InMux
    port map (
            O => \N__41064\,
            I => \N__41037\
        );

    \I__9156\ : InMux
    port map (
            O => \N__41063\,
            I => \N__41037\
        );

    \I__9155\ : InMux
    port map (
            O => \N__41062\,
            I => \N__41037\
        );

    \I__9154\ : InMux
    port map (
            O => \N__41061\,
            I => \N__41030\
        );

    \I__9153\ : InMux
    port map (
            O => \N__41060\,
            I => \N__41030\
        );

    \I__9152\ : InMux
    port map (
            O => \N__41059\,
            I => \N__41030\
        );

    \I__9151\ : InMux
    port map (
            O => \N__41058\,
            I => \N__41023\
        );

    \I__9150\ : InMux
    port map (
            O => \N__41055\,
            I => \N__41018\
        );

    \I__9149\ : InMux
    port map (
            O => \N__41054\,
            I => \N__41015\
        );

    \I__9148\ : InMux
    port map (
            O => \N__41053\,
            I => \N__41012\
        );

    \I__9147\ : LocalMux
    port map (
            O => \N__41046\,
            I => \N__41009\
        );

    \I__9146\ : LocalMux
    port map (
            O => \N__41037\,
            I => \N__41004\
        );

    \I__9145\ : LocalMux
    port map (
            O => \N__41030\,
            I => \N__41004\
        );

    \I__9144\ : CascadeMux
    port map (
            O => \N__41029\,
            I => \N__41001\
        );

    \I__9143\ : InMux
    port map (
            O => \N__41028\,
            I => \N__40991\
        );

    \I__9142\ : InMux
    port map (
            O => \N__41027\,
            I => \N__40991\
        );

    \I__9141\ : InMux
    port map (
            O => \N__41026\,
            I => \N__40991\
        );

    \I__9140\ : LocalMux
    port map (
            O => \N__41023\,
            I => \N__40988\
        );

    \I__9139\ : InMux
    port map (
            O => \N__41022\,
            I => \N__40985\
        );

    \I__9138\ : InMux
    port map (
            O => \N__41021\,
            I => \N__40982\
        );

    \I__9137\ : LocalMux
    port map (
            O => \N__41018\,
            I => \N__40970\
        );

    \I__9136\ : LocalMux
    port map (
            O => \N__41015\,
            I => \N__40970\
        );

    \I__9135\ : LocalMux
    port map (
            O => \N__41012\,
            I => \N__40970\
        );

    \I__9134\ : Span4Mux_v
    port map (
            O => \N__41009\,
            I => \N__40970\
        );

    \I__9133\ : Span4Mux_v
    port map (
            O => \N__41004\,
            I => \N__40970\
        );

    \I__9132\ : InMux
    port map (
            O => \N__41001\,
            I => \N__40961\
        );

    \I__9131\ : InMux
    port map (
            O => \N__41000\,
            I => \N__40961\
        );

    \I__9130\ : InMux
    port map (
            O => \N__40999\,
            I => \N__40961\
        );

    \I__9129\ : InMux
    port map (
            O => \N__40998\,
            I => \N__40961\
        );

    \I__9128\ : LocalMux
    port map (
            O => \N__40991\,
            I => \N__40956\
        );

    \I__9127\ : Span4Mux_v
    port map (
            O => \N__40988\,
            I => \N__40956\
        );

    \I__9126\ : LocalMux
    port map (
            O => \N__40985\,
            I => \N__40953\
        );

    \I__9125\ : LocalMux
    port map (
            O => \N__40982\,
            I => \N__40950\
        );

    \I__9124\ : InMux
    port map (
            O => \N__40981\,
            I => \N__40947\
        );

    \I__9123\ : Span4Mux_v
    port map (
            O => \N__40970\,
            I => \N__40942\
        );

    \I__9122\ : LocalMux
    port map (
            O => \N__40961\,
            I => \N__40942\
        );

    \I__9121\ : Span4Mux_v
    port map (
            O => \N__40956\,
            I => \N__40937\
        );

    \I__9120\ : Span4Mux_h
    port map (
            O => \N__40953\,
            I => \N__40937\
        );

    \I__9119\ : Span4Mux_v
    port map (
            O => \N__40950\,
            I => \N__40934\
        );

    \I__9118\ : LocalMux
    port map (
            O => \N__40947\,
            I => \N__40929\
        );

    \I__9117\ : Span4Mux_v
    port map (
            O => \N__40942\,
            I => \N__40929\
        );

    \I__9116\ : Span4Mux_v
    port map (
            O => \N__40937\,
            I => \N__40926\
        );

    \I__9115\ : Odrv4
    port map (
            O => \N__40934\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__9114\ : Odrv4
    port map (
            O => \N__40929\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__9113\ : Odrv4
    port map (
            O => \N__40926\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__9112\ : CascadeMux
    port map (
            O => \N__40919\,
            I => \N__40911\
        );

    \I__9111\ : CascadeMux
    port map (
            O => \N__40918\,
            I => \N__40906\
        );

    \I__9110\ : CascadeMux
    port map (
            O => \N__40917\,
            I => \N__40903\
        );

    \I__9109\ : CascadeMux
    port map (
            O => \N__40916\,
            I => \N__40896\
        );

    \I__9108\ : CascadeMux
    port map (
            O => \N__40915\,
            I => \N__40891\
        );

    \I__9107\ : CascadeMux
    port map (
            O => \N__40914\,
            I => \N__40888\
        );

    \I__9106\ : InMux
    port map (
            O => \N__40911\,
            I => \N__40885\
        );

    \I__9105\ : CascadeMux
    port map (
            O => \N__40910\,
            I => \N__40882\
        );

    \I__9104\ : CascadeMux
    port map (
            O => \N__40909\,
            I => \N__40879\
        );

    \I__9103\ : InMux
    port map (
            O => \N__40906\,
            I => \N__40876\
        );

    \I__9102\ : InMux
    port map (
            O => \N__40903\,
            I => \N__40873\
        );

    \I__9101\ : CascadeMux
    port map (
            O => \N__40902\,
            I => \N__40869\
        );

    \I__9100\ : CascadeMux
    port map (
            O => \N__40901\,
            I => \N__40866\
        );

    \I__9099\ : CascadeMux
    port map (
            O => \N__40900\,
            I => \N__40863\
        );

    \I__9098\ : CascadeMux
    port map (
            O => \N__40899\,
            I => \N__40854\
        );

    \I__9097\ : InMux
    port map (
            O => \N__40896\,
            I => \N__40849\
        );

    \I__9096\ : InMux
    port map (
            O => \N__40895\,
            I => \N__40842\
        );

    \I__9095\ : InMux
    port map (
            O => \N__40894\,
            I => \N__40842\
        );

    \I__9094\ : InMux
    port map (
            O => \N__40891\,
            I => \N__40842\
        );

    \I__9093\ : InMux
    port map (
            O => \N__40888\,
            I => \N__40839\
        );

    \I__9092\ : LocalMux
    port map (
            O => \N__40885\,
            I => \N__40836\
        );

    \I__9091\ : InMux
    port map (
            O => \N__40882\,
            I => \N__40831\
        );

    \I__9090\ : InMux
    port map (
            O => \N__40879\,
            I => \N__40831\
        );

    \I__9089\ : LocalMux
    port map (
            O => \N__40876\,
            I => \N__40826\
        );

    \I__9088\ : LocalMux
    port map (
            O => \N__40873\,
            I => \N__40826\
        );

    \I__9087\ : InMux
    port map (
            O => \N__40872\,
            I => \N__40821\
        );

    \I__9086\ : InMux
    port map (
            O => \N__40869\,
            I => \N__40821\
        );

    \I__9085\ : InMux
    port map (
            O => \N__40866\,
            I => \N__40812\
        );

    \I__9084\ : InMux
    port map (
            O => \N__40863\,
            I => \N__40812\
        );

    \I__9083\ : InMux
    port map (
            O => \N__40862\,
            I => \N__40812\
        );

    \I__9082\ : InMux
    port map (
            O => \N__40861\,
            I => \N__40812\
        );

    \I__9081\ : InMux
    port map (
            O => \N__40860\,
            I => \N__40803\
        );

    \I__9080\ : InMux
    port map (
            O => \N__40859\,
            I => \N__40803\
        );

    \I__9079\ : InMux
    port map (
            O => \N__40858\,
            I => \N__40803\
        );

    \I__9078\ : InMux
    port map (
            O => \N__40857\,
            I => \N__40803\
        );

    \I__9077\ : InMux
    port map (
            O => \N__40854\,
            I => \N__40795\
        );

    \I__9076\ : InMux
    port map (
            O => \N__40853\,
            I => \N__40795\
        );

    \I__9075\ : InMux
    port map (
            O => \N__40852\,
            I => \N__40795\
        );

    \I__9074\ : LocalMux
    port map (
            O => \N__40849\,
            I => \N__40792\
        );

    \I__9073\ : LocalMux
    port map (
            O => \N__40842\,
            I => \N__40789\
        );

    \I__9072\ : LocalMux
    port map (
            O => \N__40839\,
            I => \N__40784\
        );

    \I__9071\ : Span4Mux_h
    port map (
            O => \N__40836\,
            I => \N__40784\
        );

    \I__9070\ : LocalMux
    port map (
            O => \N__40831\,
            I => \N__40775\
        );

    \I__9069\ : Span4Mux_h
    port map (
            O => \N__40826\,
            I => \N__40775\
        );

    \I__9068\ : LocalMux
    port map (
            O => \N__40821\,
            I => \N__40775\
        );

    \I__9067\ : LocalMux
    port map (
            O => \N__40812\,
            I => \N__40775\
        );

    \I__9066\ : LocalMux
    port map (
            O => \N__40803\,
            I => \N__40772\
        );

    \I__9065\ : InMux
    port map (
            O => \N__40802\,
            I => \N__40769\
        );

    \I__9064\ : LocalMux
    port map (
            O => \N__40795\,
            I => \N__40766\
        );

    \I__9063\ : Span4Mux_v
    port map (
            O => \N__40792\,
            I => \N__40763\
        );

    \I__9062\ : Span4Mux_h
    port map (
            O => \N__40789\,
            I => \N__40760\
        );

    \I__9061\ : Span4Mux_v
    port map (
            O => \N__40784\,
            I => \N__40755\
        );

    \I__9060\ : Span4Mux_v
    port map (
            O => \N__40775\,
            I => \N__40755\
        );

    \I__9059\ : Span4Mux_h
    port map (
            O => \N__40772\,
            I => \N__40752\
        );

    \I__9058\ : LocalMux
    port map (
            O => \N__40769\,
            I => \phase_controller_slave.start_timer_hcZ0\
        );

    \I__9057\ : Odrv12
    port map (
            O => \N__40766\,
            I => \phase_controller_slave.start_timer_hcZ0\
        );

    \I__9056\ : Odrv4
    port map (
            O => \N__40763\,
            I => \phase_controller_slave.start_timer_hcZ0\
        );

    \I__9055\ : Odrv4
    port map (
            O => \N__40760\,
            I => \phase_controller_slave.start_timer_hcZ0\
        );

    \I__9054\ : Odrv4
    port map (
            O => \N__40755\,
            I => \phase_controller_slave.start_timer_hcZ0\
        );

    \I__9053\ : Odrv4
    port map (
            O => \N__40752\,
            I => \phase_controller_slave.start_timer_hcZ0\
        );

    \I__9052\ : InMux
    port map (
            O => \N__40739\,
            I => \N__40735\
        );

    \I__9051\ : InMux
    port map (
            O => \N__40738\,
            I => \N__40732\
        );

    \I__9050\ : LocalMux
    port map (
            O => \N__40735\,
            I => \N__40729\
        );

    \I__9049\ : LocalMux
    port map (
            O => \N__40732\,
            I => \N__40725\
        );

    \I__9048\ : Span4Mux_v
    port map (
            O => \N__40729\,
            I => \N__40722\
        );

    \I__9047\ : InMux
    port map (
            O => \N__40728\,
            I => \N__40719\
        );

    \I__9046\ : Span4Mux_h
    port map (
            O => \N__40725\,
            I => \N__40713\
        );

    \I__9045\ : Span4Mux_h
    port map (
            O => \N__40722\,
            I => \N__40708\
        );

    \I__9044\ : LocalMux
    port map (
            O => \N__40719\,
            I => \N__40708\
        );

    \I__9043\ : InMux
    port map (
            O => \N__40718\,
            I => \N__40705\
        );

    \I__9042\ : InMux
    port map (
            O => \N__40717\,
            I => \N__40700\
        );

    \I__9041\ : InMux
    port map (
            O => \N__40716\,
            I => \N__40700\
        );

    \I__9040\ : Odrv4
    port map (
            O => \N__40713\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__9039\ : Odrv4
    port map (
            O => \N__40708\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__9038\ : LocalMux
    port map (
            O => \N__40705\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__9037\ : LocalMux
    port map (
            O => \N__40700\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__9036\ : CascadeMux
    port map (
            O => \N__40691\,
            I => \N__40687\
        );

    \I__9035\ : CascadeMux
    port map (
            O => \N__40690\,
            I => \N__40684\
        );

    \I__9034\ : InMux
    port map (
            O => \N__40687\,
            I => \N__40674\
        );

    \I__9033\ : InMux
    port map (
            O => \N__40684\,
            I => \N__40674\
        );

    \I__9032\ : InMux
    port map (
            O => \N__40683\,
            I => \N__40671\
        );

    \I__9031\ : InMux
    port map (
            O => \N__40682\,
            I => \N__40668\
        );

    \I__9030\ : InMux
    port map (
            O => \N__40681\,
            I => \N__40656\
        );

    \I__9029\ : InMux
    port map (
            O => \N__40680\,
            I => \N__40656\
        );

    \I__9028\ : InMux
    port map (
            O => \N__40679\,
            I => \N__40656\
        );

    \I__9027\ : LocalMux
    port map (
            O => \N__40674\,
            I => \N__40650\
        );

    \I__9026\ : LocalMux
    port map (
            O => \N__40671\,
            I => \N__40650\
        );

    \I__9025\ : LocalMux
    port map (
            O => \N__40668\,
            I => \N__40647\
        );

    \I__9024\ : CascadeMux
    port map (
            O => \N__40667\,
            I => \N__40644\
        );

    \I__9023\ : CascadeMux
    port map (
            O => \N__40666\,
            I => \N__40641\
        );

    \I__9022\ : CascadeMux
    port map (
            O => \N__40665\,
            I => \N__40637\
        );

    \I__9021\ : InMux
    port map (
            O => \N__40664\,
            I => \N__40625\
        );

    \I__9020\ : InMux
    port map (
            O => \N__40663\,
            I => \N__40622\
        );

    \I__9019\ : LocalMux
    port map (
            O => \N__40656\,
            I => \N__40619\
        );

    \I__9018\ : InMux
    port map (
            O => \N__40655\,
            I => \N__40616\
        );

    \I__9017\ : Span4Mux_v
    port map (
            O => \N__40650\,
            I => \N__40611\
        );

    \I__9016\ : Span4Mux_v
    port map (
            O => \N__40647\,
            I => \N__40611\
        );

    \I__9015\ : InMux
    port map (
            O => \N__40644\,
            I => \N__40604\
        );

    \I__9014\ : InMux
    port map (
            O => \N__40641\,
            I => \N__40604\
        );

    \I__9013\ : InMux
    port map (
            O => \N__40640\,
            I => \N__40604\
        );

    \I__9012\ : InMux
    port map (
            O => \N__40637\,
            I => \N__40595\
        );

    \I__9011\ : InMux
    port map (
            O => \N__40636\,
            I => \N__40595\
        );

    \I__9010\ : InMux
    port map (
            O => \N__40635\,
            I => \N__40595\
        );

    \I__9009\ : InMux
    port map (
            O => \N__40634\,
            I => \N__40595\
        );

    \I__9008\ : InMux
    port map (
            O => \N__40633\,
            I => \N__40588\
        );

    \I__9007\ : InMux
    port map (
            O => \N__40632\,
            I => \N__40588\
        );

    \I__9006\ : InMux
    port map (
            O => \N__40631\,
            I => \N__40588\
        );

    \I__9005\ : InMux
    port map (
            O => \N__40630\,
            I => \N__40583\
        );

    \I__9004\ : InMux
    port map (
            O => \N__40629\,
            I => \N__40583\
        );

    \I__9003\ : InMux
    port map (
            O => \N__40628\,
            I => \N__40580\
        );

    \I__9002\ : LocalMux
    port map (
            O => \N__40625\,
            I => \N__40572\
        );

    \I__9001\ : LocalMux
    port map (
            O => \N__40622\,
            I => \N__40572\
        );

    \I__9000\ : Span4Mux_v
    port map (
            O => \N__40619\,
            I => \N__40572\
        );

    \I__8999\ : LocalMux
    port map (
            O => \N__40616\,
            I => \N__40569\
        );

    \I__8998\ : Span4Mux_v
    port map (
            O => \N__40611\,
            I => \N__40564\
        );

    \I__8997\ : LocalMux
    port map (
            O => \N__40604\,
            I => \N__40564\
        );

    \I__8996\ : LocalMux
    port map (
            O => \N__40595\,
            I => \N__40557\
        );

    \I__8995\ : LocalMux
    port map (
            O => \N__40588\,
            I => \N__40557\
        );

    \I__8994\ : LocalMux
    port map (
            O => \N__40583\,
            I => \N__40557\
        );

    \I__8993\ : LocalMux
    port map (
            O => \N__40580\,
            I => \N__40554\
        );

    \I__8992\ : InMux
    port map (
            O => \N__40579\,
            I => \N__40551\
        );

    \I__8991\ : Span4Mux_v
    port map (
            O => \N__40572\,
            I => \N__40548\
        );

    \I__8990\ : Span4Mux_h
    port map (
            O => \N__40569\,
            I => \N__40543\
        );

    \I__8989\ : Span4Mux_h
    port map (
            O => \N__40564\,
            I => \N__40543\
        );

    \I__8988\ : Span4Mux_v
    port map (
            O => \N__40557\,
            I => \N__40538\
        );

    \I__8987\ : Span4Mux_h
    port map (
            O => \N__40554\,
            I => \N__40538\
        );

    \I__8986\ : LocalMux
    port map (
            O => \N__40551\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__8985\ : Odrv4
    port map (
            O => \N__40548\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__8984\ : Odrv4
    port map (
            O => \N__40543\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__8983\ : Odrv4
    port map (
            O => \N__40538\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__8982\ : IoInMux
    port map (
            O => \N__40529\,
            I => \N__40526\
        );

    \I__8981\ : LocalMux
    port map (
            O => \N__40526\,
            I => \N__40523\
        );

    \I__8980\ : Span4Mux_s2_v
    port map (
            O => \N__40523\,
            I => \N__40519\
        );

    \I__8979\ : CEMux
    port map (
            O => \N__40522\,
            I => \N__40515\
        );

    \I__8978\ : Span4Mux_h
    port map (
            O => \N__40519\,
            I => \N__40511\
        );

    \I__8977\ : CEMux
    port map (
            O => \N__40518\,
            I => \N__40508\
        );

    \I__8976\ : LocalMux
    port map (
            O => \N__40515\,
            I => \N__40505\
        );

    \I__8975\ : CEMux
    port map (
            O => \N__40514\,
            I => \N__40502\
        );

    \I__8974\ : Span4Mux_v
    port map (
            O => \N__40511\,
            I => \N__40499\
        );

    \I__8973\ : LocalMux
    port map (
            O => \N__40508\,
            I => \N__40496\
        );

    \I__8972\ : Span4Mux_v
    port map (
            O => \N__40505\,
            I => \N__40491\
        );

    \I__8971\ : LocalMux
    port map (
            O => \N__40502\,
            I => \N__40491\
        );

    \I__8970\ : Span4Mux_v
    port map (
            O => \N__40499\,
            I => \N__40488\
        );

    \I__8969\ : Sp12to4
    port map (
            O => \N__40496\,
            I => \N__40485\
        );

    \I__8968\ : Span4Mux_v
    port map (
            O => \N__40491\,
            I => \N__40482\
        );

    \I__8967\ : Odrv4
    port map (
            O => \N__40488\,
            I => red_c_i
        );

    \I__8966\ : Odrv12
    port map (
            O => \N__40485\,
            I => red_c_i
        );

    \I__8965\ : Odrv4
    port map (
            O => \N__40482\,
            I => red_c_i
        );

    \I__8964\ : CascadeMux
    port map (
            O => \N__40475\,
            I => \N__40472\
        );

    \I__8963\ : InMux
    port map (
            O => \N__40472\,
            I => \N__40469\
        );

    \I__8962\ : LocalMux
    port map (
            O => \N__40469\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_17\
        );

    \I__8961\ : CascadeMux
    port map (
            O => \N__40466\,
            I => \N__40463\
        );

    \I__8960\ : InMux
    port map (
            O => \N__40463\,
            I => \N__40460\
        );

    \I__8959\ : LocalMux
    port map (
            O => \N__40460\,
            I => \N__40457\
        );

    \I__8958\ : Odrv4
    port map (
            O => \N__40457\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_8\
        );

    \I__8957\ : InMux
    port map (
            O => \N__40454\,
            I => \N__40450\
        );

    \I__8956\ : InMux
    port map (
            O => \N__40453\,
            I => \N__40447\
        );

    \I__8955\ : LocalMux
    port map (
            O => \N__40450\,
            I => \N__40444\
        );

    \I__8954\ : LocalMux
    port map (
            O => \N__40447\,
            I => \N__40441\
        );

    \I__8953\ : Span4Mux_v
    port map (
            O => \N__40444\,
            I => \N__40436\
        );

    \I__8952\ : Span4Mux_v
    port map (
            O => \N__40441\,
            I => \N__40433\
        );

    \I__8951\ : InMux
    port map (
            O => \N__40440\,
            I => \N__40430\
        );

    \I__8950\ : CascadeMux
    port map (
            O => \N__40439\,
            I => \N__40426\
        );

    \I__8949\ : Span4Mux_v
    port map (
            O => \N__40436\,
            I => \N__40419\
        );

    \I__8948\ : Span4Mux_h
    port map (
            O => \N__40433\,
            I => \N__40419\
        );

    \I__8947\ : LocalMux
    port map (
            O => \N__40430\,
            I => \N__40419\
        );

    \I__8946\ : InMux
    port map (
            O => \N__40429\,
            I => \N__40414\
        );

    \I__8945\ : InMux
    port map (
            O => \N__40426\,
            I => \N__40414\
        );

    \I__8944\ : Odrv4
    port map (
            O => \N__40419\,
            I => measured_delay_hc_16
        );

    \I__8943\ : LocalMux
    port map (
            O => \N__40414\,
            I => measured_delay_hc_16
        );

    \I__8942\ : CascadeMux
    port map (
            O => \N__40409\,
            I => \N__40406\
        );

    \I__8941\ : InMux
    port map (
            O => \N__40406\,
            I => \N__40403\
        );

    \I__8940\ : LocalMux
    port map (
            O => \N__40403\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_16\
        );

    \I__8939\ : InMux
    port map (
            O => \N__40400\,
            I => \N__40397\
        );

    \I__8938\ : LocalMux
    port map (
            O => \N__40397\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_18\
        );

    \I__8937\ : InMux
    port map (
            O => \N__40394\,
            I => \N__40390\
        );

    \I__8936\ : InMux
    port map (
            O => \N__40393\,
            I => \N__40386\
        );

    \I__8935\ : LocalMux
    port map (
            O => \N__40390\,
            I => \N__40383\
        );

    \I__8934\ : InMux
    port map (
            O => \N__40389\,
            I => \N__40380\
        );

    \I__8933\ : LocalMux
    port map (
            O => \N__40386\,
            I => \N__40377\
        );

    \I__8932\ : Span4Mux_h
    port map (
            O => \N__40383\,
            I => \N__40374\
        );

    \I__8931\ : LocalMux
    port map (
            O => \N__40380\,
            I => \N__40371\
        );

    \I__8930\ : Span4Mux_h
    port map (
            O => \N__40377\,
            I => \N__40368\
        );

    \I__8929\ : Span4Mux_v
    port map (
            O => \N__40374\,
            I => \N__40365\
        );

    \I__8928\ : Span4Mux_h
    port map (
            O => \N__40371\,
            I => \N__40360\
        );

    \I__8927\ : Span4Mux_v
    port map (
            O => \N__40368\,
            I => \N__40360\
        );

    \I__8926\ : Odrv4
    port map (
            O => \N__40365\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1\
        );

    \I__8925\ : Odrv4
    port map (
            O => \N__40360\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1\
        );

    \I__8924\ : CascadeMux
    port map (
            O => \N__40355\,
            I => \N__40352\
        );

    \I__8923\ : InMux
    port map (
            O => \N__40352\,
            I => \N__40349\
        );

    \I__8922\ : LocalMux
    port map (
            O => \N__40349\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_19\
        );

    \I__8921\ : InMux
    port map (
            O => \N__40346\,
            I => \N__40337\
        );

    \I__8920\ : InMux
    port map (
            O => \N__40345\,
            I => \N__40337\
        );

    \I__8919\ : InMux
    port map (
            O => \N__40344\,
            I => \N__40332\
        );

    \I__8918\ : CascadeMux
    port map (
            O => \N__40343\,
            I => \N__40329\
        );

    \I__8917\ : InMux
    port map (
            O => \N__40342\,
            I => \N__40323\
        );

    \I__8916\ : LocalMux
    port map (
            O => \N__40337\,
            I => \N__40320\
        );

    \I__8915\ : InMux
    port map (
            O => \N__40336\,
            I => \N__40311\
        );

    \I__8914\ : InMux
    port map (
            O => \N__40335\,
            I => \N__40311\
        );

    \I__8913\ : LocalMux
    port map (
            O => \N__40332\,
            I => \N__40308\
        );

    \I__8912\ : InMux
    port map (
            O => \N__40329\,
            I => \N__40299\
        );

    \I__8911\ : InMux
    port map (
            O => \N__40328\,
            I => \N__40299\
        );

    \I__8910\ : InMux
    port map (
            O => \N__40327\,
            I => \N__40299\
        );

    \I__8909\ : InMux
    port map (
            O => \N__40326\,
            I => \N__40299\
        );

    \I__8908\ : LocalMux
    port map (
            O => \N__40323\,
            I => \N__40296\
        );

    \I__8907\ : Span4Mux_h
    port map (
            O => \N__40320\,
            I => \N__40293\
        );

    \I__8906\ : InMux
    port map (
            O => \N__40319\,
            I => \N__40284\
        );

    \I__8905\ : InMux
    port map (
            O => \N__40318\,
            I => \N__40284\
        );

    \I__8904\ : InMux
    port map (
            O => \N__40317\,
            I => \N__40284\
        );

    \I__8903\ : InMux
    port map (
            O => \N__40316\,
            I => \N__40284\
        );

    \I__8902\ : LocalMux
    port map (
            O => \N__40311\,
            I => \N__40281\
        );

    \I__8901\ : Span4Mux_v
    port map (
            O => \N__40308\,
            I => \N__40278\
        );

    \I__8900\ : LocalMux
    port map (
            O => \N__40299\,
            I => \N__40275\
        );

    \I__8899\ : Span4Mux_v
    port map (
            O => \N__40296\,
            I => \N__40272\
        );

    \I__8898\ : Span4Mux_v
    port map (
            O => \N__40293\,
            I => \N__40269\
        );

    \I__8897\ : LocalMux
    port map (
            O => \N__40284\,
            I => \N__40262\
        );

    \I__8896\ : Span4Mux_v
    port map (
            O => \N__40281\,
            I => \N__40262\
        );

    \I__8895\ : Span4Mux_v
    port map (
            O => \N__40278\,
            I => \N__40262\
        );

    \I__8894\ : Span12Mux_h
    port map (
            O => \N__40275\,
            I => \N__40259\
        );

    \I__8893\ : Odrv4
    port map (
            O => \N__40272\,
            I => \phase_controller_inst1.stoper_hc.un2_startlt31\
        );

    \I__8892\ : Odrv4
    port map (
            O => \N__40269\,
            I => \phase_controller_inst1.stoper_hc.un2_startlt31\
        );

    \I__8891\ : Odrv4
    port map (
            O => \N__40262\,
            I => \phase_controller_inst1.stoper_hc.un2_startlt31\
        );

    \I__8890\ : Odrv12
    port map (
            O => \N__40259\,
            I => \phase_controller_inst1.stoper_hc.un2_startlt31\
        );

    \I__8889\ : InMux
    port map (
            O => \N__40250\,
            I => \N__40245\
        );

    \I__8888\ : InMux
    port map (
            O => \N__40249\,
            I => \N__40242\
        );

    \I__8887\ : InMux
    port map (
            O => \N__40248\,
            I => \N__40239\
        );

    \I__8886\ : LocalMux
    port map (
            O => \N__40245\,
            I => \N__40236\
        );

    \I__8885\ : LocalMux
    port map (
            O => \N__40242\,
            I => \N__40233\
        );

    \I__8884\ : LocalMux
    port map (
            O => \N__40239\,
            I => \N__40230\
        );

    \I__8883\ : Span4Mux_v
    port map (
            O => \N__40236\,
            I => \N__40225\
        );

    \I__8882\ : Span4Mux_h
    port map (
            O => \N__40233\,
            I => \N__40225\
        );

    \I__8881\ : Span12Mux_v
    port map (
            O => \N__40230\,
            I => \N__40222\
        );

    \I__8880\ : Odrv4
    port map (
            O => \N__40225\,
            I => measured_delay_tr_6
        );

    \I__8879\ : Odrv12
    port map (
            O => \N__40222\,
            I => measured_delay_tr_6
        );

    \I__8878\ : InMux
    port map (
            O => \N__40217\,
            I => \N__40210\
        );

    \I__8877\ : InMux
    port map (
            O => \N__40216\,
            I => \N__40210\
        );

    \I__8876\ : CascadeMux
    port map (
            O => \N__40215\,
            I => \N__40207\
        );

    \I__8875\ : LocalMux
    port map (
            O => \N__40210\,
            I => \N__40202\
        );

    \I__8874\ : InMux
    port map (
            O => \N__40207\,
            I => \N__40195\
        );

    \I__8873\ : InMux
    port map (
            O => \N__40206\,
            I => \N__40195\
        );

    \I__8872\ : InMux
    port map (
            O => \N__40205\,
            I => \N__40195\
        );

    \I__8871\ : Span4Mux_v
    port map (
            O => \N__40202\,
            I => \N__40192\
        );

    \I__8870\ : LocalMux
    port map (
            O => \N__40195\,
            I => \N__40189\
        );

    \I__8869\ : Span4Mux_h
    port map (
            O => \N__40192\,
            I => \N__40186\
        );

    \I__8868\ : Span4Mux_v
    port map (
            O => \N__40189\,
            I => \N__40183\
        );

    \I__8867\ : Odrv4
    port map (
            O => \N__40186\,
            I => measured_delay_tr_3
        );

    \I__8866\ : Odrv4
    port map (
            O => \N__40183\,
            I => measured_delay_tr_3
        );

    \I__8865\ : InMux
    port map (
            O => \N__40178\,
            I => \N__40174\
        );

    \I__8864\ : CascadeMux
    port map (
            O => \N__40177\,
            I => \N__40171\
        );

    \I__8863\ : LocalMux
    port map (
            O => \N__40174\,
            I => \N__40168\
        );

    \I__8862\ : InMux
    port map (
            O => \N__40171\,
            I => \N__40165\
        );

    \I__8861\ : Span4Mux_v
    port map (
            O => \N__40168\,
            I => \N__40161\
        );

    \I__8860\ : LocalMux
    port map (
            O => \N__40165\,
            I => \N__40158\
        );

    \I__8859\ : InMux
    port map (
            O => \N__40164\,
            I => \N__40155\
        );

    \I__8858\ : Span4Mux_h
    port map (
            O => \N__40161\,
            I => \N__40150\
        );

    \I__8857\ : Span4Mux_v
    port map (
            O => \N__40158\,
            I => \N__40150\
        );

    \I__8856\ : LocalMux
    port map (
            O => \N__40155\,
            I => \N__40147\
        );

    \I__8855\ : Sp12to4
    port map (
            O => \N__40150\,
            I => \N__40142\
        );

    \I__8854\ : Span12Mux_h
    port map (
            O => \N__40147\,
            I => \N__40142\
        );

    \I__8853\ : Odrv12
    port map (
            O => \N__40142\,
            I => measured_delay_tr_5
        );

    \I__8852\ : InMux
    port map (
            O => \N__40139\,
            I => \N__40135\
        );

    \I__8851\ : InMux
    port map (
            O => \N__40138\,
            I => \N__40132\
        );

    \I__8850\ : LocalMux
    port map (
            O => \N__40135\,
            I => \N__40129\
        );

    \I__8849\ : LocalMux
    port map (
            O => \N__40132\,
            I => \N__40126\
        );

    \I__8848\ : Odrv12
    port map (
            O => \N__40129\,
            I => \delay_measurement_inst.elapsed_time_tr_1\
        );

    \I__8847\ : Odrv4
    port map (
            O => \N__40126\,
            I => \delay_measurement_inst.elapsed_time_tr_1\
        );

    \I__8846\ : CascadeMux
    port map (
            O => \N__40121\,
            I => \N__40118\
        );

    \I__8845\ : InMux
    port map (
            O => \N__40118\,
            I => \N__40114\
        );

    \I__8844\ : InMux
    port map (
            O => \N__40117\,
            I => \N__40111\
        );

    \I__8843\ : LocalMux
    port map (
            O => \N__40114\,
            I => \N__40108\
        );

    \I__8842\ : LocalMux
    port map (
            O => \N__40111\,
            I => \N__40105\
        );

    \I__8841\ : Span4Mux_v
    port map (
            O => \N__40108\,
            I => \N__40102\
        );

    \I__8840\ : Span4Mux_v
    port map (
            O => \N__40105\,
            I => \N__40099\
        );

    \I__8839\ : Odrv4
    port map (
            O => \N__40102\,
            I => measured_delay_tr_1
        );

    \I__8838\ : Odrv4
    port map (
            O => \N__40099\,
            I => measured_delay_tr_1
        );

    \I__8837\ : InMux
    port map (
            O => \N__40094\,
            I => \N__40089\
        );

    \I__8836\ : InMux
    port map (
            O => \N__40093\,
            I => \N__40084\
        );

    \I__8835\ : InMux
    port map (
            O => \N__40092\,
            I => \N__40084\
        );

    \I__8834\ : LocalMux
    port map (
            O => \N__40089\,
            I => \N__40081\
        );

    \I__8833\ : LocalMux
    port map (
            O => \N__40084\,
            I => \N__40078\
        );

    \I__8832\ : Span4Mux_h
    port map (
            O => \N__40081\,
            I => \N__40075\
        );

    \I__8831\ : Span4Mux_v
    port map (
            O => \N__40078\,
            I => \N__40072\
        );

    \I__8830\ : Odrv4
    port map (
            O => \N__40075\,
            I => measured_delay_tr_2
        );

    \I__8829\ : Odrv4
    port map (
            O => \N__40072\,
            I => measured_delay_tr_2
        );

    \I__8828\ : InMux
    port map (
            O => \N__40067\,
            I => \N__40061\
        );

    \I__8827\ : InMux
    port map (
            O => \N__40066\,
            I => \N__40056\
        );

    \I__8826\ : InMux
    port map (
            O => \N__40065\,
            I => \N__40056\
        );

    \I__8825\ : InMux
    port map (
            O => \N__40064\,
            I => \N__40053\
        );

    \I__8824\ : LocalMux
    port map (
            O => \N__40061\,
            I => \N__40050\
        );

    \I__8823\ : LocalMux
    port map (
            O => \N__40056\,
            I => \N__40047\
        );

    \I__8822\ : LocalMux
    port map (
            O => \N__40053\,
            I => \N__40044\
        );

    \I__8821\ : Span4Mux_h
    port map (
            O => \N__40050\,
            I => \N__40041\
        );

    \I__8820\ : Span12Mux_h
    port map (
            O => \N__40047\,
            I => \N__40036\
        );

    \I__8819\ : Span4Mux_h
    port map (
            O => \N__40044\,
            I => \N__40031\
        );

    \I__8818\ : Span4Mux_v
    port map (
            O => \N__40041\,
            I => \N__40031\
        );

    \I__8817\ : InMux
    port map (
            O => \N__40040\,
            I => \N__40026\
        );

    \I__8816\ : InMux
    port map (
            O => \N__40039\,
            I => \N__40026\
        );

    \I__8815\ : Odrv12
    port map (
            O => \N__40036\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__8814\ : Odrv4
    port map (
            O => \N__40031\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__8813\ : LocalMux
    port map (
            O => \N__40026\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__8812\ : CascadeMux
    port map (
            O => \N__40019\,
            I => \N__40008\
        );

    \I__8811\ : CascadeMux
    port map (
            O => \N__40018\,
            I => \N__40003\
        );

    \I__8810\ : CascadeMux
    port map (
            O => \N__40017\,
            I => \N__39998\
        );

    \I__8809\ : CascadeMux
    port map (
            O => \N__40016\,
            I => \N__39995\
        );

    \I__8808\ : CascadeMux
    port map (
            O => \N__40015\,
            I => \N__39991\
        );

    \I__8807\ : CascadeMux
    port map (
            O => \N__40014\,
            I => \N__39985\
        );

    \I__8806\ : CascadeMux
    port map (
            O => \N__40013\,
            I => \N__39982\
        );

    \I__8805\ : CascadeMux
    port map (
            O => \N__40012\,
            I => \N__39979\
        );

    \I__8804\ : InMux
    port map (
            O => \N__40011\,
            I => \N__39972\
        );

    \I__8803\ : InMux
    port map (
            O => \N__40008\,
            I => \N__39972\
        );

    \I__8802\ : CascadeMux
    port map (
            O => \N__40007\,
            I => \N__39969\
        );

    \I__8801\ : CascadeMux
    port map (
            O => \N__40006\,
            I => \N__39966\
        );

    \I__8800\ : InMux
    port map (
            O => \N__40003\,
            I => \N__39963\
        );

    \I__8799\ : InMux
    port map (
            O => \N__40002\,
            I => \N__39946\
        );

    \I__8798\ : InMux
    port map (
            O => \N__40001\,
            I => \N__39946\
        );

    \I__8797\ : InMux
    port map (
            O => \N__39998\,
            I => \N__39946\
        );

    \I__8796\ : InMux
    port map (
            O => \N__39995\,
            I => \N__39946\
        );

    \I__8795\ : InMux
    port map (
            O => \N__39994\,
            I => \N__39946\
        );

    \I__8794\ : InMux
    port map (
            O => \N__39991\,
            I => \N__39946\
        );

    \I__8793\ : InMux
    port map (
            O => \N__39990\,
            I => \N__39946\
        );

    \I__8792\ : InMux
    port map (
            O => \N__39989\,
            I => \N__39933\
        );

    \I__8791\ : InMux
    port map (
            O => \N__39988\,
            I => \N__39933\
        );

    \I__8790\ : InMux
    port map (
            O => \N__39985\,
            I => \N__39933\
        );

    \I__8789\ : InMux
    port map (
            O => \N__39982\,
            I => \N__39933\
        );

    \I__8788\ : InMux
    port map (
            O => \N__39979\,
            I => \N__39933\
        );

    \I__8787\ : InMux
    port map (
            O => \N__39978\,
            I => \N__39933\
        );

    \I__8786\ : CascadeMux
    port map (
            O => \N__39977\,
            I => \N__39929\
        );

    \I__8785\ : LocalMux
    port map (
            O => \N__39972\,
            I => \N__39925\
        );

    \I__8784\ : InMux
    port map (
            O => \N__39969\,
            I => \N__39920\
        );

    \I__8783\ : InMux
    port map (
            O => \N__39966\,
            I => \N__39920\
        );

    \I__8782\ : LocalMux
    port map (
            O => \N__39963\,
            I => \N__39917\
        );

    \I__8781\ : InMux
    port map (
            O => \N__39962\,
            I => \N__39914\
        );

    \I__8780\ : InMux
    port map (
            O => \N__39961\,
            I => \N__39911\
        );

    \I__8779\ : LocalMux
    port map (
            O => \N__39946\,
            I => \N__39907\
        );

    \I__8778\ : LocalMux
    port map (
            O => \N__39933\,
            I => \N__39904\
        );

    \I__8777\ : InMux
    port map (
            O => \N__39932\,
            I => \N__39899\
        );

    \I__8776\ : InMux
    port map (
            O => \N__39929\,
            I => \N__39899\
        );

    \I__8775\ : CascadeMux
    port map (
            O => \N__39928\,
            I => \N__39896\
        );

    \I__8774\ : Span4Mux_v
    port map (
            O => \N__39925\,
            I => \N__39893\
        );

    \I__8773\ : LocalMux
    port map (
            O => \N__39920\,
            I => \N__39890\
        );

    \I__8772\ : Span4Mux_v
    port map (
            O => \N__39917\,
            I => \N__39883\
        );

    \I__8771\ : LocalMux
    port map (
            O => \N__39914\,
            I => \N__39883\
        );

    \I__8770\ : LocalMux
    port map (
            O => \N__39911\,
            I => \N__39883\
        );

    \I__8769\ : InMux
    port map (
            O => \N__39910\,
            I => \N__39880\
        );

    \I__8768\ : Span4Mux_v
    port map (
            O => \N__39907\,
            I => \N__39873\
        );

    \I__8767\ : Span4Mux_v
    port map (
            O => \N__39904\,
            I => \N__39873\
        );

    \I__8766\ : LocalMux
    port map (
            O => \N__39899\,
            I => \N__39873\
        );

    \I__8765\ : InMux
    port map (
            O => \N__39896\,
            I => \N__39870\
        );

    \I__8764\ : Span4Mux_h
    port map (
            O => \N__39893\,
            I => \N__39863\
        );

    \I__8763\ : Span4Mux_h
    port map (
            O => \N__39890\,
            I => \N__39863\
        );

    \I__8762\ : Span4Mux_h
    port map (
            O => \N__39883\,
            I => \N__39863\
        );

    \I__8761\ : LocalMux
    port map (
            O => \N__39880\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__8760\ : Odrv4
    port map (
            O => \N__39873\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__8759\ : LocalMux
    port map (
            O => \N__39870\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__8758\ : Odrv4
    port map (
            O => \N__39863\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__8757\ : CascadeMux
    port map (
            O => \N__39854\,
            I => \N__39842\
        );

    \I__8756\ : CascadeMux
    port map (
            O => \N__39853\,
            I => \N__39839\
        );

    \I__8755\ : CascadeMux
    port map (
            O => \N__39852\,
            I => \N__39836\
        );

    \I__8754\ : CascadeMux
    port map (
            O => \N__39851\,
            I => \N__39833\
        );

    \I__8753\ : CascadeMux
    port map (
            O => \N__39850\,
            I => \N__39830\
        );

    \I__8752\ : CascadeMux
    port map (
            O => \N__39849\,
            I => \N__39827\
        );

    \I__8751\ : CascadeMux
    port map (
            O => \N__39848\,
            I => \N__39824\
        );

    \I__8750\ : InMux
    port map (
            O => \N__39847\,
            I => \N__39813\
        );

    \I__8749\ : InMux
    port map (
            O => \N__39846\,
            I => \N__39813\
        );

    \I__8748\ : InMux
    port map (
            O => \N__39845\,
            I => \N__39808\
        );

    \I__8747\ : InMux
    port map (
            O => \N__39842\,
            I => \N__39799\
        );

    \I__8746\ : InMux
    port map (
            O => \N__39839\,
            I => \N__39799\
        );

    \I__8745\ : InMux
    port map (
            O => \N__39836\,
            I => \N__39799\
        );

    \I__8744\ : InMux
    port map (
            O => \N__39833\,
            I => \N__39799\
        );

    \I__8743\ : InMux
    port map (
            O => \N__39830\,
            I => \N__39792\
        );

    \I__8742\ : InMux
    port map (
            O => \N__39827\,
            I => \N__39792\
        );

    \I__8741\ : InMux
    port map (
            O => \N__39824\,
            I => \N__39792\
        );

    \I__8740\ : InMux
    port map (
            O => \N__39823\,
            I => \N__39785\
        );

    \I__8739\ : InMux
    port map (
            O => \N__39822\,
            I => \N__39785\
        );

    \I__8738\ : InMux
    port map (
            O => \N__39821\,
            I => \N__39785\
        );

    \I__8737\ : InMux
    port map (
            O => \N__39820\,
            I => \N__39778\
        );

    \I__8736\ : InMux
    port map (
            O => \N__39819\,
            I => \N__39778\
        );

    \I__8735\ : InMux
    port map (
            O => \N__39818\,
            I => \N__39778\
        );

    \I__8734\ : LocalMux
    port map (
            O => \N__39813\,
            I => \N__39775\
        );

    \I__8733\ : InMux
    port map (
            O => \N__39812\,
            I => \N__39770\
        );

    \I__8732\ : InMux
    port map (
            O => \N__39811\,
            I => \N__39770\
        );

    \I__8731\ : LocalMux
    port map (
            O => \N__39808\,
            I => \N__39755\
        );

    \I__8730\ : LocalMux
    port map (
            O => \N__39799\,
            I => \N__39755\
        );

    \I__8729\ : LocalMux
    port map (
            O => \N__39792\,
            I => \N__39755\
        );

    \I__8728\ : LocalMux
    port map (
            O => \N__39785\,
            I => \N__39755\
        );

    \I__8727\ : LocalMux
    port map (
            O => \N__39778\,
            I => \N__39755\
        );

    \I__8726\ : Span4Mux_v
    port map (
            O => \N__39775\,
            I => \N__39750\
        );

    \I__8725\ : LocalMux
    port map (
            O => \N__39770\,
            I => \N__39750\
        );

    \I__8724\ : InMux
    port map (
            O => \N__39769\,
            I => \N__39747\
        );

    \I__8723\ : InMux
    port map (
            O => \N__39768\,
            I => \N__39744\
        );

    \I__8722\ : InMux
    port map (
            O => \N__39767\,
            I => \N__39739\
        );

    \I__8721\ : InMux
    port map (
            O => \N__39766\,
            I => \N__39739\
        );

    \I__8720\ : Span4Mux_h
    port map (
            O => \N__39755\,
            I => \N__39735\
        );

    \I__8719\ : Span4Mux_h
    port map (
            O => \N__39750\,
            I => \N__39732\
        );

    \I__8718\ : LocalMux
    port map (
            O => \N__39747\,
            I => \N__39729\
        );

    \I__8717\ : LocalMux
    port map (
            O => \N__39744\,
            I => \N__39726\
        );

    \I__8716\ : LocalMux
    port map (
            O => \N__39739\,
            I => \N__39723\
        );

    \I__8715\ : CascadeMux
    port map (
            O => \N__39738\,
            I => \N__39720\
        );

    \I__8714\ : Span4Mux_v
    port map (
            O => \N__39735\,
            I => \N__39716\
        );

    \I__8713\ : Span4Mux_v
    port map (
            O => \N__39732\,
            I => \N__39713\
        );

    \I__8712\ : Span4Mux_h
    port map (
            O => \N__39729\,
            I => \N__39710\
        );

    \I__8711\ : Span4Mux_v
    port map (
            O => \N__39726\,
            I => \N__39705\
        );

    \I__8710\ : Span4Mux_h
    port map (
            O => \N__39723\,
            I => \N__39705\
        );

    \I__8709\ : InMux
    port map (
            O => \N__39720\,
            I => \N__39700\
        );

    \I__8708\ : InMux
    port map (
            O => \N__39719\,
            I => \N__39700\
        );

    \I__8707\ : Span4Mux_h
    port map (
            O => \N__39716\,
            I => \N__39697\
        );

    \I__8706\ : Span4Mux_h
    port map (
            O => \N__39713\,
            I => \N__39694\
        );

    \I__8705\ : Span4Mux_h
    port map (
            O => \N__39710\,
            I => \N__39689\
        );

    \I__8704\ : Span4Mux_h
    port map (
            O => \N__39705\,
            I => \N__39689\
        );

    \I__8703\ : LocalMux
    port map (
            O => \N__39700\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__8702\ : Odrv4
    port map (
            O => \N__39697\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__8701\ : Odrv4
    port map (
            O => \N__39694\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__8700\ : Odrv4
    port map (
            O => \N__39689\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__8699\ : CascadeMux
    port map (
            O => \N__39680\,
            I => \N__39675\
        );

    \I__8698\ : InMux
    port map (
            O => \N__39679\,
            I => \N__39670\
        );

    \I__8697\ : InMux
    port map (
            O => \N__39678\,
            I => \N__39670\
        );

    \I__8696\ : InMux
    port map (
            O => \N__39675\,
            I => \N__39651\
        );

    \I__8695\ : LocalMux
    port map (
            O => \N__39670\,
            I => \N__39648\
        );

    \I__8694\ : InMux
    port map (
            O => \N__39669\,
            I => \N__39645\
        );

    \I__8693\ : InMux
    port map (
            O => \N__39668\,
            I => \N__39642\
        );

    \I__8692\ : InMux
    port map (
            O => \N__39667\,
            I => \N__39629\
        );

    \I__8691\ : InMux
    port map (
            O => \N__39666\,
            I => \N__39629\
        );

    \I__8690\ : InMux
    port map (
            O => \N__39665\,
            I => \N__39629\
        );

    \I__8689\ : InMux
    port map (
            O => \N__39664\,
            I => \N__39629\
        );

    \I__8688\ : InMux
    port map (
            O => \N__39663\,
            I => \N__39629\
        );

    \I__8687\ : InMux
    port map (
            O => \N__39662\,
            I => \N__39629\
        );

    \I__8686\ : InMux
    port map (
            O => \N__39661\,
            I => \N__39614\
        );

    \I__8685\ : InMux
    port map (
            O => \N__39660\,
            I => \N__39614\
        );

    \I__8684\ : InMux
    port map (
            O => \N__39659\,
            I => \N__39614\
        );

    \I__8683\ : InMux
    port map (
            O => \N__39658\,
            I => \N__39614\
        );

    \I__8682\ : InMux
    port map (
            O => \N__39657\,
            I => \N__39614\
        );

    \I__8681\ : InMux
    port map (
            O => \N__39656\,
            I => \N__39614\
        );

    \I__8680\ : InMux
    port map (
            O => \N__39655\,
            I => \N__39614\
        );

    \I__8679\ : InMux
    port map (
            O => \N__39654\,
            I => \N__39611\
        );

    \I__8678\ : LocalMux
    port map (
            O => \N__39651\,
            I => \N__39601\
        );

    \I__8677\ : Span4Mux_v
    port map (
            O => \N__39648\,
            I => \N__39601\
        );

    \I__8676\ : LocalMux
    port map (
            O => \N__39645\,
            I => \N__39601\
        );

    \I__8675\ : LocalMux
    port map (
            O => \N__39642\,
            I => \N__39594\
        );

    \I__8674\ : LocalMux
    port map (
            O => \N__39629\,
            I => \N__39594\
        );

    \I__8673\ : LocalMux
    port map (
            O => \N__39614\,
            I => \N__39594\
        );

    \I__8672\ : LocalMux
    port map (
            O => \N__39611\,
            I => \N__39591\
        );

    \I__8671\ : InMux
    port map (
            O => \N__39610\,
            I => \N__39588\
        );

    \I__8670\ : InMux
    port map (
            O => \N__39609\,
            I => \N__39583\
        );

    \I__8669\ : InMux
    port map (
            O => \N__39608\,
            I => \N__39583\
        );

    \I__8668\ : Span4Mux_h
    port map (
            O => \N__39601\,
            I => \N__39580\
        );

    \I__8667\ : Span4Mux_h
    port map (
            O => \N__39594\,
            I => \N__39577\
        );

    \I__8666\ : Span4Mux_v
    port map (
            O => \N__39591\,
            I => \N__39570\
        );

    \I__8665\ : LocalMux
    port map (
            O => \N__39588\,
            I => \N__39570\
        );

    \I__8664\ : LocalMux
    port map (
            O => \N__39583\,
            I => \N__39570\
        );

    \I__8663\ : Span4Mux_v
    port map (
            O => \N__39580\,
            I => \N__39565\
        );

    \I__8662\ : Span4Mux_v
    port map (
            O => \N__39577\,
            I => \N__39562\
        );

    \I__8661\ : Span4Mux_h
    port map (
            O => \N__39570\,
            I => \N__39559\
        );

    \I__8660\ : InMux
    port map (
            O => \N__39569\,
            I => \N__39554\
        );

    \I__8659\ : InMux
    port map (
            O => \N__39568\,
            I => \N__39554\
        );

    \I__8658\ : Span4Mux_h
    port map (
            O => \N__39565\,
            I => \N__39551\
        );

    \I__8657\ : Span4Mux_h
    port map (
            O => \N__39562\,
            I => \N__39548\
        );

    \I__8656\ : Span4Mux_h
    port map (
            O => \N__39559\,
            I => \N__39545\
        );

    \I__8655\ : LocalMux
    port map (
            O => \N__39554\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__8654\ : Odrv4
    port map (
            O => \N__39551\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__8653\ : Odrv4
    port map (
            O => \N__39548\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__8652\ : Odrv4
    port map (
            O => \N__39545\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__8651\ : InMux
    port map (
            O => \N__39536\,
            I => \N__39532\
        );

    \I__8650\ : InMux
    port map (
            O => \N__39535\,
            I => \N__39529\
        );

    \I__8649\ : LocalMux
    port map (
            O => \N__39532\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10\
        );

    \I__8648\ : LocalMux
    port map (
            O => \N__39529\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10\
        );

    \I__8647\ : CascadeMux
    port map (
            O => \N__39524\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10_cascade_\
        );

    \I__8646\ : CascadeMux
    port map (
            O => \N__39521\,
            I => \delay_measurement_inst.delay_tr_timer.N_400_cascade_\
        );

    \I__8645\ : CascadeMux
    port map (
            O => \N__39518\,
            I => \delay_measurement_inst.N_394_1_cascade_\
        );

    \I__8644\ : InMux
    port map (
            O => \N__39515\,
            I => \N__39503\
        );

    \I__8643\ : InMux
    port map (
            O => \N__39514\,
            I => \N__39503\
        );

    \I__8642\ : InMux
    port map (
            O => \N__39513\,
            I => \N__39503\
        );

    \I__8641\ : InMux
    port map (
            O => \N__39512\,
            I => \N__39503\
        );

    \I__8640\ : LocalMux
    port map (
            O => \N__39503\,
            I => \delay_measurement_inst.N_394_1\
        );

    \I__8639\ : InMux
    port map (
            O => \N__39500\,
            I => \N__39497\
        );

    \I__8638\ : LocalMux
    port map (
            O => \N__39497\,
            I => \N__39493\
        );

    \I__8637\ : InMux
    port map (
            O => \N__39496\,
            I => \N__39490\
        );

    \I__8636\ : Span4Mux_v
    port map (
            O => \N__39493\,
            I => \N__39486\
        );

    \I__8635\ : LocalMux
    port map (
            O => \N__39490\,
            I => \N__39483\
        );

    \I__8634\ : InMux
    port map (
            O => \N__39489\,
            I => \N__39480\
        );

    \I__8633\ : Odrv4
    port map (
            O => \N__39486\,
            I => measured_delay_tr_12
        );

    \I__8632\ : Odrv4
    port map (
            O => \N__39483\,
            I => measured_delay_tr_12
        );

    \I__8631\ : LocalMux
    port map (
            O => \N__39480\,
            I => measured_delay_tr_12
        );

    \I__8630\ : InMux
    port map (
            O => \N__39473\,
            I => \N__39470\
        );

    \I__8629\ : LocalMux
    port map (
            O => \N__39470\,
            I => \N__39466\
        );

    \I__8628\ : InMux
    port map (
            O => \N__39469\,
            I => \N__39463\
        );

    \I__8627\ : Span4Mux_h
    port map (
            O => \N__39466\,
            I => \N__39459\
        );

    \I__8626\ : LocalMux
    port map (
            O => \N__39463\,
            I => \N__39456\
        );

    \I__8625\ : InMux
    port map (
            O => \N__39462\,
            I => \N__39453\
        );

    \I__8624\ : Odrv4
    port map (
            O => \N__39459\,
            I => measured_delay_tr_10
        );

    \I__8623\ : Odrv4
    port map (
            O => \N__39456\,
            I => measured_delay_tr_10
        );

    \I__8622\ : LocalMux
    port map (
            O => \N__39453\,
            I => measured_delay_tr_10
        );

    \I__8621\ : InMux
    port map (
            O => \N__39446\,
            I => \N__39443\
        );

    \I__8620\ : LocalMux
    port map (
            O => \N__39443\,
            I => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_4\
        );

    \I__8619\ : CascadeMux
    port map (
            O => \N__39440\,
            I => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_6_cascade_\
        );

    \I__8618\ : InMux
    port map (
            O => \N__39437\,
            I => \N__39434\
        );

    \I__8617\ : LocalMux
    port map (
            O => \N__39434\,
            I => \delay_measurement_inst.delay_tr_timer.N_364\
        );

    \I__8616\ : InMux
    port map (
            O => \N__39431\,
            I => \N__39428\
        );

    \I__8615\ : LocalMux
    port map (
            O => \N__39428\,
            I => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_5\
        );

    \I__8614\ : CascadeMux
    port map (
            O => \N__39425\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_6_19_cascade_\
        );

    \I__8613\ : InMux
    port map (
            O => \N__39422\,
            I => \N__39419\
        );

    \I__8612\ : LocalMux
    port map (
            O => \N__39419\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_0_19\
        );

    \I__8611\ : CascadeMux
    port map (
            O => \N__39416\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20_cascade_\
        );

    \I__8610\ : InMux
    port map (
            O => \N__39413\,
            I => \N__39410\
        );

    \I__8609\ : LocalMux
    port map (
            O => \N__39410\,
            I => \delay_measurement_inst.delay_tr_timer.N_409\
        );

    \I__8608\ : InMux
    port map (
            O => \N__39407\,
            I => \N__39402\
        );

    \I__8607\ : InMux
    port map (
            O => \N__39406\,
            I => \N__39398\
        );

    \I__8606\ : CascadeMux
    port map (
            O => \N__39405\,
            I => \N__39395\
        );

    \I__8605\ : LocalMux
    port map (
            O => \N__39402\,
            I => \N__39392\
        );

    \I__8604\ : InMux
    port map (
            O => \N__39401\,
            I => \N__39389\
        );

    \I__8603\ : LocalMux
    port map (
            O => \N__39398\,
            I => \N__39386\
        );

    \I__8602\ : InMux
    port map (
            O => \N__39395\,
            I => \N__39383\
        );

    \I__8601\ : Span4Mux_v
    port map (
            O => \N__39392\,
            I => \N__39380\
        );

    \I__8600\ : LocalMux
    port map (
            O => \N__39389\,
            I => \N__39376\
        );

    \I__8599\ : Span4Mux_v
    port map (
            O => \N__39386\,
            I => \N__39373\
        );

    \I__8598\ : LocalMux
    port map (
            O => \N__39383\,
            I => \N__39368\
        );

    \I__8597\ : Span4Mux_h
    port map (
            O => \N__39380\,
            I => \N__39368\
        );

    \I__8596\ : InMux
    port map (
            O => \N__39379\,
            I => \N__39365\
        );

    \I__8595\ : Span4Mux_v
    port map (
            O => \N__39376\,
            I => \N__39362\
        );

    \I__8594\ : Odrv4
    port map (
            O => \N__39373\,
            I => measured_delay_hc_12
        );

    \I__8593\ : Odrv4
    port map (
            O => \N__39368\,
            I => measured_delay_hc_12
        );

    \I__8592\ : LocalMux
    port map (
            O => \N__39365\,
            I => measured_delay_hc_12
        );

    \I__8591\ : Odrv4
    port map (
            O => \N__39362\,
            I => measured_delay_hc_12
        );

    \I__8590\ : InMux
    port map (
            O => \N__39353\,
            I => \N__39347\
        );

    \I__8589\ : InMux
    port map (
            O => \N__39352\,
            I => \N__39344\
        );

    \I__8588\ : InMux
    port map (
            O => \N__39351\,
            I => \N__39341\
        );

    \I__8587\ : CascadeMux
    port map (
            O => \N__39350\,
            I => \N__39338\
        );

    \I__8586\ : LocalMux
    port map (
            O => \N__39347\,
            I => \N__39335\
        );

    \I__8585\ : LocalMux
    port map (
            O => \N__39344\,
            I => \N__39332\
        );

    \I__8584\ : LocalMux
    port map (
            O => \N__39341\,
            I => \N__39328\
        );

    \I__8583\ : InMux
    port map (
            O => \N__39338\,
            I => \N__39325\
        );

    \I__8582\ : Span4Mux_v
    port map (
            O => \N__39335\,
            I => \N__39322\
        );

    \I__8581\ : Span4Mux_h
    port map (
            O => \N__39332\,
            I => \N__39319\
        );

    \I__8580\ : InMux
    port map (
            O => \N__39331\,
            I => \N__39316\
        );

    \I__8579\ : Span4Mux_v
    port map (
            O => \N__39328\,
            I => \N__39313\
        );

    \I__8578\ : LocalMux
    port map (
            O => \N__39325\,
            I => measured_delay_hc_11
        );

    \I__8577\ : Odrv4
    port map (
            O => \N__39322\,
            I => measured_delay_hc_11
        );

    \I__8576\ : Odrv4
    port map (
            O => \N__39319\,
            I => measured_delay_hc_11
        );

    \I__8575\ : LocalMux
    port map (
            O => \N__39316\,
            I => measured_delay_hc_11
        );

    \I__8574\ : Odrv4
    port map (
            O => \N__39313\,
            I => measured_delay_hc_11
        );

    \I__8573\ : InMux
    port map (
            O => \N__39302\,
            I => \N__39299\
        );

    \I__8572\ : LocalMux
    port map (
            O => \N__39299\,
            I => \N__39296\
        );

    \I__8571\ : Odrv4
    port map (
            O => \N__39296\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9\
        );

    \I__8570\ : InMux
    port map (
            O => \N__39293\,
            I => \N__39290\
        );

    \I__8569\ : LocalMux
    port map (
            O => \N__39290\,
            I => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_5\
        );

    \I__8568\ : CascadeMux
    port map (
            O => \N__39287\,
            I => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_6_cascade_\
        );

    \I__8567\ : InMux
    port map (
            O => \N__39284\,
            I => \N__39281\
        );

    \I__8566\ : LocalMux
    port map (
            O => \N__39281\,
            I => \N__39278\
        );

    \I__8565\ : Span4Mux_h
    port map (
            O => \N__39278\,
            I => \N__39275\
        );

    \I__8564\ : Odrv4
    port map (
            O => \N__39275\,
            I => \delay_measurement_inst.tr_state_RNIMR6LZ0Z_0\
        );

    \I__8563\ : CascadeMux
    port map (
            O => \N__39272\,
            I => \delay_measurement_inst.delay_tr_timer.N_375_cascade_\
        );

    \I__8562\ : CascadeMux
    port map (
            O => \N__39269\,
            I => \delay_measurement_inst.N_265_i_cascade_\
        );

    \I__8561\ : InMux
    port map (
            O => \N__39266\,
            I => \N__39263\
        );

    \I__8560\ : LocalMux
    port map (
            O => \N__39263\,
            I => \N__39260\
        );

    \I__8559\ : Span4Mux_v
    port map (
            O => \N__39260\,
            I => \N__39256\
        );

    \I__8558\ : InMux
    port map (
            O => \N__39259\,
            I => \N__39251\
        );

    \I__8557\ : Span4Mux_v
    port map (
            O => \N__39256\,
            I => \N__39248\
        );

    \I__8556\ : InMux
    port map (
            O => \N__39255\,
            I => \N__39243\
        );

    \I__8555\ : InMux
    port map (
            O => \N__39254\,
            I => \N__39243\
        );

    \I__8554\ : LocalMux
    port map (
            O => \N__39251\,
            I => \N__39240\
        );

    \I__8553\ : Odrv4
    port map (
            O => \N__39248\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__8552\ : LocalMux
    port map (
            O => \N__39243\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__8551\ : Odrv4
    port map (
            O => \N__39240\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__8550\ : CascadeMux
    port map (
            O => \N__39233\,
            I => \N__39228\
        );

    \I__8549\ : CascadeMux
    port map (
            O => \N__39232\,
            I => \N__39225\
        );

    \I__8548\ : InMux
    port map (
            O => \N__39231\,
            I => \N__39222\
        );

    \I__8547\ : InMux
    port map (
            O => \N__39228\,
            I => \N__39217\
        );

    \I__8546\ : InMux
    port map (
            O => \N__39225\,
            I => \N__39217\
        );

    \I__8545\ : LocalMux
    port map (
            O => \N__39222\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__8544\ : LocalMux
    port map (
            O => \N__39217\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__8543\ : InMux
    port map (
            O => \N__39212\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_21\
        );

    \I__8542\ : CascadeMux
    port map (
            O => \N__39209\,
            I => \N__39204\
        );

    \I__8541\ : CascadeMux
    port map (
            O => \N__39208\,
            I => \N__39201\
        );

    \I__8540\ : InMux
    port map (
            O => \N__39207\,
            I => \N__39198\
        );

    \I__8539\ : InMux
    port map (
            O => \N__39204\,
            I => \N__39193\
        );

    \I__8538\ : InMux
    port map (
            O => \N__39201\,
            I => \N__39193\
        );

    \I__8537\ : LocalMux
    port map (
            O => \N__39198\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__8536\ : LocalMux
    port map (
            O => \N__39193\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__8535\ : InMux
    port map (
            O => \N__39188\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_22\
        );

    \I__8534\ : InMux
    port map (
            O => \N__39185\,
            I => \N__39180\
        );

    \I__8533\ : InMux
    port map (
            O => \N__39184\,
            I => \N__39177\
        );

    \I__8532\ : InMux
    port map (
            O => \N__39183\,
            I => \N__39174\
        );

    \I__8531\ : LocalMux
    port map (
            O => \N__39180\,
            I => \N__39171\
        );

    \I__8530\ : LocalMux
    port map (
            O => \N__39177\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__8529\ : LocalMux
    port map (
            O => \N__39174\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__8528\ : Odrv4
    port map (
            O => \N__39171\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__8527\ : InMux
    port map (
            O => \N__39164\,
            I => \bfn_16_10_0_\
        );

    \I__8526\ : InMux
    port map (
            O => \N__39161\,
            I => \N__39156\
        );

    \I__8525\ : InMux
    port map (
            O => \N__39160\,
            I => \N__39153\
        );

    \I__8524\ : InMux
    port map (
            O => \N__39159\,
            I => \N__39150\
        );

    \I__8523\ : LocalMux
    port map (
            O => \N__39156\,
            I => \N__39147\
        );

    \I__8522\ : LocalMux
    port map (
            O => \N__39153\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__8521\ : LocalMux
    port map (
            O => \N__39150\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__8520\ : Odrv4
    port map (
            O => \N__39147\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__8519\ : InMux
    port map (
            O => \N__39140\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_24\
        );

    \I__8518\ : CascadeMux
    port map (
            O => \N__39137\,
            I => \N__39132\
        );

    \I__8517\ : CascadeMux
    port map (
            O => \N__39136\,
            I => \N__39129\
        );

    \I__8516\ : InMux
    port map (
            O => \N__39135\,
            I => \N__39126\
        );

    \I__8515\ : InMux
    port map (
            O => \N__39132\,
            I => \N__39121\
        );

    \I__8514\ : InMux
    port map (
            O => \N__39129\,
            I => \N__39121\
        );

    \I__8513\ : LocalMux
    port map (
            O => \N__39126\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__8512\ : LocalMux
    port map (
            O => \N__39121\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__8511\ : InMux
    port map (
            O => \N__39116\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_25\
        );

    \I__8510\ : CascadeMux
    port map (
            O => \N__39113\,
            I => \N__39108\
        );

    \I__8509\ : CascadeMux
    port map (
            O => \N__39112\,
            I => \N__39105\
        );

    \I__8508\ : InMux
    port map (
            O => \N__39111\,
            I => \N__39102\
        );

    \I__8507\ : InMux
    port map (
            O => \N__39108\,
            I => \N__39097\
        );

    \I__8506\ : InMux
    port map (
            O => \N__39105\,
            I => \N__39097\
        );

    \I__8505\ : LocalMux
    port map (
            O => \N__39102\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__8504\ : LocalMux
    port map (
            O => \N__39097\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__8503\ : InMux
    port map (
            O => \N__39092\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_26\
        );

    \I__8502\ : InMux
    port map (
            O => \N__39089\,
            I => \N__39085\
        );

    \I__8501\ : InMux
    port map (
            O => \N__39088\,
            I => \N__39082\
        );

    \I__8500\ : LocalMux
    port map (
            O => \N__39085\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__8499\ : LocalMux
    port map (
            O => \N__39082\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__8498\ : InMux
    port map (
            O => \N__39077\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_27\
        );

    \I__8497\ : InMux
    port map (
            O => \N__39074\,
            I => \N__39044\
        );

    \I__8496\ : InMux
    port map (
            O => \N__39073\,
            I => \N__39044\
        );

    \I__8495\ : InMux
    port map (
            O => \N__39072\,
            I => \N__39035\
        );

    \I__8494\ : InMux
    port map (
            O => \N__39071\,
            I => \N__39035\
        );

    \I__8493\ : InMux
    port map (
            O => \N__39070\,
            I => \N__39035\
        );

    \I__8492\ : InMux
    port map (
            O => \N__39069\,
            I => \N__39035\
        );

    \I__8491\ : InMux
    port map (
            O => \N__39068\,
            I => \N__39022\
        );

    \I__8490\ : InMux
    port map (
            O => \N__39067\,
            I => \N__39022\
        );

    \I__8489\ : InMux
    port map (
            O => \N__39066\,
            I => \N__39022\
        );

    \I__8488\ : InMux
    port map (
            O => \N__39065\,
            I => \N__39022\
        );

    \I__8487\ : InMux
    port map (
            O => \N__39064\,
            I => \N__39013\
        );

    \I__8486\ : InMux
    port map (
            O => \N__39063\,
            I => \N__39013\
        );

    \I__8485\ : InMux
    port map (
            O => \N__39062\,
            I => \N__39013\
        );

    \I__8484\ : InMux
    port map (
            O => \N__39061\,
            I => \N__39013\
        );

    \I__8483\ : InMux
    port map (
            O => \N__39060\,
            I => \N__39004\
        );

    \I__8482\ : InMux
    port map (
            O => \N__39059\,
            I => \N__39004\
        );

    \I__8481\ : InMux
    port map (
            O => \N__39058\,
            I => \N__39004\
        );

    \I__8480\ : InMux
    port map (
            O => \N__39057\,
            I => \N__39004\
        );

    \I__8479\ : InMux
    port map (
            O => \N__39056\,
            I => \N__38995\
        );

    \I__8478\ : InMux
    port map (
            O => \N__39055\,
            I => \N__38995\
        );

    \I__8477\ : InMux
    port map (
            O => \N__39054\,
            I => \N__38995\
        );

    \I__8476\ : InMux
    port map (
            O => \N__39053\,
            I => \N__38995\
        );

    \I__8475\ : InMux
    port map (
            O => \N__39052\,
            I => \N__38986\
        );

    \I__8474\ : InMux
    port map (
            O => \N__39051\,
            I => \N__38986\
        );

    \I__8473\ : InMux
    port map (
            O => \N__39050\,
            I => \N__38986\
        );

    \I__8472\ : InMux
    port map (
            O => \N__39049\,
            I => \N__38986\
        );

    \I__8471\ : LocalMux
    port map (
            O => \N__39044\,
            I => \N__38983\
        );

    \I__8470\ : LocalMux
    port map (
            O => \N__39035\,
            I => \N__38980\
        );

    \I__8469\ : InMux
    port map (
            O => \N__39034\,
            I => \N__38971\
        );

    \I__8468\ : InMux
    port map (
            O => \N__39033\,
            I => \N__38971\
        );

    \I__8467\ : InMux
    port map (
            O => \N__39032\,
            I => \N__38971\
        );

    \I__8466\ : InMux
    port map (
            O => \N__39031\,
            I => \N__38971\
        );

    \I__8465\ : LocalMux
    port map (
            O => \N__39022\,
            I => \N__38962\
        );

    \I__8464\ : LocalMux
    port map (
            O => \N__39013\,
            I => \N__38962\
        );

    \I__8463\ : LocalMux
    port map (
            O => \N__39004\,
            I => \N__38962\
        );

    \I__8462\ : LocalMux
    port map (
            O => \N__38995\,
            I => \N__38962\
        );

    \I__8461\ : LocalMux
    port map (
            O => \N__38986\,
            I => \N__38959\
        );

    \I__8460\ : Span4Mux_h
    port map (
            O => \N__38983\,
            I => \N__38956\
        );

    \I__8459\ : Span4Mux_h
    port map (
            O => \N__38980\,
            I => \N__38953\
        );

    \I__8458\ : LocalMux
    port map (
            O => \N__38971\,
            I => \N__38948\
        );

    \I__8457\ : Span4Mux_v
    port map (
            O => \N__38962\,
            I => \N__38948\
        );

    \I__8456\ : Odrv12
    port map (
            O => \N__38959\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__8455\ : Odrv4
    port map (
            O => \N__38956\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__8454\ : Odrv4
    port map (
            O => \N__38953\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__8453\ : Odrv4
    port map (
            O => \N__38948\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__8452\ : InMux
    port map (
            O => \N__38939\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_28\
        );

    \I__8451\ : InMux
    port map (
            O => \N__38936\,
            I => \N__38932\
        );

    \I__8450\ : InMux
    port map (
            O => \N__38935\,
            I => \N__38929\
        );

    \I__8449\ : LocalMux
    port map (
            O => \N__38932\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__8448\ : LocalMux
    port map (
            O => \N__38929\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__8447\ : CEMux
    port map (
            O => \N__38924\,
            I => \N__38921\
        );

    \I__8446\ : LocalMux
    port map (
            O => \N__38921\,
            I => \N__38918\
        );

    \I__8445\ : Span4Mux_v
    port map (
            O => \N__38918\,
            I => \N__38913\
        );

    \I__8444\ : CEMux
    port map (
            O => \N__38917\,
            I => \N__38910\
        );

    \I__8443\ : CEMux
    port map (
            O => \N__38916\,
            I => \N__38906\
        );

    \I__8442\ : Span4Mux_h
    port map (
            O => \N__38913\,
            I => \N__38901\
        );

    \I__8441\ : LocalMux
    port map (
            O => \N__38910\,
            I => \N__38901\
        );

    \I__8440\ : CEMux
    port map (
            O => \N__38909\,
            I => \N__38898\
        );

    \I__8439\ : LocalMux
    port map (
            O => \N__38906\,
            I => \N__38895\
        );

    \I__8438\ : Span4Mux_v
    port map (
            O => \N__38901\,
            I => \N__38890\
        );

    \I__8437\ : LocalMux
    port map (
            O => \N__38898\,
            I => \N__38890\
        );

    \I__8436\ : Span4Mux_h
    port map (
            O => \N__38895\,
            I => \N__38887\
        );

    \I__8435\ : Span4Mux_v
    port map (
            O => \N__38890\,
            I => \N__38884\
        );

    \I__8434\ : Odrv4
    port map (
            O => \N__38887\,
            I => \delay_measurement_inst.delay_hc_timer.N_322_i\
        );

    \I__8433\ : Odrv4
    port map (
            O => \N__38884\,
            I => \delay_measurement_inst.delay_hc_timer.N_322_i\
        );

    \I__8432\ : CascadeMux
    port map (
            O => \N__38879\,
            I => \N__38874\
        );

    \I__8431\ : CascadeMux
    port map (
            O => \N__38878\,
            I => \N__38871\
        );

    \I__8430\ : InMux
    port map (
            O => \N__38877\,
            I => \N__38868\
        );

    \I__8429\ : InMux
    port map (
            O => \N__38874\,
            I => \N__38863\
        );

    \I__8428\ : InMux
    port map (
            O => \N__38871\,
            I => \N__38863\
        );

    \I__8427\ : LocalMux
    port map (
            O => \N__38868\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__8426\ : LocalMux
    port map (
            O => \N__38863\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__8425\ : InMux
    port map (
            O => \N__38858\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_13\
        );

    \I__8424\ : CascadeMux
    port map (
            O => \N__38855\,
            I => \N__38850\
        );

    \I__8423\ : CascadeMux
    port map (
            O => \N__38854\,
            I => \N__38847\
        );

    \I__8422\ : InMux
    port map (
            O => \N__38853\,
            I => \N__38844\
        );

    \I__8421\ : InMux
    port map (
            O => \N__38850\,
            I => \N__38839\
        );

    \I__8420\ : InMux
    port map (
            O => \N__38847\,
            I => \N__38839\
        );

    \I__8419\ : LocalMux
    port map (
            O => \N__38844\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__8418\ : LocalMux
    port map (
            O => \N__38839\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__8417\ : InMux
    port map (
            O => \N__38834\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_14\
        );

    \I__8416\ : InMux
    port map (
            O => \N__38831\,
            I => \N__38826\
        );

    \I__8415\ : InMux
    port map (
            O => \N__38830\,
            I => \N__38823\
        );

    \I__8414\ : InMux
    port map (
            O => \N__38829\,
            I => \N__38820\
        );

    \I__8413\ : LocalMux
    port map (
            O => \N__38826\,
            I => \N__38817\
        );

    \I__8412\ : LocalMux
    port map (
            O => \N__38823\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__8411\ : LocalMux
    port map (
            O => \N__38820\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__8410\ : Odrv4
    port map (
            O => \N__38817\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__8409\ : InMux
    port map (
            O => \N__38810\,
            I => \bfn_16_9_0_\
        );

    \I__8408\ : InMux
    port map (
            O => \N__38807\,
            I => \N__38802\
        );

    \I__8407\ : InMux
    port map (
            O => \N__38806\,
            I => \N__38799\
        );

    \I__8406\ : InMux
    port map (
            O => \N__38805\,
            I => \N__38796\
        );

    \I__8405\ : LocalMux
    port map (
            O => \N__38802\,
            I => \N__38793\
        );

    \I__8404\ : LocalMux
    port map (
            O => \N__38799\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__8403\ : LocalMux
    port map (
            O => \N__38796\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__8402\ : Odrv4
    port map (
            O => \N__38793\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__8401\ : InMux
    port map (
            O => \N__38786\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_16\
        );

    \I__8400\ : CascadeMux
    port map (
            O => \N__38783\,
            I => \N__38778\
        );

    \I__8399\ : CascadeMux
    port map (
            O => \N__38782\,
            I => \N__38775\
        );

    \I__8398\ : InMux
    port map (
            O => \N__38781\,
            I => \N__38772\
        );

    \I__8397\ : InMux
    port map (
            O => \N__38778\,
            I => \N__38767\
        );

    \I__8396\ : InMux
    port map (
            O => \N__38775\,
            I => \N__38767\
        );

    \I__8395\ : LocalMux
    port map (
            O => \N__38772\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__8394\ : LocalMux
    port map (
            O => \N__38767\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__8393\ : InMux
    port map (
            O => \N__38762\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_17\
        );

    \I__8392\ : CascadeMux
    port map (
            O => \N__38759\,
            I => \N__38754\
        );

    \I__8391\ : CascadeMux
    port map (
            O => \N__38758\,
            I => \N__38751\
        );

    \I__8390\ : InMux
    port map (
            O => \N__38757\,
            I => \N__38748\
        );

    \I__8389\ : InMux
    port map (
            O => \N__38754\,
            I => \N__38743\
        );

    \I__8388\ : InMux
    port map (
            O => \N__38751\,
            I => \N__38743\
        );

    \I__8387\ : LocalMux
    port map (
            O => \N__38748\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__8386\ : LocalMux
    port map (
            O => \N__38743\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__8385\ : InMux
    port map (
            O => \N__38738\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_18\
        );

    \I__8384\ : InMux
    port map (
            O => \N__38735\,
            I => \N__38730\
        );

    \I__8383\ : InMux
    port map (
            O => \N__38734\,
            I => \N__38725\
        );

    \I__8382\ : InMux
    port map (
            O => \N__38733\,
            I => \N__38725\
        );

    \I__8381\ : LocalMux
    port map (
            O => \N__38730\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__8380\ : LocalMux
    port map (
            O => \N__38725\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__8379\ : InMux
    port map (
            O => \N__38720\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_19\
        );

    \I__8378\ : InMux
    port map (
            O => \N__38717\,
            I => \N__38712\
        );

    \I__8377\ : InMux
    port map (
            O => \N__38716\,
            I => \N__38707\
        );

    \I__8376\ : InMux
    port map (
            O => \N__38715\,
            I => \N__38707\
        );

    \I__8375\ : LocalMux
    port map (
            O => \N__38712\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__8374\ : LocalMux
    port map (
            O => \N__38707\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__8373\ : InMux
    port map (
            O => \N__38702\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_20\
        );

    \I__8372\ : CascadeMux
    port map (
            O => \N__38699\,
            I => \N__38694\
        );

    \I__8371\ : CascadeMux
    port map (
            O => \N__38698\,
            I => \N__38691\
        );

    \I__8370\ : InMux
    port map (
            O => \N__38697\,
            I => \N__38688\
        );

    \I__8369\ : InMux
    port map (
            O => \N__38694\,
            I => \N__38683\
        );

    \I__8368\ : InMux
    port map (
            O => \N__38691\,
            I => \N__38683\
        );

    \I__8367\ : LocalMux
    port map (
            O => \N__38688\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__8366\ : LocalMux
    port map (
            O => \N__38683\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__8365\ : InMux
    port map (
            O => \N__38678\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_5\
        );

    \I__8364\ : CascadeMux
    port map (
            O => \N__38675\,
            I => \N__38670\
        );

    \I__8363\ : CascadeMux
    port map (
            O => \N__38674\,
            I => \N__38667\
        );

    \I__8362\ : InMux
    port map (
            O => \N__38673\,
            I => \N__38664\
        );

    \I__8361\ : InMux
    port map (
            O => \N__38670\,
            I => \N__38659\
        );

    \I__8360\ : InMux
    port map (
            O => \N__38667\,
            I => \N__38659\
        );

    \I__8359\ : LocalMux
    port map (
            O => \N__38664\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__8358\ : LocalMux
    port map (
            O => \N__38659\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__8357\ : InMux
    port map (
            O => \N__38654\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_6\
        );

    \I__8356\ : InMux
    port map (
            O => \N__38651\,
            I => \N__38646\
        );

    \I__8355\ : InMux
    port map (
            O => \N__38650\,
            I => \N__38643\
        );

    \I__8354\ : InMux
    port map (
            O => \N__38649\,
            I => \N__38640\
        );

    \I__8353\ : LocalMux
    port map (
            O => \N__38646\,
            I => \N__38637\
        );

    \I__8352\ : LocalMux
    port map (
            O => \N__38643\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__8351\ : LocalMux
    port map (
            O => \N__38640\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__8350\ : Odrv4
    port map (
            O => \N__38637\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__8349\ : InMux
    port map (
            O => \N__38630\,
            I => \bfn_16_8_0_\
        );

    \I__8348\ : InMux
    port map (
            O => \N__38627\,
            I => \N__38622\
        );

    \I__8347\ : InMux
    port map (
            O => \N__38626\,
            I => \N__38619\
        );

    \I__8346\ : InMux
    port map (
            O => \N__38625\,
            I => \N__38616\
        );

    \I__8345\ : LocalMux
    port map (
            O => \N__38622\,
            I => \N__38613\
        );

    \I__8344\ : LocalMux
    port map (
            O => \N__38619\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__8343\ : LocalMux
    port map (
            O => \N__38616\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__8342\ : Odrv4
    port map (
            O => \N__38613\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__8341\ : InMux
    port map (
            O => \N__38606\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_8\
        );

    \I__8340\ : CascadeMux
    port map (
            O => \N__38603\,
            I => \N__38598\
        );

    \I__8339\ : CascadeMux
    port map (
            O => \N__38602\,
            I => \N__38595\
        );

    \I__8338\ : InMux
    port map (
            O => \N__38601\,
            I => \N__38592\
        );

    \I__8337\ : InMux
    port map (
            O => \N__38598\,
            I => \N__38587\
        );

    \I__8336\ : InMux
    port map (
            O => \N__38595\,
            I => \N__38587\
        );

    \I__8335\ : LocalMux
    port map (
            O => \N__38592\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__8334\ : LocalMux
    port map (
            O => \N__38587\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__8333\ : InMux
    port map (
            O => \N__38582\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_9\
        );

    \I__8332\ : CascadeMux
    port map (
            O => \N__38579\,
            I => \N__38574\
        );

    \I__8331\ : CascadeMux
    port map (
            O => \N__38578\,
            I => \N__38571\
        );

    \I__8330\ : InMux
    port map (
            O => \N__38577\,
            I => \N__38568\
        );

    \I__8329\ : InMux
    port map (
            O => \N__38574\,
            I => \N__38563\
        );

    \I__8328\ : InMux
    port map (
            O => \N__38571\,
            I => \N__38563\
        );

    \I__8327\ : LocalMux
    port map (
            O => \N__38568\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__8326\ : LocalMux
    port map (
            O => \N__38563\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__8325\ : InMux
    port map (
            O => \N__38558\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_10\
        );

    \I__8324\ : InMux
    port map (
            O => \N__38555\,
            I => \N__38550\
        );

    \I__8323\ : InMux
    port map (
            O => \N__38554\,
            I => \N__38545\
        );

    \I__8322\ : InMux
    port map (
            O => \N__38553\,
            I => \N__38545\
        );

    \I__8321\ : LocalMux
    port map (
            O => \N__38550\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__8320\ : LocalMux
    port map (
            O => \N__38545\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__8319\ : InMux
    port map (
            O => \N__38540\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_11\
        );

    \I__8318\ : InMux
    port map (
            O => \N__38537\,
            I => \N__38532\
        );

    \I__8317\ : InMux
    port map (
            O => \N__38536\,
            I => \N__38527\
        );

    \I__8316\ : InMux
    port map (
            O => \N__38535\,
            I => \N__38527\
        );

    \I__8315\ : LocalMux
    port map (
            O => \N__38532\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__8314\ : LocalMux
    port map (
            O => \N__38527\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__8313\ : InMux
    port map (
            O => \N__38522\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_12\
        );

    \I__8312\ : InMux
    port map (
            O => \N__38519\,
            I => \N__38516\
        );

    \I__8311\ : LocalMux
    port map (
            O => \N__38516\,
            I => \N__38513\
        );

    \I__8310\ : Odrv4
    port map (
            O => \N__38513\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9\
        );

    \I__8309\ : InMux
    port map (
            O => \N__38510\,
            I => \N__38506\
        );

    \I__8308\ : InMux
    port map (
            O => \N__38509\,
            I => \N__38503\
        );

    \I__8307\ : LocalMux
    port map (
            O => \N__38506\,
            I => \N__38500\
        );

    \I__8306\ : LocalMux
    port map (
            O => \N__38503\,
            I => \N__38497\
        );

    \I__8305\ : Span4Mux_v
    port map (
            O => \N__38500\,
            I => \N__38494\
        );

    \I__8304\ : Odrv4
    port map (
            O => \N__38497\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__8303\ : Odrv4
    port map (
            O => \N__38494\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__8302\ : CascadeMux
    port map (
            O => \N__38489\,
            I => \N__38486\
        );

    \I__8301\ : InMux
    port map (
            O => \N__38486\,
            I => \N__38483\
        );

    \I__8300\ : LocalMux
    port map (
            O => \N__38483\,
            I => \N__38480\
        );

    \I__8299\ : Odrv12
    port map (
            O => \N__38480\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15\
        );

    \I__8298\ : InMux
    port map (
            O => \N__38477\,
            I => \N__38473\
        );

    \I__8297\ : InMux
    port map (
            O => \N__38476\,
            I => \N__38470\
        );

    \I__8296\ : LocalMux
    port map (
            O => \N__38473\,
            I => \N__38467\
        );

    \I__8295\ : LocalMux
    port map (
            O => \N__38470\,
            I => \N__38464\
        );

    \I__8294\ : Span4Mux_v
    port map (
            O => \N__38467\,
            I => \N__38461\
        );

    \I__8293\ : Odrv12
    port map (
            O => \N__38464\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__8292\ : Odrv4
    port map (
            O => \N__38461\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__8291\ : InMux
    port map (
            O => \N__38456\,
            I => \N__38451\
        );

    \I__8290\ : InMux
    port map (
            O => \N__38455\,
            I => \N__38448\
        );

    \I__8289\ : InMux
    port map (
            O => \N__38454\,
            I => \N__38445\
        );

    \I__8288\ : LocalMux
    port map (
            O => \N__38451\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__8287\ : LocalMux
    port map (
            O => \N__38448\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__8286\ : LocalMux
    port map (
            O => \N__38445\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__8285\ : InMux
    port map (
            O => \N__38438\,
            I => \bfn_16_7_0_\
        );

    \I__8284\ : InMux
    port map (
            O => \N__38435\,
            I => \N__38430\
        );

    \I__8283\ : InMux
    port map (
            O => \N__38434\,
            I => \N__38427\
        );

    \I__8282\ : InMux
    port map (
            O => \N__38433\,
            I => \N__38424\
        );

    \I__8281\ : LocalMux
    port map (
            O => \N__38430\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__8280\ : LocalMux
    port map (
            O => \N__38427\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__38424\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__8278\ : InMux
    port map (
            O => \N__38417\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_0\
        );

    \I__8277\ : CascadeMux
    port map (
            O => \N__38414\,
            I => \N__38409\
        );

    \I__8276\ : CascadeMux
    port map (
            O => \N__38413\,
            I => \N__38406\
        );

    \I__8275\ : InMux
    port map (
            O => \N__38412\,
            I => \N__38403\
        );

    \I__8274\ : InMux
    port map (
            O => \N__38409\,
            I => \N__38398\
        );

    \I__8273\ : InMux
    port map (
            O => \N__38406\,
            I => \N__38398\
        );

    \I__8272\ : LocalMux
    port map (
            O => \N__38403\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__8271\ : LocalMux
    port map (
            O => \N__38398\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__8270\ : InMux
    port map (
            O => \N__38393\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_1\
        );

    \I__8269\ : CascadeMux
    port map (
            O => \N__38390\,
            I => \N__38385\
        );

    \I__8268\ : CascadeMux
    port map (
            O => \N__38389\,
            I => \N__38382\
        );

    \I__8267\ : InMux
    port map (
            O => \N__38388\,
            I => \N__38379\
        );

    \I__8266\ : InMux
    port map (
            O => \N__38385\,
            I => \N__38374\
        );

    \I__8265\ : InMux
    port map (
            O => \N__38382\,
            I => \N__38374\
        );

    \I__8264\ : LocalMux
    port map (
            O => \N__38379\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__8263\ : LocalMux
    port map (
            O => \N__38374\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__8262\ : InMux
    port map (
            O => \N__38369\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_2\
        );

    \I__8261\ : InMux
    port map (
            O => \N__38366\,
            I => \N__38361\
        );

    \I__8260\ : InMux
    port map (
            O => \N__38365\,
            I => \N__38356\
        );

    \I__8259\ : InMux
    port map (
            O => \N__38364\,
            I => \N__38356\
        );

    \I__8258\ : LocalMux
    port map (
            O => \N__38361\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__8257\ : LocalMux
    port map (
            O => \N__38356\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__8256\ : InMux
    port map (
            O => \N__38351\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_3\
        );

    \I__8255\ : InMux
    port map (
            O => \N__38348\,
            I => \N__38343\
        );

    \I__8254\ : InMux
    port map (
            O => \N__38347\,
            I => \N__38338\
        );

    \I__8253\ : InMux
    port map (
            O => \N__38346\,
            I => \N__38338\
        );

    \I__8252\ : LocalMux
    port map (
            O => \N__38343\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__8251\ : LocalMux
    port map (
            O => \N__38338\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__8250\ : InMux
    port map (
            O => \N__38333\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_4\
        );

    \I__8249\ : InMux
    port map (
            O => \N__38330\,
            I => \N__38327\
        );

    \I__8248\ : LocalMux
    port map (
            O => \N__38327\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14\
        );

    \I__8247\ : InMux
    port map (
            O => \N__38324\,
            I => \N__38321\
        );

    \I__8246\ : LocalMux
    port map (
            O => \N__38321\,
            I => \N__38317\
        );

    \I__8245\ : InMux
    port map (
            O => \N__38320\,
            I => \N__38314\
        );

    \I__8244\ : Span4Mux_h
    port map (
            O => \N__38317\,
            I => \N__38311\
        );

    \I__8243\ : LocalMux
    port map (
            O => \N__38314\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__8242\ : Odrv4
    port map (
            O => \N__38311\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__8241\ : CascadeMux
    port map (
            O => \N__38306\,
            I => \N__38303\
        );

    \I__8240\ : InMux
    port map (
            O => \N__38303\,
            I => \N__38300\
        );

    \I__8239\ : LocalMux
    port map (
            O => \N__38300\,
            I => \N__38297\
        );

    \I__8238\ : Span4Mux_v
    port map (
            O => \N__38297\,
            I => \N__38294\
        );

    \I__8237\ : Odrv4
    port map (
            O => \N__38294\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0\
        );

    \I__8236\ : CascadeMux
    port map (
            O => \N__38291\,
            I => \N__38288\
        );

    \I__8235\ : InMux
    port map (
            O => \N__38288\,
            I => \N__38283\
        );

    \I__8234\ : InMux
    port map (
            O => \N__38287\,
            I => \N__38280\
        );

    \I__8233\ : InMux
    port map (
            O => \N__38286\,
            I => \N__38277\
        );

    \I__8232\ : LocalMux
    port map (
            O => \N__38283\,
            I => \N__38274\
        );

    \I__8231\ : LocalMux
    port map (
            O => \N__38280\,
            I => \N__38269\
        );

    \I__8230\ : LocalMux
    port map (
            O => \N__38277\,
            I => \N__38269\
        );

    \I__8229\ : Odrv4
    port map (
            O => \N__38274\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__8228\ : Odrv12
    port map (
            O => \N__38269\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__8227\ : InMux
    port map (
            O => \N__38264\,
            I => \N__38261\
        );

    \I__8226\ : LocalMux
    port map (
            O => \N__38261\,
            I => \N__38258\
        );

    \I__8225\ : Span4Mux_h
    port map (
            O => \N__38258\,
            I => \N__38255\
        );

    \I__8224\ : Odrv4
    port map (
            O => \N__38255\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2\
        );

    \I__8223\ : InMux
    port map (
            O => \N__38252\,
            I => \N__38248\
        );

    \I__8222\ : InMux
    port map (
            O => \N__38251\,
            I => \N__38245\
        );

    \I__8221\ : LocalMux
    port map (
            O => \N__38248\,
            I => \N__38242\
        );

    \I__8220\ : LocalMux
    port map (
            O => \N__38245\,
            I => \N__38239\
        );

    \I__8219\ : Odrv4
    port map (
            O => \N__38242\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__8218\ : Odrv12
    port map (
            O => \N__38239\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__8217\ : CascadeMux
    port map (
            O => \N__38234\,
            I => \N__38231\
        );

    \I__8216\ : InMux
    port map (
            O => \N__38231\,
            I => \N__38228\
        );

    \I__8215\ : LocalMux
    port map (
            O => \N__38228\,
            I => \N__38225\
        );

    \I__8214\ : Odrv4
    port map (
            O => \N__38225\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17\
        );

    \I__8213\ : InMux
    port map (
            O => \N__38222\,
            I => \N__38219\
        );

    \I__8212\ : LocalMux
    port map (
            O => \N__38219\,
            I => \N__38215\
        );

    \I__8211\ : InMux
    port map (
            O => \N__38218\,
            I => \N__38212\
        );

    \I__8210\ : Span4Mux_h
    port map (
            O => \N__38215\,
            I => \N__38209\
        );

    \I__8209\ : LocalMux
    port map (
            O => \N__38212\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__8208\ : Odrv4
    port map (
            O => \N__38209\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__8207\ : InMux
    port map (
            O => \N__38204\,
            I => \N__38201\
        );

    \I__8206\ : LocalMux
    port map (
            O => \N__38201\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18\
        );

    \I__8205\ : InMux
    port map (
            O => \N__38198\,
            I => \N__38195\
        );

    \I__8204\ : LocalMux
    port map (
            O => \N__38195\,
            I => \N__38191\
        );

    \I__8203\ : InMux
    port map (
            O => \N__38194\,
            I => \N__38188\
        );

    \I__8202\ : Span4Mux_h
    port map (
            O => \N__38191\,
            I => \N__38185\
        );

    \I__8201\ : LocalMux
    port map (
            O => \N__38188\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__8200\ : Odrv4
    port map (
            O => \N__38185\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__8199\ : CascadeMux
    port map (
            O => \N__38180\,
            I => \N__38170\
        );

    \I__8198\ : CascadeMux
    port map (
            O => \N__38179\,
            I => \N__38167\
        );

    \I__8197\ : InMux
    port map (
            O => \N__38178\,
            I => \N__38148\
        );

    \I__8196\ : InMux
    port map (
            O => \N__38177\,
            I => \N__38148\
        );

    \I__8195\ : InMux
    port map (
            O => \N__38176\,
            I => \N__38148\
        );

    \I__8194\ : InMux
    port map (
            O => \N__38175\,
            I => \N__38148\
        );

    \I__8193\ : InMux
    port map (
            O => \N__38174\,
            I => \N__38148\
        );

    \I__8192\ : InMux
    port map (
            O => \N__38173\,
            I => \N__38127\
        );

    \I__8191\ : InMux
    port map (
            O => \N__38170\,
            I => \N__38127\
        );

    \I__8190\ : InMux
    port map (
            O => \N__38167\,
            I => \N__38127\
        );

    \I__8189\ : InMux
    port map (
            O => \N__38166\,
            I => \N__38127\
        );

    \I__8188\ : InMux
    port map (
            O => \N__38165\,
            I => \N__38127\
        );

    \I__8187\ : InMux
    port map (
            O => \N__38164\,
            I => \N__38127\
        );

    \I__8186\ : InMux
    port map (
            O => \N__38163\,
            I => \N__38127\
        );

    \I__8185\ : InMux
    port map (
            O => \N__38162\,
            I => \N__38118\
        );

    \I__8184\ : InMux
    port map (
            O => \N__38161\,
            I => \N__38118\
        );

    \I__8183\ : InMux
    port map (
            O => \N__38160\,
            I => \N__38118\
        );

    \I__8182\ : InMux
    port map (
            O => \N__38159\,
            I => \N__38118\
        );

    \I__8181\ : LocalMux
    port map (
            O => \N__38148\,
            I => \N__38114\
        );

    \I__8180\ : InMux
    port map (
            O => \N__38147\,
            I => \N__38107\
        );

    \I__8179\ : InMux
    port map (
            O => \N__38146\,
            I => \N__38107\
        );

    \I__8178\ : InMux
    port map (
            O => \N__38145\,
            I => \N__38107\
        );

    \I__8177\ : CascadeMux
    port map (
            O => \N__38144\,
            I => \N__38104\
        );

    \I__8176\ : InMux
    port map (
            O => \N__38143\,
            I => \N__38098\
        );

    \I__8175\ : InMux
    port map (
            O => \N__38142\,
            I => \N__38098\
        );

    \I__8174\ : LocalMux
    port map (
            O => \N__38127\,
            I => \N__38093\
        );

    \I__8173\ : LocalMux
    port map (
            O => \N__38118\,
            I => \N__38093\
        );

    \I__8172\ : InMux
    port map (
            O => \N__38117\,
            I => \N__38090\
        );

    \I__8171\ : Span4Mux_h
    port map (
            O => \N__38114\,
            I => \N__38085\
        );

    \I__8170\ : LocalMux
    port map (
            O => \N__38107\,
            I => \N__38085\
        );

    \I__8169\ : InMux
    port map (
            O => \N__38104\,
            I => \N__38080\
        );

    \I__8168\ : InMux
    port map (
            O => \N__38103\,
            I => \N__38080\
        );

    \I__8167\ : LocalMux
    port map (
            O => \N__38098\,
            I => \N__38075\
        );

    \I__8166\ : Span4Mux_v
    port map (
            O => \N__38093\,
            I => \N__38075\
        );

    \I__8165\ : LocalMux
    port map (
            O => \N__38090\,
            I => \N__38072\
        );

    \I__8164\ : Span4Mux_v
    port map (
            O => \N__38085\,
            I => \N__38069\
        );

    \I__8163\ : LocalMux
    port map (
            O => \N__38080\,
            I => \N__38064\
        );

    \I__8162\ : Span4Mux_v
    port map (
            O => \N__38075\,
            I => \N__38064\
        );

    \I__8161\ : Span4Mux_h
    port map (
            O => \N__38072\,
            I => \N__38061\
        );

    \I__8160\ : Span4Mux_v
    port map (
            O => \N__38069\,
            I => \N__38058\
        );

    \I__8159\ : Odrv4
    port map (
            O => \N__38064\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__8158\ : Odrv4
    port map (
            O => \N__38061\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__8157\ : Odrv4
    port map (
            O => \N__38058\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__8156\ : CascadeMux
    port map (
            O => \N__38051\,
            I => \N__38040\
        );

    \I__8155\ : CascadeMux
    port map (
            O => \N__38050\,
            I => \N__38034\
        );

    \I__8154\ : CascadeMux
    port map (
            O => \N__38049\,
            I => \N__38031\
        );

    \I__8153\ : CascadeMux
    port map (
            O => \N__38048\,
            I => \N__38028\
        );

    \I__8152\ : CascadeMux
    port map (
            O => \N__38047\,
            I => \N__38025\
        );

    \I__8151\ : CascadeMux
    port map (
            O => \N__38046\,
            I => \N__38019\
        );

    \I__8150\ : InMux
    port map (
            O => \N__38045\,
            I => \N__38012\
        );

    \I__8149\ : CascadeMux
    port map (
            O => \N__38044\,
            I => \N__38009\
        );

    \I__8148\ : CascadeMux
    port map (
            O => \N__38043\,
            I => \N__38006\
        );

    \I__8147\ : InMux
    port map (
            O => \N__38040\,
            I => \N__37999\
        );

    \I__8146\ : InMux
    port map (
            O => \N__38039\,
            I => \N__37999\
        );

    \I__8145\ : InMux
    port map (
            O => \N__38038\,
            I => \N__37987\
        );

    \I__8144\ : InMux
    port map (
            O => \N__38037\,
            I => \N__37987\
        );

    \I__8143\ : InMux
    port map (
            O => \N__38034\,
            I => \N__37987\
        );

    \I__8142\ : InMux
    port map (
            O => \N__38031\,
            I => \N__37987\
        );

    \I__8141\ : InMux
    port map (
            O => \N__38028\,
            I => \N__37987\
        );

    \I__8140\ : InMux
    port map (
            O => \N__38025\,
            I => \N__37982\
        );

    \I__8139\ : InMux
    port map (
            O => \N__38024\,
            I => \N__37982\
        );

    \I__8138\ : InMux
    port map (
            O => \N__38023\,
            I => \N__37967\
        );

    \I__8137\ : InMux
    port map (
            O => \N__38022\,
            I => \N__37967\
        );

    \I__8136\ : InMux
    port map (
            O => \N__38019\,
            I => \N__37967\
        );

    \I__8135\ : InMux
    port map (
            O => \N__38018\,
            I => \N__37967\
        );

    \I__8134\ : InMux
    port map (
            O => \N__38017\,
            I => \N__37967\
        );

    \I__8133\ : InMux
    port map (
            O => \N__38016\,
            I => \N__37967\
        );

    \I__8132\ : InMux
    port map (
            O => \N__38015\,
            I => \N__37967\
        );

    \I__8131\ : LocalMux
    port map (
            O => \N__38012\,
            I => \N__37964\
        );

    \I__8130\ : InMux
    port map (
            O => \N__38009\,
            I => \N__37955\
        );

    \I__8129\ : InMux
    port map (
            O => \N__38006\,
            I => \N__37955\
        );

    \I__8128\ : InMux
    port map (
            O => \N__38005\,
            I => \N__37955\
        );

    \I__8127\ : InMux
    port map (
            O => \N__38004\,
            I => \N__37955\
        );

    \I__8126\ : LocalMux
    port map (
            O => \N__37999\,
            I => \N__37952\
        );

    \I__8125\ : CascadeMux
    port map (
            O => \N__37998\,
            I => \N__37948\
        );

    \I__8124\ : LocalMux
    port map (
            O => \N__37987\,
            I => \N__37944\
        );

    \I__8123\ : LocalMux
    port map (
            O => \N__37982\,
            I => \N__37937\
        );

    \I__8122\ : LocalMux
    port map (
            O => \N__37967\,
            I => \N__37937\
        );

    \I__8121\ : Span4Mux_v
    port map (
            O => \N__37964\,
            I => \N__37937\
        );

    \I__8120\ : LocalMux
    port map (
            O => \N__37955\,
            I => \N__37934\
        );

    \I__8119\ : Sp12to4
    port map (
            O => \N__37952\,
            I => \N__37931\
        );

    \I__8118\ : InMux
    port map (
            O => \N__37951\,
            I => \N__37924\
        );

    \I__8117\ : InMux
    port map (
            O => \N__37948\,
            I => \N__37924\
        );

    \I__8116\ : InMux
    port map (
            O => \N__37947\,
            I => \N__37924\
        );

    \I__8115\ : Span4Mux_h
    port map (
            O => \N__37944\,
            I => \N__37919\
        );

    \I__8114\ : Span4Mux_v
    port map (
            O => \N__37937\,
            I => \N__37919\
        );

    \I__8113\ : Odrv4
    port map (
            O => \N__37934\,
            I => \phase_controller_slave.start_timer_trZ0\
        );

    \I__8112\ : Odrv12
    port map (
            O => \N__37931\,
            I => \phase_controller_slave.start_timer_trZ0\
        );

    \I__8111\ : LocalMux
    port map (
            O => \N__37924\,
            I => \phase_controller_slave.start_timer_trZ0\
        );

    \I__8110\ : Odrv4
    port map (
            O => \N__37919\,
            I => \phase_controller_slave.start_timer_trZ0\
        );

    \I__8109\ : CascadeMux
    port map (
            O => \N__37910\,
            I => \N__37907\
        );

    \I__8108\ : InMux
    port map (
            O => \N__37907\,
            I => \N__37904\
        );

    \I__8107\ : LocalMux
    port map (
            O => \N__37904\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19\
        );

    \I__8106\ : CascadeMux
    port map (
            O => \N__37901\,
            I => \N__37889\
        );

    \I__8105\ : CascadeMux
    port map (
            O => \N__37900\,
            I => \N__37886\
        );

    \I__8104\ : CascadeMux
    port map (
            O => \N__37899\,
            I => \N__37881\
        );

    \I__8103\ : CascadeMux
    port map (
            O => \N__37898\,
            I => \N__37878\
        );

    \I__8102\ : InMux
    port map (
            O => \N__37897\,
            I => \N__37862\
        );

    \I__8101\ : InMux
    port map (
            O => \N__37896\,
            I => \N__37862\
        );

    \I__8100\ : InMux
    port map (
            O => \N__37895\,
            I => \N__37862\
        );

    \I__8099\ : InMux
    port map (
            O => \N__37894\,
            I => \N__37862\
        );

    \I__8098\ : InMux
    port map (
            O => \N__37893\,
            I => \N__37862\
        );

    \I__8097\ : InMux
    port map (
            O => \N__37892\,
            I => \N__37855\
        );

    \I__8096\ : InMux
    port map (
            O => \N__37889\,
            I => \N__37850\
        );

    \I__8095\ : InMux
    port map (
            O => \N__37886\,
            I => \N__37850\
        );

    \I__8094\ : InMux
    port map (
            O => \N__37885\,
            I => \N__37845\
        );

    \I__8093\ : InMux
    port map (
            O => \N__37884\,
            I => \N__37845\
        );

    \I__8092\ : InMux
    port map (
            O => \N__37881\,
            I => \N__37830\
        );

    \I__8091\ : InMux
    port map (
            O => \N__37878\,
            I => \N__37830\
        );

    \I__8090\ : InMux
    port map (
            O => \N__37877\,
            I => \N__37830\
        );

    \I__8089\ : InMux
    port map (
            O => \N__37876\,
            I => \N__37830\
        );

    \I__8088\ : InMux
    port map (
            O => \N__37875\,
            I => \N__37830\
        );

    \I__8087\ : InMux
    port map (
            O => \N__37874\,
            I => \N__37830\
        );

    \I__8086\ : InMux
    port map (
            O => \N__37873\,
            I => \N__37830\
        );

    \I__8085\ : LocalMux
    port map (
            O => \N__37862\,
            I => \N__37827\
        );

    \I__8084\ : InMux
    port map (
            O => \N__37861\,
            I => \N__37823\
        );

    \I__8083\ : InMux
    port map (
            O => \N__37860\,
            I => \N__37818\
        );

    \I__8082\ : InMux
    port map (
            O => \N__37859\,
            I => \N__37818\
        );

    \I__8081\ : InMux
    port map (
            O => \N__37858\,
            I => \N__37815\
        );

    \I__8080\ : LocalMux
    port map (
            O => \N__37855\,
            I => \N__37812\
        );

    \I__8079\ : LocalMux
    port map (
            O => \N__37850\,
            I => \N__37803\
        );

    \I__8078\ : LocalMux
    port map (
            O => \N__37845\,
            I => \N__37803\
        );

    \I__8077\ : LocalMux
    port map (
            O => \N__37830\,
            I => \N__37803\
        );

    \I__8076\ : Span4Mux_v
    port map (
            O => \N__37827\,
            I => \N__37803\
        );

    \I__8075\ : InMux
    port map (
            O => \N__37826\,
            I => \N__37800\
        );

    \I__8074\ : LocalMux
    port map (
            O => \N__37823\,
            I => \N__37795\
        );

    \I__8073\ : LocalMux
    port map (
            O => \N__37818\,
            I => \N__37795\
        );

    \I__8072\ : LocalMux
    port map (
            O => \N__37815\,
            I => \N__37786\
        );

    \I__8071\ : Span4Mux_h
    port map (
            O => \N__37812\,
            I => \N__37786\
        );

    \I__8070\ : Span4Mux_v
    port map (
            O => \N__37803\,
            I => \N__37786\
        );

    \I__8069\ : LocalMux
    port map (
            O => \N__37800\,
            I => \N__37783\
        );

    \I__8068\ : Span4Mux_v
    port map (
            O => \N__37795\,
            I => \N__37780\
        );

    \I__8067\ : InMux
    port map (
            O => \N__37794\,
            I => \N__37775\
        );

    \I__8066\ : InMux
    port map (
            O => \N__37793\,
            I => \N__37775\
        );

    \I__8065\ : Span4Mux_v
    port map (
            O => \N__37786\,
            I => \N__37770\
        );

    \I__8064\ : Span4Mux_v
    port map (
            O => \N__37783\,
            I => \N__37770\
        );

    \I__8063\ : Span4Mux_v
    port map (
            O => \N__37780\,
            I => \N__37767\
        );

    \I__8062\ : LocalMux
    port map (
            O => \N__37775\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__8061\ : Odrv4
    port map (
            O => \N__37770\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__8060\ : Odrv4
    port map (
            O => \N__37767\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__8059\ : InMux
    port map (
            O => \N__37760\,
            I => \N__37757\
        );

    \I__8058\ : LocalMux
    port map (
            O => \N__37757\,
            I => \N__37753\
        );

    \I__8057\ : InMux
    port map (
            O => \N__37756\,
            I => \N__37750\
        );

    \I__8056\ : Span4Mux_h
    port map (
            O => \N__37753\,
            I => \N__37747\
        );

    \I__8055\ : LocalMux
    port map (
            O => \N__37750\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__8054\ : Odrv4
    port map (
            O => \N__37747\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__8053\ : InMux
    port map (
            O => \N__37742\,
            I => \N__37739\
        );

    \I__8052\ : LocalMux
    port map (
            O => \N__37739\,
            I => \N__37736\
        );

    \I__8051\ : Odrv4
    port map (
            O => \N__37736\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10\
        );

    \I__8050\ : InMux
    port map (
            O => \N__37733\,
            I => \N__37729\
        );

    \I__8049\ : InMux
    port map (
            O => \N__37732\,
            I => \N__37726\
        );

    \I__8048\ : LocalMux
    port map (
            O => \N__37729\,
            I => \N__37723\
        );

    \I__8047\ : LocalMux
    port map (
            O => \N__37726\,
            I => \N__37720\
        );

    \I__8046\ : Odrv12
    port map (
            O => \N__37723\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__8045\ : Odrv12
    port map (
            O => \N__37720\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__8044\ : InMux
    port map (
            O => \N__37715\,
            I => \N__37712\
        );

    \I__8043\ : LocalMux
    port map (
            O => \N__37712\,
            I => \N__37709\
        );

    \I__8042\ : Odrv4
    port map (
            O => \N__37709\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11\
        );

    \I__8041\ : InMux
    port map (
            O => \N__37706\,
            I => \N__37702\
        );

    \I__8040\ : InMux
    port map (
            O => \N__37705\,
            I => \N__37699\
        );

    \I__8039\ : LocalMux
    port map (
            O => \N__37702\,
            I => \N__37696\
        );

    \I__8038\ : LocalMux
    port map (
            O => \N__37699\,
            I => \N__37693\
        );

    \I__8037\ : Span4Mux_v
    port map (
            O => \N__37696\,
            I => \N__37690\
        );

    \I__8036\ : Odrv4
    port map (
            O => \N__37693\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__8035\ : Odrv4
    port map (
            O => \N__37690\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__8034\ : InMux
    port map (
            O => \N__37685\,
            I => \N__37682\
        );

    \I__8033\ : LocalMux
    port map (
            O => \N__37682\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15\
        );

    \I__8032\ : InMux
    port map (
            O => \N__37679\,
            I => \N__37676\
        );

    \I__8031\ : LocalMux
    port map (
            O => \N__37676\,
            I => \N__37672\
        );

    \I__8030\ : InMux
    port map (
            O => \N__37675\,
            I => \N__37669\
        );

    \I__8029\ : Span4Mux_h
    port map (
            O => \N__37672\,
            I => \N__37666\
        );

    \I__8028\ : LocalMux
    port map (
            O => \N__37669\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__8027\ : Odrv4
    port map (
            O => \N__37666\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__8026\ : InMux
    port map (
            O => \N__37661\,
            I => \N__37658\
        );

    \I__8025\ : LocalMux
    port map (
            O => \N__37658\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12\
        );

    \I__8024\ : InMux
    port map (
            O => \N__37655\,
            I => \N__37652\
        );

    \I__8023\ : LocalMux
    port map (
            O => \N__37652\,
            I => \N__37648\
        );

    \I__8022\ : InMux
    port map (
            O => \N__37651\,
            I => \N__37645\
        );

    \I__8021\ : Span4Mux_v
    port map (
            O => \N__37648\,
            I => \N__37642\
        );

    \I__8020\ : LocalMux
    port map (
            O => \N__37645\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__8019\ : Odrv4
    port map (
            O => \N__37642\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__8018\ : InMux
    port map (
            O => \N__37637\,
            I => \N__37634\
        );

    \I__8017\ : LocalMux
    port map (
            O => \N__37634\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16\
        );

    \I__8016\ : InMux
    port map (
            O => \N__37631\,
            I => \N__37628\
        );

    \I__8015\ : LocalMux
    port map (
            O => \N__37628\,
            I => \N__37624\
        );

    \I__8014\ : InMux
    port map (
            O => \N__37627\,
            I => \N__37621\
        );

    \I__8013\ : Span4Mux_v
    port map (
            O => \N__37624\,
            I => \N__37618\
        );

    \I__8012\ : LocalMux
    port map (
            O => \N__37621\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__8011\ : Odrv4
    port map (
            O => \N__37618\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__8010\ : InMux
    port map (
            O => \N__37613\,
            I => \N__37610\
        );

    \I__8009\ : LocalMux
    port map (
            O => \N__37610\,
            I => \N__37607\
        );

    \I__8008\ : Span4Mux_h
    port map (
            O => \N__37607\,
            I => \N__37604\
        );

    \I__8007\ : Odrv4
    port map (
            O => \N__37604\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4\
        );

    \I__8006\ : InMux
    port map (
            O => \N__37601\,
            I => \N__37598\
        );

    \I__8005\ : LocalMux
    port map (
            O => \N__37598\,
            I => \N__37594\
        );

    \I__8004\ : InMux
    port map (
            O => \N__37597\,
            I => \N__37591\
        );

    \I__8003\ : Span4Mux_v
    port map (
            O => \N__37594\,
            I => \N__37588\
        );

    \I__8002\ : LocalMux
    port map (
            O => \N__37591\,
            I => \N__37585\
        );

    \I__8001\ : Odrv4
    port map (
            O => \N__37588\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__8000\ : Odrv12
    port map (
            O => \N__37585\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__7999\ : InMux
    port map (
            O => \N__37580\,
            I => \N__37577\
        );

    \I__7998\ : LocalMux
    port map (
            O => \N__37577\,
            I => \N__37574\
        );

    \I__7997\ : Span4Mux_h
    port map (
            O => \N__37574\,
            I => \N__37571\
        );

    \I__7996\ : Odrv4
    port map (
            O => \N__37571\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5\
        );

    \I__7995\ : InMux
    port map (
            O => \N__37568\,
            I => \N__37565\
        );

    \I__7994\ : LocalMux
    port map (
            O => \N__37565\,
            I => \N__37561\
        );

    \I__7993\ : InMux
    port map (
            O => \N__37564\,
            I => \N__37558\
        );

    \I__7992\ : Span4Mux_h
    port map (
            O => \N__37561\,
            I => \N__37555\
        );

    \I__7991\ : LocalMux
    port map (
            O => \N__37558\,
            I => \N__37552\
        );

    \I__7990\ : Odrv4
    port map (
            O => \N__37555\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__7989\ : Odrv12
    port map (
            O => \N__37552\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__7988\ : InMux
    port map (
            O => \N__37547\,
            I => \N__37544\
        );

    \I__7987\ : LocalMux
    port map (
            O => \N__37544\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13\
        );

    \I__7986\ : InMux
    port map (
            O => \N__37541\,
            I => \N__37538\
        );

    \I__7985\ : LocalMux
    port map (
            O => \N__37538\,
            I => \N__37534\
        );

    \I__7984\ : InMux
    port map (
            O => \N__37537\,
            I => \N__37531\
        );

    \I__7983\ : Span4Mux_h
    port map (
            O => \N__37534\,
            I => \N__37528\
        );

    \I__7982\ : LocalMux
    port map (
            O => \N__37531\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__7981\ : Odrv4
    port map (
            O => \N__37528\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__7980\ : InMux
    port map (
            O => \N__37523\,
            I => \N__37520\
        );

    \I__7979\ : LocalMux
    port map (
            O => \N__37520\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9\
        );

    \I__7978\ : InMux
    port map (
            O => \N__37517\,
            I => \N__37514\
        );

    \I__7977\ : LocalMux
    port map (
            O => \N__37514\,
            I => \N__37510\
        );

    \I__7976\ : InMux
    port map (
            O => \N__37513\,
            I => \N__37507\
        );

    \I__7975\ : Span4Mux_h
    port map (
            O => \N__37510\,
            I => \N__37504\
        );

    \I__7974\ : LocalMux
    port map (
            O => \N__37507\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__7973\ : Odrv4
    port map (
            O => \N__37504\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__7972\ : CascadeMux
    port map (
            O => \N__37499\,
            I => \N__37496\
        );

    \I__7971\ : InMux
    port map (
            O => \N__37496\,
            I => \N__37493\
        );

    \I__7970\ : LocalMux
    port map (
            O => \N__37493\,
            I => \N__37490\
        );

    \I__7969\ : Odrv12
    port map (
            O => \N__37490\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6\
        );

    \I__7968\ : InMux
    port map (
            O => \N__37487\,
            I => \N__37483\
        );

    \I__7967\ : InMux
    port map (
            O => \N__37486\,
            I => \N__37480\
        );

    \I__7966\ : LocalMux
    port map (
            O => \N__37483\,
            I => \N__37477\
        );

    \I__7965\ : LocalMux
    port map (
            O => \N__37480\,
            I => \N__37474\
        );

    \I__7964\ : Odrv4
    port map (
            O => \N__37477\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__7963\ : Odrv12
    port map (
            O => \N__37474\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__7962\ : CascadeMux
    port map (
            O => \N__37469\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1_cascade_\
        );

    \I__7961\ : InMux
    port map (
            O => \N__37466\,
            I => \N__37457\
        );

    \I__7960\ : InMux
    port map (
            O => \N__37465\,
            I => \N__37457\
        );

    \I__7959\ : InMux
    port map (
            O => \N__37464\,
            I => \N__37457\
        );

    \I__7958\ : LocalMux
    port map (
            O => \N__37457\,
            I => \N__37451\
        );

    \I__7957\ : InMux
    port map (
            O => \N__37456\,
            I => \N__37444\
        );

    \I__7956\ : InMux
    port map (
            O => \N__37455\,
            I => \N__37444\
        );

    \I__7955\ : InMux
    port map (
            O => \N__37454\,
            I => \N__37444\
        );

    \I__7954\ : Odrv4
    port map (
            O => \N__37451\,
            I => \phase_controller_inst1.stoper_tr.N_20_li\
        );

    \I__7953\ : LocalMux
    port map (
            O => \N__37444\,
            I => \phase_controller_inst1.stoper_tr.N_20_li\
        );

    \I__7952\ : InMux
    port map (
            O => \N__37439\,
            I => \N__37434\
        );

    \I__7951\ : InMux
    port map (
            O => \N__37438\,
            I => \N__37429\
        );

    \I__7950\ : InMux
    port map (
            O => \N__37437\,
            I => \N__37429\
        );

    \I__7949\ : LocalMux
    port map (
            O => \N__37434\,
            I => \N__37424\
        );

    \I__7948\ : LocalMux
    port map (
            O => \N__37429\,
            I => \N__37424\
        );

    \I__7947\ : Span4Mux_h
    port map (
            O => \N__37424\,
            I => \N__37419\
        );

    \I__7946\ : InMux
    port map (
            O => \N__37423\,
            I => \N__37414\
        );

    \I__7945\ : InMux
    port map (
            O => \N__37422\,
            I => \N__37414\
        );

    \I__7944\ : Odrv4
    port map (
            O => \N__37419\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3\
        );

    \I__7943\ : LocalMux
    port map (
            O => \N__37414\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3\
        );

    \I__7942\ : InMux
    port map (
            O => \N__37409\,
            I => \N__37406\
        );

    \I__7941\ : LocalMux
    port map (
            O => \N__37406\,
            I => \N__37402\
        );

    \I__7940\ : CascadeMux
    port map (
            O => \N__37405\,
            I => \N__37399\
        );

    \I__7939\ : Span4Mux_v
    port map (
            O => \N__37402\,
            I => \N__37395\
        );

    \I__7938\ : InMux
    port map (
            O => \N__37399\,
            I => \N__37390\
        );

    \I__7937\ : InMux
    port map (
            O => \N__37398\,
            I => \N__37390\
        );

    \I__7936\ : Odrv4
    port map (
            O => \N__37395\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__7935\ : LocalMux
    port map (
            O => \N__37390\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__7934\ : InMux
    port map (
            O => \N__37385\,
            I => \N__37382\
        );

    \I__7933\ : LocalMux
    port map (
            O => \N__37382\,
            I => \N__37379\
        );

    \I__7932\ : Span4Mux_v
    port map (
            O => \N__37379\,
            I => \N__37375\
        );

    \I__7931\ : InMux
    port map (
            O => \N__37378\,
            I => \N__37372\
        );

    \I__7930\ : Span4Mux_v
    port map (
            O => \N__37375\,
            I => \N__37369\
        );

    \I__7929\ : LocalMux
    port map (
            O => \N__37372\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__7928\ : Odrv4
    port map (
            O => \N__37369\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__7927\ : InMux
    port map (
            O => \N__37364\,
            I => \N__37354\
        );

    \I__7926\ : InMux
    port map (
            O => \N__37363\,
            I => \N__37354\
        );

    \I__7925\ : InMux
    port map (
            O => \N__37362\,
            I => \N__37354\
        );

    \I__7924\ : InMux
    port map (
            O => \N__37361\,
            I => \N__37351\
        );

    \I__7923\ : LocalMux
    port map (
            O => \N__37354\,
            I => \N__37346\
        );

    \I__7922\ : LocalMux
    port map (
            O => \N__37351\,
            I => \N__37343\
        );

    \I__7921\ : InMux
    port map (
            O => \N__37350\,
            I => \N__37338\
        );

    \I__7920\ : InMux
    port map (
            O => \N__37349\,
            I => \N__37338\
        );

    \I__7919\ : Span4Mux_v
    port map (
            O => \N__37346\,
            I => \N__37333\
        );

    \I__7918\ : Span4Mux_h
    port map (
            O => \N__37343\,
            I => \N__37333\
        );

    \I__7917\ : LocalMux
    port map (
            O => \N__37338\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6\
        );

    \I__7916\ : Odrv4
    port map (
            O => \N__37333\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6\
        );

    \I__7915\ : InMux
    port map (
            O => \N__37328\,
            I => \N__37323\
        );

    \I__7914\ : InMux
    port map (
            O => \N__37327\,
            I => \N__37320\
        );

    \I__7913\ : InMux
    port map (
            O => \N__37326\,
            I => \N__37317\
        );

    \I__7912\ : LocalMux
    port map (
            O => \N__37323\,
            I => \N__37314\
        );

    \I__7911\ : LocalMux
    port map (
            O => \N__37320\,
            I => \N__37310\
        );

    \I__7910\ : LocalMux
    port map (
            O => \N__37317\,
            I => \N__37307\
        );

    \I__7909\ : Span4Mux_v
    port map (
            O => \N__37314\,
            I => \N__37304\
        );

    \I__7908\ : CascadeMux
    port map (
            O => \N__37313\,
            I => \N__37301\
        );

    \I__7907\ : Span4Mux_v
    port map (
            O => \N__37310\,
            I => \N__37296\
        );

    \I__7906\ : Span4Mux_h
    port map (
            O => \N__37307\,
            I => \N__37296\
        );

    \I__7905\ : Span4Mux_v
    port map (
            O => \N__37304\,
            I => \N__37293\
        );

    \I__7904\ : InMux
    port map (
            O => \N__37301\,
            I => \N__37290\
        );

    \I__7903\ : Span4Mux_v
    port map (
            O => \N__37296\,
            I => \N__37287\
        );

    \I__7902\ : Odrv4
    port map (
            O => \N__37293\,
            I => measured_delay_tr_7
        );

    \I__7901\ : LocalMux
    port map (
            O => \N__37290\,
            I => measured_delay_tr_7
        );

    \I__7900\ : Odrv4
    port map (
            O => \N__37287\,
            I => measured_delay_tr_7
        );

    \I__7899\ : InMux
    port map (
            O => \N__37280\,
            I => \N__37264\
        );

    \I__7898\ : InMux
    port map (
            O => \N__37279\,
            I => \N__37264\
        );

    \I__7897\ : InMux
    port map (
            O => \N__37278\,
            I => \N__37264\
        );

    \I__7896\ : InMux
    port map (
            O => \N__37277\,
            I => \N__37264\
        );

    \I__7895\ : InMux
    port map (
            O => \N__37276\,
            I => \N__37264\
        );

    \I__7894\ : InMux
    port map (
            O => \N__37275\,
            I => \N__37261\
        );

    \I__7893\ : LocalMux
    port map (
            O => \N__37264\,
            I => \N__37257\
        );

    \I__7892\ : LocalMux
    port map (
            O => \N__37261\,
            I => \N__37251\
        );

    \I__7891\ : InMux
    port map (
            O => \N__37260\,
            I => \N__37248\
        );

    \I__7890\ : Span4Mux_h
    port map (
            O => \N__37257\,
            I => \N__37245\
        );

    \I__7889\ : InMux
    port map (
            O => \N__37256\,
            I => \N__37238\
        );

    \I__7888\ : InMux
    port map (
            O => \N__37255\,
            I => \N__37238\
        );

    \I__7887\ : InMux
    port map (
            O => \N__37254\,
            I => \N__37238\
        );

    \I__7886\ : Span4Mux_h
    port map (
            O => \N__37251\,
            I => \N__37235\
        );

    \I__7885\ : LocalMux
    port map (
            O => \N__37248\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6\
        );

    \I__7884\ : Odrv4
    port map (
            O => \N__37245\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6\
        );

    \I__7883\ : LocalMux
    port map (
            O => \N__37238\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6\
        );

    \I__7882\ : Odrv4
    port map (
            O => \N__37235\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6\
        );

    \I__7881\ : InMux
    port map (
            O => \N__37226\,
            I => \N__37221\
        );

    \I__7880\ : InMux
    port map (
            O => \N__37225\,
            I => \N__37218\
        );

    \I__7879\ : InMux
    port map (
            O => \N__37224\,
            I => \N__37215\
        );

    \I__7878\ : LocalMux
    port map (
            O => \N__37221\,
            I => \N__37212\
        );

    \I__7877\ : LocalMux
    port map (
            O => \N__37218\,
            I => \N__37209\
        );

    \I__7876\ : LocalMux
    port map (
            O => \N__37215\,
            I => \N__37206\
        );

    \I__7875\ : Span4Mux_h
    port map (
            O => \N__37212\,
            I => \N__37203\
        );

    \I__7874\ : Span4Mux_v
    port map (
            O => \N__37209\,
            I => \N__37197\
        );

    \I__7873\ : Span4Mux_h
    port map (
            O => \N__37206\,
            I => \N__37197\
        );

    \I__7872\ : Span4Mux_v
    port map (
            O => \N__37203\,
            I => \N__37194\
        );

    \I__7871\ : InMux
    port map (
            O => \N__37202\,
            I => \N__37191\
        );

    \I__7870\ : Span4Mux_v
    port map (
            O => \N__37197\,
            I => \N__37188\
        );

    \I__7869\ : Odrv4
    port map (
            O => \N__37194\,
            I => measured_delay_tr_8
        );

    \I__7868\ : LocalMux
    port map (
            O => \N__37191\,
            I => measured_delay_tr_8
        );

    \I__7867\ : Odrv4
    port map (
            O => \N__37188\,
            I => measured_delay_tr_8
        );

    \I__7866\ : InMux
    port map (
            O => \N__37181\,
            I => \N__37178\
        );

    \I__7865\ : LocalMux
    port map (
            O => \N__37178\,
            I => \N__37175\
        );

    \I__7864\ : Span4Mux_v
    port map (
            O => \N__37175\,
            I => \N__37171\
        );

    \I__7863\ : InMux
    port map (
            O => \N__37174\,
            I => \N__37168\
        );

    \I__7862\ : Span4Mux_h
    port map (
            O => \N__37171\,
            I => \N__37165\
        );

    \I__7861\ : LocalMux
    port map (
            O => \N__37168\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__7860\ : Odrv4
    port map (
            O => \N__37165\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__7859\ : InMux
    port map (
            O => \N__37160\,
            I => \N__37157\
        );

    \I__7858\ : LocalMux
    port map (
            O => \N__37157\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_16\
        );

    \I__7857\ : InMux
    port map (
            O => \N__37154\,
            I => \N__37151\
        );

    \I__7856\ : LocalMux
    port map (
            O => \N__37151\,
            I => \N__37147\
        );

    \I__7855\ : InMux
    port map (
            O => \N__37150\,
            I => \N__37144\
        );

    \I__7854\ : Span4Mux_v
    port map (
            O => \N__37147\,
            I => \N__37141\
        );

    \I__7853\ : LocalMux
    port map (
            O => \N__37144\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__7852\ : Odrv4
    port map (
            O => \N__37141\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__7851\ : InMux
    port map (
            O => \N__37136\,
            I => \N__37133\
        );

    \I__7850\ : LocalMux
    port map (
            O => \N__37133\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_17\
        );

    \I__7849\ : InMux
    port map (
            O => \N__37130\,
            I => \N__37127\
        );

    \I__7848\ : LocalMux
    port map (
            O => \N__37127\,
            I => \N__37123\
        );

    \I__7847\ : InMux
    port map (
            O => \N__37126\,
            I => \N__37120\
        );

    \I__7846\ : Span4Mux_v
    port map (
            O => \N__37123\,
            I => \N__37117\
        );

    \I__7845\ : LocalMux
    port map (
            O => \N__37120\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__7844\ : Odrv4
    port map (
            O => \N__37117\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__7843\ : CascadeMux
    port map (
            O => \N__37112\,
            I => \N__37109\
        );

    \I__7842\ : InMux
    port map (
            O => \N__37109\,
            I => \N__37106\
        );

    \I__7841\ : LocalMux
    port map (
            O => \N__37106\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_18\
        );

    \I__7840\ : InMux
    port map (
            O => \N__37103\,
            I => \N__37100\
        );

    \I__7839\ : LocalMux
    port map (
            O => \N__37100\,
            I => \N__37096\
        );

    \I__7838\ : InMux
    port map (
            O => \N__37099\,
            I => \N__37093\
        );

    \I__7837\ : Span12Mux_v
    port map (
            O => \N__37096\,
            I => \N__37090\
        );

    \I__7836\ : LocalMux
    port map (
            O => \N__37093\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__7835\ : Odrv12
    port map (
            O => \N__37090\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__7834\ : InMux
    port map (
            O => \N__37085\,
            I => \N__37082\
        );

    \I__7833\ : LocalMux
    port map (
            O => \N__37082\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_19\
        );

    \I__7832\ : InMux
    port map (
            O => \N__37079\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__7831\ : InMux
    port map (
            O => \N__37076\,
            I => \N__37072\
        );

    \I__7830\ : InMux
    port map (
            O => \N__37075\,
            I => \N__37069\
        );

    \I__7829\ : LocalMux
    port map (
            O => \N__37072\,
            I => \N__37066\
        );

    \I__7828\ : LocalMux
    port map (
            O => \N__37069\,
            I => \N__37063\
        );

    \I__7827\ : Span4Mux_v
    port map (
            O => \N__37066\,
            I => \N__37059\
        );

    \I__7826\ : Span4Mux_h
    port map (
            O => \N__37063\,
            I => \N__37056\
        );

    \I__7825\ : InMux
    port map (
            O => \N__37062\,
            I => \N__37053\
        );

    \I__7824\ : Odrv4
    port map (
            O => \N__37059\,
            I => \phase_controller_slave.stoper_hc.time_passed11\
        );

    \I__7823\ : Odrv4
    port map (
            O => \N__37056\,
            I => \phase_controller_slave.stoper_hc.time_passed11\
        );

    \I__7822\ : LocalMux
    port map (
            O => \N__37053\,
            I => \phase_controller_slave.stoper_hc.time_passed11\
        );

    \I__7821\ : InMux
    port map (
            O => \N__37046\,
            I => \N__37043\
        );

    \I__7820\ : LocalMux
    port map (
            O => \N__37043\,
            I => \N__37040\
        );

    \I__7819\ : Span4Mux_v
    port map (
            O => \N__37040\,
            I => \N__37037\
        );

    \I__7818\ : Odrv4
    port map (
            O => \N__37037\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1\
        );

    \I__7817\ : InMux
    port map (
            O => \N__37034\,
            I => \N__37031\
        );

    \I__7816\ : LocalMux
    port map (
            O => \N__37031\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_9\
        );

    \I__7815\ : CascadeMux
    port map (
            O => \N__37028\,
            I => \N__37025\
        );

    \I__7814\ : InMux
    port map (
            O => \N__37025\,
            I => \N__37022\
        );

    \I__7813\ : LocalMux
    port map (
            O => \N__37022\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_9\
        );

    \I__7812\ : CascadeMux
    port map (
            O => \N__37019\,
            I => \N__37016\
        );

    \I__7811\ : InMux
    port map (
            O => \N__37016\,
            I => \N__37013\
        );

    \I__7810\ : LocalMux
    port map (
            O => \N__37013\,
            I => \N__37010\
        );

    \I__7809\ : Span4Mux_h
    port map (
            O => \N__37010\,
            I => \N__37007\
        );

    \I__7808\ : Odrv4
    port map (
            O => \N__37007\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_10\
        );

    \I__7807\ : InMux
    port map (
            O => \N__37004\,
            I => \N__37001\
        );

    \I__7806\ : LocalMux
    port map (
            O => \N__37001\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_10\
        );

    \I__7805\ : CascadeMux
    port map (
            O => \N__36998\,
            I => \N__36995\
        );

    \I__7804\ : InMux
    port map (
            O => \N__36995\,
            I => \N__36992\
        );

    \I__7803\ : LocalMux
    port map (
            O => \N__36992\,
            I => \N__36989\
        );

    \I__7802\ : Odrv4
    port map (
            O => \N__36989\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_11\
        );

    \I__7801\ : InMux
    port map (
            O => \N__36986\,
            I => \N__36983\
        );

    \I__7800\ : LocalMux
    port map (
            O => \N__36983\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_11\
        );

    \I__7799\ : CascadeMux
    port map (
            O => \N__36980\,
            I => \N__36977\
        );

    \I__7798\ : InMux
    port map (
            O => \N__36977\,
            I => \N__36974\
        );

    \I__7797\ : LocalMux
    port map (
            O => \N__36974\,
            I => \N__36971\
        );

    \I__7796\ : Odrv4
    port map (
            O => \N__36971\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_12\
        );

    \I__7795\ : InMux
    port map (
            O => \N__36968\,
            I => \N__36965\
        );

    \I__7794\ : LocalMux
    port map (
            O => \N__36965\,
            I => \N__36962\
        );

    \I__7793\ : Span4Mux_h
    port map (
            O => \N__36962\,
            I => \N__36958\
        );

    \I__7792\ : InMux
    port map (
            O => \N__36961\,
            I => \N__36955\
        );

    \I__7791\ : Span4Mux_v
    port map (
            O => \N__36958\,
            I => \N__36952\
        );

    \I__7790\ : LocalMux
    port map (
            O => \N__36955\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__7789\ : Odrv4
    port map (
            O => \N__36952\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__7788\ : InMux
    port map (
            O => \N__36947\,
            I => \N__36944\
        );

    \I__7787\ : LocalMux
    port map (
            O => \N__36944\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_12\
        );

    \I__7786\ : InMux
    port map (
            O => \N__36941\,
            I => \N__36938\
        );

    \I__7785\ : LocalMux
    port map (
            O => \N__36938\,
            I => \N__36935\
        );

    \I__7784\ : Span4Mux_h
    port map (
            O => \N__36935\,
            I => \N__36931\
        );

    \I__7783\ : InMux
    port map (
            O => \N__36934\,
            I => \N__36928\
        );

    \I__7782\ : Span4Mux_v
    port map (
            O => \N__36931\,
            I => \N__36925\
        );

    \I__7781\ : LocalMux
    port map (
            O => \N__36928\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__7780\ : Odrv4
    port map (
            O => \N__36925\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__7779\ : InMux
    port map (
            O => \N__36920\,
            I => \N__36917\
        );

    \I__7778\ : LocalMux
    port map (
            O => \N__36917\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_13\
        );

    \I__7777\ : CascadeMux
    port map (
            O => \N__36914\,
            I => \N__36911\
        );

    \I__7776\ : InMux
    port map (
            O => \N__36911\,
            I => \N__36908\
        );

    \I__7775\ : LocalMux
    port map (
            O => \N__36908\,
            I => \N__36905\
        );

    \I__7774\ : Span4Mux_v
    port map (
            O => \N__36905\,
            I => \N__36902\
        );

    \I__7773\ : Odrv4
    port map (
            O => \N__36902\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_14\
        );

    \I__7772\ : InMux
    port map (
            O => \N__36899\,
            I => \N__36896\
        );

    \I__7771\ : LocalMux
    port map (
            O => \N__36896\,
            I => \N__36892\
        );

    \I__7770\ : InMux
    port map (
            O => \N__36895\,
            I => \N__36889\
        );

    \I__7769\ : Span12Mux_h
    port map (
            O => \N__36892\,
            I => \N__36886\
        );

    \I__7768\ : LocalMux
    port map (
            O => \N__36889\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__7767\ : Odrv12
    port map (
            O => \N__36886\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__7766\ : InMux
    port map (
            O => \N__36881\,
            I => \N__36878\
        );

    \I__7765\ : LocalMux
    port map (
            O => \N__36878\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_14\
        );

    \I__7764\ : CascadeMux
    port map (
            O => \N__36875\,
            I => \N__36872\
        );

    \I__7763\ : InMux
    port map (
            O => \N__36872\,
            I => \N__36869\
        );

    \I__7762\ : LocalMux
    port map (
            O => \N__36869\,
            I => \N__36866\
        );

    \I__7761\ : Span4Mux_h
    port map (
            O => \N__36866\,
            I => \N__36863\
        );

    \I__7760\ : Odrv4
    port map (
            O => \N__36863\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_15\
        );

    \I__7759\ : InMux
    port map (
            O => \N__36860\,
            I => \N__36857\
        );

    \I__7758\ : LocalMux
    port map (
            O => \N__36857\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_15\
        );

    \I__7757\ : InMux
    port map (
            O => \N__36854\,
            I => \N__36851\
        );

    \I__7756\ : LocalMux
    port map (
            O => \N__36851\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_1\
        );

    \I__7755\ : CascadeMux
    port map (
            O => \N__36848\,
            I => \N__36845\
        );

    \I__7754\ : InMux
    port map (
            O => \N__36845\,
            I => \N__36842\
        );

    \I__7753\ : LocalMux
    port map (
            O => \N__36842\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_2\
        );

    \I__7752\ : InMux
    port map (
            O => \N__36839\,
            I => \N__36836\
        );

    \I__7751\ : LocalMux
    port map (
            O => \N__36836\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_2\
        );

    \I__7750\ : CascadeMux
    port map (
            O => \N__36833\,
            I => \N__36830\
        );

    \I__7749\ : InMux
    port map (
            O => \N__36830\,
            I => \N__36827\
        );

    \I__7748\ : LocalMux
    port map (
            O => \N__36827\,
            I => \N__36823\
        );

    \I__7747\ : InMux
    port map (
            O => \N__36826\,
            I => \N__36820\
        );

    \I__7746\ : Span4Mux_v
    port map (
            O => \N__36823\,
            I => \N__36817\
        );

    \I__7745\ : LocalMux
    port map (
            O => \N__36820\,
            I => \N__36814\
        );

    \I__7744\ : Odrv4
    port map (
            O => \N__36817\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__7743\ : Odrv4
    port map (
            O => \N__36814\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__7742\ : CascadeMux
    port map (
            O => \N__36809\,
            I => \N__36806\
        );

    \I__7741\ : InMux
    port map (
            O => \N__36806\,
            I => \N__36803\
        );

    \I__7740\ : LocalMux
    port map (
            O => \N__36803\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_3\
        );

    \I__7739\ : InMux
    port map (
            O => \N__36800\,
            I => \N__36797\
        );

    \I__7738\ : LocalMux
    port map (
            O => \N__36797\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_3\
        );

    \I__7737\ : CascadeMux
    port map (
            O => \N__36794\,
            I => \N__36791\
        );

    \I__7736\ : InMux
    port map (
            O => \N__36791\,
            I => \N__36788\
        );

    \I__7735\ : LocalMux
    port map (
            O => \N__36788\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_4\
        );

    \I__7734\ : InMux
    port map (
            O => \N__36785\,
            I => \N__36782\
        );

    \I__7733\ : LocalMux
    port map (
            O => \N__36782\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_4\
        );

    \I__7732\ : InMux
    port map (
            O => \N__36779\,
            I => \N__36776\
        );

    \I__7731\ : LocalMux
    port map (
            O => \N__36776\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_5\
        );

    \I__7730\ : CascadeMux
    port map (
            O => \N__36773\,
            I => \N__36770\
        );

    \I__7729\ : InMux
    port map (
            O => \N__36770\,
            I => \N__36767\
        );

    \I__7728\ : LocalMux
    port map (
            O => \N__36767\,
            I => \phase_controller_slave.stoper_hc.target_timeZ1Z_6\
        );

    \I__7727\ : InMux
    port map (
            O => \N__36764\,
            I => \N__36761\
        );

    \I__7726\ : LocalMux
    port map (
            O => \N__36761\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_6\
        );

    \I__7725\ : CascadeMux
    port map (
            O => \N__36758\,
            I => \N__36755\
        );

    \I__7724\ : InMux
    port map (
            O => \N__36755\,
            I => \N__36752\
        );

    \I__7723\ : LocalMux
    port map (
            O => \N__36752\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_7\
        );

    \I__7722\ : InMux
    port map (
            O => \N__36749\,
            I => \N__36746\
        );

    \I__7721\ : LocalMux
    port map (
            O => \N__36746\,
            I => \N__36743\
        );

    \I__7720\ : Sp12to4
    port map (
            O => \N__36743\,
            I => \N__36739\
        );

    \I__7719\ : InMux
    port map (
            O => \N__36742\,
            I => \N__36736\
        );

    \I__7718\ : Odrv12
    port map (
            O => \N__36739\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__7717\ : LocalMux
    port map (
            O => \N__36736\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__7716\ : InMux
    port map (
            O => \N__36731\,
            I => \N__36728\
        );

    \I__7715\ : LocalMux
    port map (
            O => \N__36728\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_7\
        );

    \I__7714\ : InMux
    port map (
            O => \N__36725\,
            I => \N__36722\
        );

    \I__7713\ : LocalMux
    port map (
            O => \N__36722\,
            I => \N__36719\
        );

    \I__7712\ : Span4Mux_v
    port map (
            O => \N__36719\,
            I => \N__36715\
        );

    \I__7711\ : InMux
    port map (
            O => \N__36718\,
            I => \N__36712\
        );

    \I__7710\ : Odrv4
    port map (
            O => \N__36715\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__7709\ : LocalMux
    port map (
            O => \N__36712\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__7708\ : InMux
    port map (
            O => \N__36707\,
            I => \N__36704\
        );

    \I__7707\ : LocalMux
    port map (
            O => \N__36704\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_8\
        );

    \I__7706\ : CascadeMux
    port map (
            O => \N__36701\,
            I => \N__36697\
        );

    \I__7705\ : CascadeMux
    port map (
            O => \N__36700\,
            I => \N__36694\
        );

    \I__7704\ : InMux
    port map (
            O => \N__36697\,
            I => \N__36688\
        );

    \I__7703\ : InMux
    port map (
            O => \N__36694\,
            I => \N__36688\
        );

    \I__7702\ : InMux
    port map (
            O => \N__36693\,
            I => \N__36685\
        );

    \I__7701\ : LocalMux
    port map (
            O => \N__36688\,
            I => \N__36682\
        );

    \I__7700\ : LocalMux
    port map (
            O => \N__36685\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__7699\ : Odrv12
    port map (
            O => \N__36682\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__7698\ : InMux
    port map (
            O => \N__36677\,
            I => \current_shift_inst.timer_s1.counter_cry_22\
        );

    \I__7697\ : InMux
    port map (
            O => \N__36674\,
            I => \N__36670\
        );

    \I__7696\ : InMux
    port map (
            O => \N__36673\,
            I => \N__36666\
        );

    \I__7695\ : LocalMux
    port map (
            O => \N__36670\,
            I => \N__36663\
        );

    \I__7694\ : InMux
    port map (
            O => \N__36669\,
            I => \N__36660\
        );

    \I__7693\ : LocalMux
    port map (
            O => \N__36666\,
            I => \N__36655\
        );

    \I__7692\ : Span4Mux_v
    port map (
            O => \N__36663\,
            I => \N__36655\
        );

    \I__7691\ : LocalMux
    port map (
            O => \N__36660\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__7690\ : Odrv4
    port map (
            O => \N__36655\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__7689\ : InMux
    port map (
            O => \N__36650\,
            I => \bfn_15_16_0_\
        );

    \I__7688\ : InMux
    port map (
            O => \N__36647\,
            I => \N__36643\
        );

    \I__7687\ : InMux
    port map (
            O => \N__36646\,
            I => \N__36639\
        );

    \I__7686\ : LocalMux
    port map (
            O => \N__36643\,
            I => \N__36636\
        );

    \I__7685\ : InMux
    port map (
            O => \N__36642\,
            I => \N__36633\
        );

    \I__7684\ : LocalMux
    port map (
            O => \N__36639\,
            I => \N__36628\
        );

    \I__7683\ : Span4Mux_v
    port map (
            O => \N__36636\,
            I => \N__36628\
        );

    \I__7682\ : LocalMux
    port map (
            O => \N__36633\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__7681\ : Odrv4
    port map (
            O => \N__36628\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__7680\ : InMux
    port map (
            O => \N__36623\,
            I => \current_shift_inst.timer_s1.counter_cry_24\
        );

    \I__7679\ : CascadeMux
    port map (
            O => \N__36620\,
            I => \N__36616\
        );

    \I__7678\ : CascadeMux
    port map (
            O => \N__36619\,
            I => \N__36613\
        );

    \I__7677\ : InMux
    port map (
            O => \N__36616\,
            I => \N__36607\
        );

    \I__7676\ : InMux
    port map (
            O => \N__36613\,
            I => \N__36607\
        );

    \I__7675\ : InMux
    port map (
            O => \N__36612\,
            I => \N__36604\
        );

    \I__7674\ : LocalMux
    port map (
            O => \N__36607\,
            I => \N__36601\
        );

    \I__7673\ : LocalMux
    port map (
            O => \N__36604\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__7672\ : Odrv4
    port map (
            O => \N__36601\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__7671\ : InMux
    port map (
            O => \N__36596\,
            I => \current_shift_inst.timer_s1.counter_cry_25\
        );

    \I__7670\ : CascadeMux
    port map (
            O => \N__36593\,
            I => \N__36589\
        );

    \I__7669\ : CascadeMux
    port map (
            O => \N__36592\,
            I => \N__36586\
        );

    \I__7668\ : InMux
    port map (
            O => \N__36589\,
            I => \N__36580\
        );

    \I__7667\ : InMux
    port map (
            O => \N__36586\,
            I => \N__36580\
        );

    \I__7666\ : InMux
    port map (
            O => \N__36585\,
            I => \N__36577\
        );

    \I__7665\ : LocalMux
    port map (
            O => \N__36580\,
            I => \N__36574\
        );

    \I__7664\ : LocalMux
    port map (
            O => \N__36577\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__7663\ : Odrv4
    port map (
            O => \N__36574\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__7662\ : InMux
    port map (
            O => \N__36569\,
            I => \current_shift_inst.timer_s1.counter_cry_26\
        );

    \I__7661\ : InMux
    port map (
            O => \N__36566\,
            I => \N__36562\
        );

    \I__7660\ : InMux
    port map (
            O => \N__36565\,
            I => \N__36559\
        );

    \I__7659\ : LocalMux
    port map (
            O => \N__36562\,
            I => \N__36556\
        );

    \I__7658\ : LocalMux
    port map (
            O => \N__36559\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__7657\ : Odrv12
    port map (
            O => \N__36556\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__7656\ : InMux
    port map (
            O => \N__36551\,
            I => \current_shift_inst.timer_s1.counter_cry_27\
        );

    \I__7655\ : InMux
    port map (
            O => \N__36548\,
            I => \N__36510\
        );

    \I__7654\ : InMux
    port map (
            O => \N__36547\,
            I => \N__36510\
        );

    \I__7653\ : InMux
    port map (
            O => \N__36546\,
            I => \N__36510\
        );

    \I__7652\ : InMux
    port map (
            O => \N__36545\,
            I => \N__36510\
        );

    \I__7651\ : InMux
    port map (
            O => \N__36544\,
            I => \N__36501\
        );

    \I__7650\ : InMux
    port map (
            O => \N__36543\,
            I => \N__36501\
        );

    \I__7649\ : InMux
    port map (
            O => \N__36542\,
            I => \N__36501\
        );

    \I__7648\ : InMux
    port map (
            O => \N__36541\,
            I => \N__36501\
        );

    \I__7647\ : InMux
    port map (
            O => \N__36540\,
            I => \N__36492\
        );

    \I__7646\ : InMux
    port map (
            O => \N__36539\,
            I => \N__36492\
        );

    \I__7645\ : InMux
    port map (
            O => \N__36538\,
            I => \N__36492\
        );

    \I__7644\ : InMux
    port map (
            O => \N__36537\,
            I => \N__36492\
        );

    \I__7643\ : InMux
    port map (
            O => \N__36536\,
            I => \N__36483\
        );

    \I__7642\ : InMux
    port map (
            O => \N__36535\,
            I => \N__36483\
        );

    \I__7641\ : InMux
    port map (
            O => \N__36534\,
            I => \N__36483\
        );

    \I__7640\ : InMux
    port map (
            O => \N__36533\,
            I => \N__36483\
        );

    \I__7639\ : InMux
    port map (
            O => \N__36532\,
            I => \N__36478\
        );

    \I__7638\ : InMux
    port map (
            O => \N__36531\,
            I => \N__36478\
        );

    \I__7637\ : InMux
    port map (
            O => \N__36530\,
            I => \N__36469\
        );

    \I__7636\ : InMux
    port map (
            O => \N__36529\,
            I => \N__36469\
        );

    \I__7635\ : InMux
    port map (
            O => \N__36528\,
            I => \N__36469\
        );

    \I__7634\ : InMux
    port map (
            O => \N__36527\,
            I => \N__36469\
        );

    \I__7633\ : InMux
    port map (
            O => \N__36526\,
            I => \N__36460\
        );

    \I__7632\ : InMux
    port map (
            O => \N__36525\,
            I => \N__36460\
        );

    \I__7631\ : InMux
    port map (
            O => \N__36524\,
            I => \N__36460\
        );

    \I__7630\ : InMux
    port map (
            O => \N__36523\,
            I => \N__36460\
        );

    \I__7629\ : InMux
    port map (
            O => \N__36522\,
            I => \N__36451\
        );

    \I__7628\ : InMux
    port map (
            O => \N__36521\,
            I => \N__36451\
        );

    \I__7627\ : InMux
    port map (
            O => \N__36520\,
            I => \N__36451\
        );

    \I__7626\ : InMux
    port map (
            O => \N__36519\,
            I => \N__36451\
        );

    \I__7625\ : LocalMux
    port map (
            O => \N__36510\,
            I => \N__36448\
        );

    \I__7624\ : LocalMux
    port map (
            O => \N__36501\,
            I => \N__36433\
        );

    \I__7623\ : LocalMux
    port map (
            O => \N__36492\,
            I => \N__36433\
        );

    \I__7622\ : LocalMux
    port map (
            O => \N__36483\,
            I => \N__36433\
        );

    \I__7621\ : LocalMux
    port map (
            O => \N__36478\,
            I => \N__36433\
        );

    \I__7620\ : LocalMux
    port map (
            O => \N__36469\,
            I => \N__36433\
        );

    \I__7619\ : LocalMux
    port map (
            O => \N__36460\,
            I => \N__36433\
        );

    \I__7618\ : LocalMux
    port map (
            O => \N__36451\,
            I => \N__36433\
        );

    \I__7617\ : Odrv4
    port map (
            O => \N__36448\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__7616\ : Odrv12
    port map (
            O => \N__36433\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__7615\ : InMux
    port map (
            O => \N__36428\,
            I => \current_shift_inst.timer_s1.counter_cry_28\
        );

    \I__7614\ : InMux
    port map (
            O => \N__36425\,
            I => \N__36421\
        );

    \I__7613\ : InMux
    port map (
            O => \N__36424\,
            I => \N__36418\
        );

    \I__7612\ : LocalMux
    port map (
            O => \N__36421\,
            I => \N__36415\
        );

    \I__7611\ : LocalMux
    port map (
            O => \N__36418\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__7610\ : Odrv12
    port map (
            O => \N__36415\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__7609\ : CEMux
    port map (
            O => \N__36410\,
            I => \N__36404\
        );

    \I__7608\ : CEMux
    port map (
            O => \N__36409\,
            I => \N__36401\
        );

    \I__7607\ : CEMux
    port map (
            O => \N__36408\,
            I => \N__36398\
        );

    \I__7606\ : CEMux
    port map (
            O => \N__36407\,
            I => \N__36395\
        );

    \I__7605\ : LocalMux
    port map (
            O => \N__36404\,
            I => \N__36390\
        );

    \I__7604\ : LocalMux
    port map (
            O => \N__36401\,
            I => \N__36390\
        );

    \I__7603\ : LocalMux
    port map (
            O => \N__36398\,
            I => \N__36385\
        );

    \I__7602\ : LocalMux
    port map (
            O => \N__36395\,
            I => \N__36385\
        );

    \I__7601\ : Span4Mux_v
    port map (
            O => \N__36390\,
            I => \N__36382\
        );

    \I__7600\ : Span4Mux_v
    port map (
            O => \N__36385\,
            I => \N__36377\
        );

    \I__7599\ : Span4Mux_h
    port map (
            O => \N__36382\,
            I => \N__36377\
        );

    \I__7598\ : Span4Mux_v
    port map (
            O => \N__36377\,
            I => \N__36374\
        );

    \I__7597\ : Odrv4
    port map (
            O => \N__36374\,
            I => \current_shift_inst.timer_s1.N_191_i\
        );

    \I__7596\ : InMux
    port map (
            O => \N__36371\,
            I => \N__36368\
        );

    \I__7595\ : LocalMux
    port map (
            O => \N__36368\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_0\
        );

    \I__7594\ : CascadeMux
    port map (
            O => \N__36365\,
            I => \N__36361\
        );

    \I__7593\ : CascadeMux
    port map (
            O => \N__36364\,
            I => \N__36358\
        );

    \I__7592\ : InMux
    port map (
            O => \N__36361\,
            I => \N__36352\
        );

    \I__7591\ : InMux
    port map (
            O => \N__36358\,
            I => \N__36352\
        );

    \I__7590\ : InMux
    port map (
            O => \N__36357\,
            I => \N__36349\
        );

    \I__7589\ : LocalMux
    port map (
            O => \N__36352\,
            I => \N__36346\
        );

    \I__7588\ : LocalMux
    port map (
            O => \N__36349\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__7587\ : Odrv12
    port map (
            O => \N__36346\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__7586\ : InMux
    port map (
            O => \N__36341\,
            I => \current_shift_inst.timer_s1.counter_cry_13\
        );

    \I__7585\ : CascadeMux
    port map (
            O => \N__36338\,
            I => \N__36334\
        );

    \I__7584\ : CascadeMux
    port map (
            O => \N__36337\,
            I => \N__36331\
        );

    \I__7583\ : InMux
    port map (
            O => \N__36334\,
            I => \N__36325\
        );

    \I__7582\ : InMux
    port map (
            O => \N__36331\,
            I => \N__36325\
        );

    \I__7581\ : InMux
    port map (
            O => \N__36330\,
            I => \N__36322\
        );

    \I__7580\ : LocalMux
    port map (
            O => \N__36325\,
            I => \N__36319\
        );

    \I__7579\ : LocalMux
    port map (
            O => \N__36322\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__7578\ : Odrv4
    port map (
            O => \N__36319\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__7577\ : InMux
    port map (
            O => \N__36314\,
            I => \current_shift_inst.timer_s1.counter_cry_14\
        );

    \I__7576\ : InMux
    port map (
            O => \N__36311\,
            I => \N__36307\
        );

    \I__7575\ : InMux
    port map (
            O => \N__36310\,
            I => \N__36304\
        );

    \I__7574\ : LocalMux
    port map (
            O => \N__36307\,
            I => \N__36300\
        );

    \I__7573\ : LocalMux
    port map (
            O => \N__36304\,
            I => \N__36297\
        );

    \I__7572\ : InMux
    port map (
            O => \N__36303\,
            I => \N__36294\
        );

    \I__7571\ : Span4Mux_h
    port map (
            O => \N__36300\,
            I => \N__36289\
        );

    \I__7570\ : Span4Mux_v
    port map (
            O => \N__36297\,
            I => \N__36289\
        );

    \I__7569\ : LocalMux
    port map (
            O => \N__36294\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__7568\ : Odrv4
    port map (
            O => \N__36289\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__7567\ : InMux
    port map (
            O => \N__36284\,
            I => \bfn_15_15_0_\
        );

    \I__7566\ : InMux
    port map (
            O => \N__36281\,
            I => \N__36277\
        );

    \I__7565\ : InMux
    port map (
            O => \N__36280\,
            I => \N__36273\
        );

    \I__7564\ : LocalMux
    port map (
            O => \N__36277\,
            I => \N__36270\
        );

    \I__7563\ : InMux
    port map (
            O => \N__36276\,
            I => \N__36267\
        );

    \I__7562\ : LocalMux
    port map (
            O => \N__36273\,
            I => \N__36262\
        );

    \I__7561\ : Span4Mux_v
    port map (
            O => \N__36270\,
            I => \N__36262\
        );

    \I__7560\ : LocalMux
    port map (
            O => \N__36267\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__7559\ : Odrv4
    port map (
            O => \N__36262\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__7558\ : InMux
    port map (
            O => \N__36257\,
            I => \current_shift_inst.timer_s1.counter_cry_16\
        );

    \I__7557\ : CascadeMux
    port map (
            O => \N__36254\,
            I => \N__36250\
        );

    \I__7556\ : CascadeMux
    port map (
            O => \N__36253\,
            I => \N__36247\
        );

    \I__7555\ : InMux
    port map (
            O => \N__36250\,
            I => \N__36241\
        );

    \I__7554\ : InMux
    port map (
            O => \N__36247\,
            I => \N__36241\
        );

    \I__7553\ : InMux
    port map (
            O => \N__36246\,
            I => \N__36238\
        );

    \I__7552\ : LocalMux
    port map (
            O => \N__36241\,
            I => \N__36235\
        );

    \I__7551\ : LocalMux
    port map (
            O => \N__36238\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__7550\ : Odrv4
    port map (
            O => \N__36235\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__7549\ : InMux
    port map (
            O => \N__36230\,
            I => \current_shift_inst.timer_s1.counter_cry_17\
        );

    \I__7548\ : CascadeMux
    port map (
            O => \N__36227\,
            I => \N__36223\
        );

    \I__7547\ : CascadeMux
    port map (
            O => \N__36226\,
            I => \N__36220\
        );

    \I__7546\ : InMux
    port map (
            O => \N__36223\,
            I => \N__36214\
        );

    \I__7545\ : InMux
    port map (
            O => \N__36220\,
            I => \N__36214\
        );

    \I__7544\ : InMux
    port map (
            O => \N__36219\,
            I => \N__36211\
        );

    \I__7543\ : LocalMux
    port map (
            O => \N__36214\,
            I => \N__36208\
        );

    \I__7542\ : LocalMux
    port map (
            O => \N__36211\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__7541\ : Odrv4
    port map (
            O => \N__36208\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__7540\ : InMux
    port map (
            O => \N__36203\,
            I => \current_shift_inst.timer_s1.counter_cry_18\
        );

    \I__7539\ : InMux
    port map (
            O => \N__36200\,
            I => \N__36193\
        );

    \I__7538\ : InMux
    port map (
            O => \N__36199\,
            I => \N__36193\
        );

    \I__7537\ : InMux
    port map (
            O => \N__36198\,
            I => \N__36190\
        );

    \I__7536\ : LocalMux
    port map (
            O => \N__36193\,
            I => \N__36187\
        );

    \I__7535\ : LocalMux
    port map (
            O => \N__36190\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__7534\ : Odrv4
    port map (
            O => \N__36187\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__7533\ : InMux
    port map (
            O => \N__36182\,
            I => \current_shift_inst.timer_s1.counter_cry_19\
        );

    \I__7532\ : InMux
    port map (
            O => \N__36179\,
            I => \N__36172\
        );

    \I__7531\ : InMux
    port map (
            O => \N__36178\,
            I => \N__36172\
        );

    \I__7530\ : InMux
    port map (
            O => \N__36177\,
            I => \N__36169\
        );

    \I__7529\ : LocalMux
    port map (
            O => \N__36172\,
            I => \N__36166\
        );

    \I__7528\ : LocalMux
    port map (
            O => \N__36169\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__7527\ : Odrv12
    port map (
            O => \N__36166\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__7526\ : InMux
    port map (
            O => \N__36161\,
            I => \current_shift_inst.timer_s1.counter_cry_20\
        );

    \I__7525\ : CascadeMux
    port map (
            O => \N__36158\,
            I => \N__36154\
        );

    \I__7524\ : CascadeMux
    port map (
            O => \N__36157\,
            I => \N__36151\
        );

    \I__7523\ : InMux
    port map (
            O => \N__36154\,
            I => \N__36145\
        );

    \I__7522\ : InMux
    port map (
            O => \N__36151\,
            I => \N__36145\
        );

    \I__7521\ : InMux
    port map (
            O => \N__36150\,
            I => \N__36142\
        );

    \I__7520\ : LocalMux
    port map (
            O => \N__36145\,
            I => \N__36139\
        );

    \I__7519\ : LocalMux
    port map (
            O => \N__36142\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__7518\ : Odrv12
    port map (
            O => \N__36139\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__7517\ : InMux
    port map (
            O => \N__36134\,
            I => \current_shift_inst.timer_s1.counter_cry_21\
        );

    \I__7516\ : InMux
    port map (
            O => \N__36131\,
            I => \N__36124\
        );

    \I__7515\ : InMux
    port map (
            O => \N__36130\,
            I => \N__36124\
        );

    \I__7514\ : InMux
    port map (
            O => \N__36129\,
            I => \N__36121\
        );

    \I__7513\ : LocalMux
    port map (
            O => \N__36124\,
            I => \N__36118\
        );

    \I__7512\ : LocalMux
    port map (
            O => \N__36121\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__7511\ : Odrv12
    port map (
            O => \N__36118\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__7510\ : InMux
    port map (
            O => \N__36113\,
            I => \current_shift_inst.timer_s1.counter_cry_5\
        );

    \I__7509\ : InMux
    port map (
            O => \N__36110\,
            I => \N__36103\
        );

    \I__7508\ : InMux
    port map (
            O => \N__36109\,
            I => \N__36103\
        );

    \I__7507\ : InMux
    port map (
            O => \N__36108\,
            I => \N__36100\
        );

    \I__7506\ : LocalMux
    port map (
            O => \N__36103\,
            I => \N__36097\
        );

    \I__7505\ : LocalMux
    port map (
            O => \N__36100\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__7504\ : Odrv12
    port map (
            O => \N__36097\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__7503\ : InMux
    port map (
            O => \N__36092\,
            I => \current_shift_inst.timer_s1.counter_cry_6\
        );

    \I__7502\ : CascadeMux
    port map (
            O => \N__36089\,
            I => \N__36086\
        );

    \I__7501\ : InMux
    port map (
            O => \N__36086\,
            I => \N__36083\
        );

    \I__7500\ : LocalMux
    port map (
            O => \N__36083\,
            I => \N__36079\
        );

    \I__7499\ : InMux
    port map (
            O => \N__36082\,
            I => \N__36075\
        );

    \I__7498\ : Span4Mux_v
    port map (
            O => \N__36079\,
            I => \N__36072\
        );

    \I__7497\ : InMux
    port map (
            O => \N__36078\,
            I => \N__36069\
        );

    \I__7496\ : LocalMux
    port map (
            O => \N__36075\,
            I => \N__36064\
        );

    \I__7495\ : Span4Mux_h
    port map (
            O => \N__36072\,
            I => \N__36064\
        );

    \I__7494\ : LocalMux
    port map (
            O => \N__36069\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__7493\ : Odrv4
    port map (
            O => \N__36064\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__7492\ : InMux
    port map (
            O => \N__36059\,
            I => \bfn_15_14_0_\
        );

    \I__7491\ : CascadeMux
    port map (
            O => \N__36056\,
            I => \N__36052\
        );

    \I__7490\ : InMux
    port map (
            O => \N__36055\,
            I => \N__36049\
        );

    \I__7489\ : InMux
    port map (
            O => \N__36052\,
            I => \N__36046\
        );

    \I__7488\ : LocalMux
    port map (
            O => \N__36049\,
            I => \N__36040\
        );

    \I__7487\ : LocalMux
    port map (
            O => \N__36046\,
            I => \N__36040\
        );

    \I__7486\ : InMux
    port map (
            O => \N__36045\,
            I => \N__36037\
        );

    \I__7485\ : Span4Mux_v
    port map (
            O => \N__36040\,
            I => \N__36034\
        );

    \I__7484\ : LocalMux
    port map (
            O => \N__36037\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__7483\ : Odrv4
    port map (
            O => \N__36034\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__7482\ : InMux
    port map (
            O => \N__36029\,
            I => \current_shift_inst.timer_s1.counter_cry_8\
        );

    \I__7481\ : CascadeMux
    port map (
            O => \N__36026\,
            I => \N__36022\
        );

    \I__7480\ : CascadeMux
    port map (
            O => \N__36025\,
            I => \N__36019\
        );

    \I__7479\ : InMux
    port map (
            O => \N__36022\,
            I => \N__36013\
        );

    \I__7478\ : InMux
    port map (
            O => \N__36019\,
            I => \N__36013\
        );

    \I__7477\ : InMux
    port map (
            O => \N__36018\,
            I => \N__36010\
        );

    \I__7476\ : LocalMux
    port map (
            O => \N__36013\,
            I => \N__36007\
        );

    \I__7475\ : LocalMux
    port map (
            O => \N__36010\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__7474\ : Odrv4
    port map (
            O => \N__36007\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__7473\ : InMux
    port map (
            O => \N__36002\,
            I => \current_shift_inst.timer_s1.counter_cry_9\
        );

    \I__7472\ : CascadeMux
    port map (
            O => \N__35999\,
            I => \N__35995\
        );

    \I__7471\ : CascadeMux
    port map (
            O => \N__35998\,
            I => \N__35992\
        );

    \I__7470\ : InMux
    port map (
            O => \N__35995\,
            I => \N__35986\
        );

    \I__7469\ : InMux
    port map (
            O => \N__35992\,
            I => \N__35986\
        );

    \I__7468\ : InMux
    port map (
            O => \N__35991\,
            I => \N__35983\
        );

    \I__7467\ : LocalMux
    port map (
            O => \N__35986\,
            I => \N__35980\
        );

    \I__7466\ : LocalMux
    port map (
            O => \N__35983\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__7465\ : Odrv12
    port map (
            O => \N__35980\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__7464\ : InMux
    port map (
            O => \N__35975\,
            I => \current_shift_inst.timer_s1.counter_cry_10\
        );

    \I__7463\ : InMux
    port map (
            O => \N__35972\,
            I => \N__35965\
        );

    \I__7462\ : InMux
    port map (
            O => \N__35971\,
            I => \N__35965\
        );

    \I__7461\ : InMux
    port map (
            O => \N__35970\,
            I => \N__35962\
        );

    \I__7460\ : LocalMux
    port map (
            O => \N__35965\,
            I => \N__35959\
        );

    \I__7459\ : LocalMux
    port map (
            O => \N__35962\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__7458\ : Odrv12
    port map (
            O => \N__35959\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__7457\ : InMux
    port map (
            O => \N__35954\,
            I => \current_shift_inst.timer_s1.counter_cry_11\
        );

    \I__7456\ : InMux
    port map (
            O => \N__35951\,
            I => \N__35944\
        );

    \I__7455\ : InMux
    port map (
            O => \N__35950\,
            I => \N__35944\
        );

    \I__7454\ : InMux
    port map (
            O => \N__35949\,
            I => \N__35941\
        );

    \I__7453\ : LocalMux
    port map (
            O => \N__35944\,
            I => \N__35938\
        );

    \I__7452\ : LocalMux
    port map (
            O => \N__35941\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__7451\ : Odrv4
    port map (
            O => \N__35938\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__7450\ : InMux
    port map (
            O => \N__35933\,
            I => \current_shift_inst.timer_s1.counter_cry_12\
        );

    \I__7449\ : InMux
    port map (
            O => \N__35930\,
            I => \N__35926\
        );

    \I__7448\ : InMux
    port map (
            O => \N__35929\,
            I => \N__35923\
        );

    \I__7447\ : LocalMux
    port map (
            O => \N__35926\,
            I => \N__35920\
        );

    \I__7446\ : LocalMux
    port map (
            O => \N__35923\,
            I => \N__35917\
        );

    \I__7445\ : Span4Mux_v
    port map (
            O => \N__35920\,
            I => \N__35911\
        );

    \I__7444\ : Span4Mux_h
    port map (
            O => \N__35917\,
            I => \N__35911\
        );

    \I__7443\ : InMux
    port map (
            O => \N__35916\,
            I => \N__35908\
        );

    \I__7442\ : Odrv4
    port map (
            O => \N__35911\,
            I => \delay_measurement_inst.hc_stateZ0Z_0\
        );

    \I__7441\ : LocalMux
    port map (
            O => \N__35908\,
            I => \delay_measurement_inst.hc_stateZ0Z_0\
        );

    \I__7440\ : InMux
    port map (
            O => \N__35903\,
            I => \N__35900\
        );

    \I__7439\ : LocalMux
    port map (
            O => \N__35900\,
            I => \N__35896\
        );

    \I__7438\ : InMux
    port map (
            O => \N__35899\,
            I => \N__35893\
        );

    \I__7437\ : Span4Mux_v
    port map (
            O => \N__35896\,
            I => \N__35888\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__35893\,
            I => \N__35888\
        );

    \I__7435\ : Span4Mux_v
    port map (
            O => \N__35888\,
            I => \N__35885\
        );

    \I__7434\ : Odrv4
    port map (
            O => \N__35885\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__7433\ : InMux
    port map (
            O => \N__35882\,
            I => \N__35878\
        );

    \I__7432\ : InMux
    port map (
            O => \N__35881\,
            I => \N__35875\
        );

    \I__7431\ : LocalMux
    port map (
            O => \N__35878\,
            I => \N__35872\
        );

    \I__7430\ : LocalMux
    port map (
            O => \N__35875\,
            I => \N__35869\
        );

    \I__7429\ : Span4Mux_v
    port map (
            O => \N__35872\,
            I => \N__35863\
        );

    \I__7428\ : Span4Mux_v
    port map (
            O => \N__35869\,
            I => \N__35863\
        );

    \I__7427\ : InMux
    port map (
            O => \N__35868\,
            I => \N__35860\
        );

    \I__7426\ : Odrv4
    port map (
            O => \N__35863\,
            I => \delay_measurement_inst.prev_hc_sigZ0\
        );

    \I__7425\ : LocalMux
    port map (
            O => \N__35860\,
            I => \delay_measurement_inst.prev_hc_sigZ0\
        );

    \I__7424\ : CascadeMux
    port map (
            O => \N__35855\,
            I => \N__35851\
        );

    \I__7423\ : InMux
    port map (
            O => \N__35854\,
            I => \N__35847\
        );

    \I__7422\ : InMux
    port map (
            O => \N__35851\,
            I => \N__35844\
        );

    \I__7421\ : InMux
    port map (
            O => \N__35850\,
            I => \N__35841\
        );

    \I__7420\ : LocalMux
    port map (
            O => \N__35847\,
            I => \N__35836\
        );

    \I__7419\ : LocalMux
    port map (
            O => \N__35844\,
            I => \N__35836\
        );

    \I__7418\ : LocalMux
    port map (
            O => \N__35841\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__7417\ : Odrv12
    port map (
            O => \N__35836\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__7416\ : InMux
    port map (
            O => \N__35831\,
            I => \bfn_15_13_0_\
        );

    \I__7415\ : CascadeMux
    port map (
            O => \N__35828\,
            I => \N__35824\
        );

    \I__7414\ : InMux
    port map (
            O => \N__35827\,
            I => \N__35821\
        );

    \I__7413\ : InMux
    port map (
            O => \N__35824\,
            I => \N__35817\
        );

    \I__7412\ : LocalMux
    port map (
            O => \N__35821\,
            I => \N__35814\
        );

    \I__7411\ : InMux
    port map (
            O => \N__35820\,
            I => \N__35811\
        );

    \I__7410\ : LocalMux
    port map (
            O => \N__35817\,
            I => \N__35808\
        );

    \I__7409\ : Odrv12
    port map (
            O => \N__35814\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__7408\ : LocalMux
    port map (
            O => \N__35811\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__7407\ : Odrv4
    port map (
            O => \N__35808\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__7406\ : InMux
    port map (
            O => \N__35801\,
            I => \current_shift_inst.timer_s1.counter_cry_0\
        );

    \I__7405\ : InMux
    port map (
            O => \N__35798\,
            I => \N__35791\
        );

    \I__7404\ : InMux
    port map (
            O => \N__35797\,
            I => \N__35791\
        );

    \I__7403\ : InMux
    port map (
            O => \N__35796\,
            I => \N__35788\
        );

    \I__7402\ : LocalMux
    port map (
            O => \N__35791\,
            I => \N__35785\
        );

    \I__7401\ : LocalMux
    port map (
            O => \N__35788\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__7400\ : Odrv4
    port map (
            O => \N__35785\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__7399\ : InMux
    port map (
            O => \N__35780\,
            I => \current_shift_inst.timer_s1.counter_cry_1\
        );

    \I__7398\ : InMux
    port map (
            O => \N__35777\,
            I => \N__35770\
        );

    \I__7397\ : InMux
    port map (
            O => \N__35776\,
            I => \N__35770\
        );

    \I__7396\ : InMux
    port map (
            O => \N__35775\,
            I => \N__35767\
        );

    \I__7395\ : LocalMux
    port map (
            O => \N__35770\,
            I => \N__35764\
        );

    \I__7394\ : LocalMux
    port map (
            O => \N__35767\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__7393\ : Odrv4
    port map (
            O => \N__35764\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__7392\ : InMux
    port map (
            O => \N__35759\,
            I => \current_shift_inst.timer_s1.counter_cry_2\
        );

    \I__7391\ : CascadeMux
    port map (
            O => \N__35756\,
            I => \N__35752\
        );

    \I__7390\ : CascadeMux
    port map (
            O => \N__35755\,
            I => \N__35749\
        );

    \I__7389\ : InMux
    port map (
            O => \N__35752\,
            I => \N__35744\
        );

    \I__7388\ : InMux
    port map (
            O => \N__35749\,
            I => \N__35744\
        );

    \I__7387\ : LocalMux
    port map (
            O => \N__35744\,
            I => \N__35740\
        );

    \I__7386\ : InMux
    port map (
            O => \N__35743\,
            I => \N__35737\
        );

    \I__7385\ : Span4Mux_h
    port map (
            O => \N__35740\,
            I => \N__35734\
        );

    \I__7384\ : LocalMux
    port map (
            O => \N__35737\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__7383\ : Odrv4
    port map (
            O => \N__35734\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__7382\ : InMux
    port map (
            O => \N__35729\,
            I => \current_shift_inst.timer_s1.counter_cry_3\
        );

    \I__7381\ : CascadeMux
    port map (
            O => \N__35726\,
            I => \N__35722\
        );

    \I__7380\ : CascadeMux
    port map (
            O => \N__35725\,
            I => \N__35719\
        );

    \I__7379\ : InMux
    port map (
            O => \N__35722\,
            I => \N__35713\
        );

    \I__7378\ : InMux
    port map (
            O => \N__35719\,
            I => \N__35713\
        );

    \I__7377\ : InMux
    port map (
            O => \N__35718\,
            I => \N__35710\
        );

    \I__7376\ : LocalMux
    port map (
            O => \N__35713\,
            I => \N__35707\
        );

    \I__7375\ : LocalMux
    port map (
            O => \N__35710\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__7374\ : Odrv12
    port map (
            O => \N__35707\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__7373\ : InMux
    port map (
            O => \N__35702\,
            I => \current_shift_inst.timer_s1.counter_cry_4\
        );

    \I__7372\ : CEMux
    port map (
            O => \N__35699\,
            I => \N__35684\
        );

    \I__7371\ : CEMux
    port map (
            O => \N__35698\,
            I => \N__35684\
        );

    \I__7370\ : CEMux
    port map (
            O => \N__35697\,
            I => \N__35684\
        );

    \I__7369\ : CEMux
    port map (
            O => \N__35696\,
            I => \N__35684\
        );

    \I__7368\ : CEMux
    port map (
            O => \N__35695\,
            I => \N__35684\
        );

    \I__7367\ : GlobalMux
    port map (
            O => \N__35684\,
            I => \N__35681\
        );

    \I__7366\ : gio2CtrlBuf
    port map (
            O => \N__35681\,
            I => \delay_measurement_inst.delay_hc_timer.N_321_i_g\
        );

    \I__7365\ : InMux
    port map (
            O => \N__35678\,
            I => \N__35674\
        );

    \I__7364\ : CascadeMux
    port map (
            O => \N__35677\,
            I => \N__35671\
        );

    \I__7363\ : LocalMux
    port map (
            O => \N__35674\,
            I => \N__35667\
        );

    \I__7362\ : InMux
    port map (
            O => \N__35671\,
            I => \N__35664\
        );

    \I__7361\ : InMux
    port map (
            O => \N__35670\,
            I => \N__35661\
        );

    \I__7360\ : Span4Mux_h
    port map (
            O => \N__35667\,
            I => \N__35658\
        );

    \I__7359\ : LocalMux
    port map (
            O => \N__35664\,
            I => \N__35651\
        );

    \I__7358\ : LocalMux
    port map (
            O => \N__35661\,
            I => \N__35651\
        );

    \I__7357\ : Span4Mux_h
    port map (
            O => \N__35658\,
            I => \N__35648\
        );

    \I__7356\ : InMux
    port map (
            O => \N__35657\,
            I => \N__35645\
        );

    \I__7355\ : InMux
    port map (
            O => \N__35656\,
            I => \N__35642\
        );

    \I__7354\ : Odrv12
    port map (
            O => \N__35651\,
            I => measured_delay_hc_10
        );

    \I__7353\ : Odrv4
    port map (
            O => \N__35648\,
            I => measured_delay_hc_10
        );

    \I__7352\ : LocalMux
    port map (
            O => \N__35645\,
            I => measured_delay_hc_10
        );

    \I__7351\ : LocalMux
    port map (
            O => \N__35642\,
            I => measured_delay_hc_10
        );

    \I__7350\ : InMux
    port map (
            O => \N__35633\,
            I => \N__35630\
        );

    \I__7349\ : LocalMux
    port map (
            O => \N__35630\,
            I => \N__35627\
        );

    \I__7348\ : Odrv4
    port map (
            O => \N__35627\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7\
        );

    \I__7347\ : InMux
    port map (
            O => \N__35624\,
            I => \N__35621\
        );

    \I__7346\ : LocalMux
    port map (
            O => \N__35621\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__7345\ : InMux
    port map (
            O => \N__35618\,
            I => \N__35615\
        );

    \I__7344\ : LocalMux
    port map (
            O => \N__35615\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__7343\ : CascadeMux
    port map (
            O => \N__35612\,
            I => \N__35609\
        );

    \I__7342\ : InMux
    port map (
            O => \N__35609\,
            I => \N__35606\
        );

    \I__7341\ : LocalMux
    port map (
            O => \N__35606\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__7340\ : InMux
    port map (
            O => \N__35603\,
            I => \N__35600\
        );

    \I__7339\ : LocalMux
    port map (
            O => \N__35600\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__7338\ : InMux
    port map (
            O => \N__35597\,
            I => \N__35594\
        );

    \I__7337\ : LocalMux
    port map (
            O => \N__35594\,
            I => \N__35589\
        );

    \I__7336\ : InMux
    port map (
            O => \N__35593\,
            I => \N__35584\
        );

    \I__7335\ : InMux
    port map (
            O => \N__35592\,
            I => \N__35584\
        );

    \I__7334\ : Span4Mux_h
    port map (
            O => \N__35589\,
            I => \N__35579\
        );

    \I__7333\ : LocalMux
    port map (
            O => \N__35584\,
            I => \N__35579\
        );

    \I__7332\ : Odrv4
    port map (
            O => \N__35579\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9\
        );

    \I__7331\ : InMux
    port map (
            O => \N__35576\,
            I => \N__35573\
        );

    \I__7330\ : LocalMux
    port map (
            O => \N__35573\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2\
        );

    \I__7329\ : InMux
    port map (
            O => \N__35570\,
            I => \N__35566\
        );

    \I__7328\ : InMux
    port map (
            O => \N__35569\,
            I => \N__35563\
        );

    \I__7327\ : LocalMux
    port map (
            O => \N__35566\,
            I => \N__35560\
        );

    \I__7326\ : LocalMux
    port map (
            O => \N__35563\,
            I => \N__35553\
        );

    \I__7325\ : Span4Mux_v
    port map (
            O => \N__35560\,
            I => \N__35553\
        );

    \I__7324\ : InMux
    port map (
            O => \N__35559\,
            I => \N__35548\
        );

    \I__7323\ : InMux
    port map (
            O => \N__35558\,
            I => \N__35548\
        );

    \I__7322\ : Odrv4
    port map (
            O => \N__35553\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__7321\ : LocalMux
    port map (
            O => \N__35548\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__7320\ : InMux
    port map (
            O => \N__35543\,
            I => \N__35540\
        );

    \I__7319\ : LocalMux
    port map (
            O => \N__35540\,
            I => \N__35535\
        );

    \I__7318\ : InMux
    port map (
            O => \N__35539\,
            I => \N__35532\
        );

    \I__7317\ : InMux
    port map (
            O => \N__35538\,
            I => \N__35529\
        );

    \I__7316\ : Odrv12
    port map (
            O => \N__35535\,
            I => \delay_measurement_inst.elapsed_time_hc_3\
        );

    \I__7315\ : LocalMux
    port map (
            O => \N__35532\,
            I => \delay_measurement_inst.elapsed_time_hc_3\
        );

    \I__7314\ : LocalMux
    port map (
            O => \N__35529\,
            I => \delay_measurement_inst.elapsed_time_hc_3\
        );

    \I__7313\ : InMux
    port map (
            O => \N__35522\,
            I => \N__35519\
        );

    \I__7312\ : LocalMux
    port map (
            O => \N__35519\,
            I => \N__35514\
        );

    \I__7311\ : CascadeMux
    port map (
            O => \N__35518\,
            I => \N__35510\
        );

    \I__7310\ : CascadeMux
    port map (
            O => \N__35517\,
            I => \N__35507\
        );

    \I__7309\ : Span4Mux_v
    port map (
            O => \N__35514\,
            I => \N__35504\
        );

    \I__7308\ : InMux
    port map (
            O => \N__35513\,
            I => \N__35501\
        );

    \I__7307\ : InMux
    port map (
            O => \N__35510\,
            I => \N__35497\
        );

    \I__7306\ : InMux
    port map (
            O => \N__35507\,
            I => \N__35494\
        );

    \I__7305\ : Span4Mux_h
    port map (
            O => \N__35504\,
            I => \N__35491\
        );

    \I__7304\ : LocalMux
    port map (
            O => \N__35501\,
            I => \N__35488\
        );

    \I__7303\ : CascadeMux
    port map (
            O => \N__35500\,
            I => \N__35485\
        );

    \I__7302\ : LocalMux
    port map (
            O => \N__35497\,
            I => \N__35482\
        );

    \I__7301\ : LocalMux
    port map (
            O => \N__35494\,
            I => \N__35479\
        );

    \I__7300\ : Span4Mux_h
    port map (
            O => \N__35491\,
            I => \N__35474\
        );

    \I__7299\ : Span4Mux_v
    port map (
            O => \N__35488\,
            I => \N__35474\
        );

    \I__7298\ : InMux
    port map (
            O => \N__35485\,
            I => \N__35471\
        );

    \I__7297\ : Sp12to4
    port map (
            O => \N__35482\,
            I => \N__35468\
        );

    \I__7296\ : Span4Mux_h
    port map (
            O => \N__35479\,
            I => \N__35465\
        );

    \I__7295\ : Span4Mux_h
    port map (
            O => \N__35474\,
            I => \N__35462\
        );

    \I__7294\ : LocalMux
    port map (
            O => \N__35471\,
            I => measured_delay_hc_3
        );

    \I__7293\ : Odrv12
    port map (
            O => \N__35468\,
            I => measured_delay_hc_3
        );

    \I__7292\ : Odrv4
    port map (
            O => \N__35465\,
            I => measured_delay_hc_3
        );

    \I__7291\ : Odrv4
    port map (
            O => \N__35462\,
            I => measured_delay_hc_3
        );

    \I__7290\ : InMux
    port map (
            O => \N__35453\,
            I => \N__35450\
        );

    \I__7289\ : LocalMux
    port map (
            O => \N__35450\,
            I => \N__35445\
        );

    \I__7288\ : InMux
    port map (
            O => \N__35449\,
            I => \N__35442\
        );

    \I__7287\ : InMux
    port map (
            O => \N__35448\,
            I => \N__35439\
        );

    \I__7286\ : Odrv12
    port map (
            O => \N__35445\,
            I => \delay_measurement_inst.elapsed_time_hc_4\
        );

    \I__7285\ : LocalMux
    port map (
            O => \N__35442\,
            I => \delay_measurement_inst.elapsed_time_hc_4\
        );

    \I__7284\ : LocalMux
    port map (
            O => \N__35439\,
            I => \delay_measurement_inst.elapsed_time_hc_4\
        );

    \I__7283\ : InMux
    port map (
            O => \N__35432\,
            I => \N__35428\
        );

    \I__7282\ : InMux
    port map (
            O => \N__35431\,
            I => \N__35423\
        );

    \I__7281\ : LocalMux
    port map (
            O => \N__35428\,
            I => \N__35419\
        );

    \I__7280\ : InMux
    port map (
            O => \N__35427\,
            I => \N__35416\
        );

    \I__7279\ : InMux
    port map (
            O => \N__35426\,
            I => \N__35413\
        );

    \I__7278\ : LocalMux
    port map (
            O => \N__35423\,
            I => \N__35410\
        );

    \I__7277\ : CascadeMux
    port map (
            O => \N__35422\,
            I => \N__35407\
        );

    \I__7276\ : Span4Mux_v
    port map (
            O => \N__35419\,
            I => \N__35404\
        );

    \I__7275\ : LocalMux
    port map (
            O => \N__35416\,
            I => \N__35401\
        );

    \I__7274\ : LocalMux
    port map (
            O => \N__35413\,
            I => \N__35398\
        );

    \I__7273\ : Span4Mux_v
    port map (
            O => \N__35410\,
            I => \N__35395\
        );

    \I__7272\ : InMux
    port map (
            O => \N__35407\,
            I => \N__35392\
        );

    \I__7271\ : Span4Mux_h
    port map (
            O => \N__35404\,
            I => \N__35389\
        );

    \I__7270\ : Sp12to4
    port map (
            O => \N__35401\,
            I => \N__35386\
        );

    \I__7269\ : Span4Mux_h
    port map (
            O => \N__35398\,
            I => \N__35383\
        );

    \I__7268\ : Span4Mux_h
    port map (
            O => \N__35395\,
            I => \N__35380\
        );

    \I__7267\ : LocalMux
    port map (
            O => \N__35392\,
            I => measured_delay_hc_4
        );

    \I__7266\ : Odrv4
    port map (
            O => \N__35389\,
            I => measured_delay_hc_4
        );

    \I__7265\ : Odrv12
    port map (
            O => \N__35386\,
            I => measured_delay_hc_4
        );

    \I__7264\ : Odrv4
    port map (
            O => \N__35383\,
            I => measured_delay_hc_4
        );

    \I__7263\ : Odrv4
    port map (
            O => \N__35380\,
            I => measured_delay_hc_4
        );

    \I__7262\ : InMux
    port map (
            O => \N__35369\,
            I => \N__35366\
        );

    \I__7261\ : LocalMux
    port map (
            O => \N__35366\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__7260\ : InMux
    port map (
            O => \N__35363\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__7259\ : InMux
    port map (
            O => \N__35360\,
            I => \N__35357\
        );

    \I__7258\ : LocalMux
    port map (
            O => \N__35357\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__7257\ : InMux
    port map (
            O => \N__35354\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__7256\ : InMux
    port map (
            O => \N__35351\,
            I => \N__35348\
        );

    \I__7255\ : LocalMux
    port map (
            O => \N__35348\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__7254\ : InMux
    port map (
            O => \N__35345\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__7253\ : CascadeMux
    port map (
            O => \N__35342\,
            I => \N__35339\
        );

    \I__7252\ : InMux
    port map (
            O => \N__35339\,
            I => \N__35336\
        );

    \I__7251\ : LocalMux
    port map (
            O => \N__35336\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__7250\ : InMux
    port map (
            O => \N__35333\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__7249\ : InMux
    port map (
            O => \N__35330\,
            I => \bfn_15_10_0_\
        );

    \I__7248\ : InMux
    port map (
            O => \N__35327\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__7247\ : InMux
    port map (
            O => \N__35324\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__7246\ : InMux
    port map (
            O => \N__35321\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__7245\ : InMux
    port map (
            O => \N__35318\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__7244\ : InMux
    port map (
            O => \N__35315\,
            I => \N__35306\
        );

    \I__7243\ : InMux
    port map (
            O => \N__35314\,
            I => \N__35306\
        );

    \I__7242\ : InMux
    port map (
            O => \N__35313\,
            I => \N__35306\
        );

    \I__7241\ : LocalMux
    port map (
            O => \N__35306\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__7240\ : InMux
    port map (
            O => \N__35303\,
            I => \N__35299\
        );

    \I__7239\ : InMux
    port map (
            O => \N__35302\,
            I => \N__35295\
        );

    \I__7238\ : LocalMux
    port map (
            O => \N__35299\,
            I => \N__35292\
        );

    \I__7237\ : InMux
    port map (
            O => \N__35298\,
            I => \N__35289\
        );

    \I__7236\ : LocalMux
    port map (
            O => \N__35295\,
            I => \N__35285\
        );

    \I__7235\ : Span4Mux_h
    port map (
            O => \N__35292\,
            I => \N__35280\
        );

    \I__7234\ : LocalMux
    port map (
            O => \N__35289\,
            I => \N__35280\
        );

    \I__7233\ : InMux
    port map (
            O => \N__35288\,
            I => \N__35277\
        );

    \I__7232\ : Odrv4
    port map (
            O => \N__35285\,
            I => \delay_measurement_inst.delay_hc_reg3lto14\
        );

    \I__7231\ : Odrv4
    port map (
            O => \N__35280\,
            I => \delay_measurement_inst.delay_hc_reg3lto14\
        );

    \I__7230\ : LocalMux
    port map (
            O => \N__35277\,
            I => \delay_measurement_inst.delay_hc_reg3lto14\
        );

    \I__7229\ : InMux
    port map (
            O => \N__35270\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__7228\ : CascadeMux
    port map (
            O => \N__35267\,
            I => \N__35264\
        );

    \I__7227\ : InMux
    port map (
            O => \N__35264\,
            I => \N__35261\
        );

    \I__7226\ : LocalMux
    port map (
            O => \N__35261\,
            I => \N__35253\
        );

    \I__7225\ : InMux
    port map (
            O => \N__35260\,
            I => \N__35250\
        );

    \I__7224\ : InMux
    port map (
            O => \N__35259\,
            I => \N__35246\
        );

    \I__7223\ : InMux
    port map (
            O => \N__35258\,
            I => \N__35243\
        );

    \I__7222\ : InMux
    port map (
            O => \N__35257\,
            I => \N__35240\
        );

    \I__7221\ : InMux
    port map (
            O => \N__35256\,
            I => \N__35237\
        );

    \I__7220\ : Span4Mux_h
    port map (
            O => \N__35253\,
            I => \N__35232\
        );

    \I__7219\ : LocalMux
    port map (
            O => \N__35250\,
            I => \N__35232\
        );

    \I__7218\ : InMux
    port map (
            O => \N__35249\,
            I => \N__35229\
        );

    \I__7217\ : LocalMux
    port map (
            O => \N__35246\,
            I => \N__35224\
        );

    \I__7216\ : LocalMux
    port map (
            O => \N__35243\,
            I => \N__35224\
        );

    \I__7215\ : LocalMux
    port map (
            O => \N__35240\,
            I => \delay_measurement_inst.delay_hc_reg3lto15\
        );

    \I__7214\ : LocalMux
    port map (
            O => \N__35237\,
            I => \delay_measurement_inst.delay_hc_reg3lto15\
        );

    \I__7213\ : Odrv4
    port map (
            O => \N__35232\,
            I => \delay_measurement_inst.delay_hc_reg3lto15\
        );

    \I__7212\ : LocalMux
    port map (
            O => \N__35229\,
            I => \delay_measurement_inst.delay_hc_reg3lto15\
        );

    \I__7211\ : Odrv4
    port map (
            O => \N__35224\,
            I => \delay_measurement_inst.delay_hc_reg3lto15\
        );

    \I__7210\ : InMux
    port map (
            O => \N__35213\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__7209\ : CascadeMux
    port map (
            O => \N__35210\,
            I => \N__35207\
        );

    \I__7208\ : InMux
    port map (
            O => \N__35207\,
            I => \N__35203\
        );

    \I__7207\ : InMux
    port map (
            O => \N__35206\,
            I => \N__35200\
        );

    \I__7206\ : LocalMux
    port map (
            O => \N__35203\,
            I => \N__35195\
        );

    \I__7205\ : LocalMux
    port map (
            O => \N__35200\,
            I => \N__35195\
        );

    \I__7204\ : Span4Mux_v
    port map (
            O => \N__35195\,
            I => \N__35191\
        );

    \I__7203\ : InMux
    port map (
            O => \N__35194\,
            I => \N__35188\
        );

    \I__7202\ : Odrv4
    port map (
            O => \N__35191\,
            I => \delay_measurement_inst.elapsed_time_hc_16\
        );

    \I__7201\ : LocalMux
    port map (
            O => \N__35188\,
            I => \delay_measurement_inst.elapsed_time_hc_16\
        );

    \I__7200\ : InMux
    port map (
            O => \N__35183\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__7199\ : InMux
    port map (
            O => \N__35180\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__7198\ : InMux
    port map (
            O => \N__35177\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__7197\ : InMux
    port map (
            O => \N__35174\,
            I => \bfn_15_9_0_\
        );

    \I__7196\ : CascadeMux
    port map (
            O => \N__35171\,
            I => \N__35167\
        );

    \I__7195\ : InMux
    port map (
            O => \N__35170\,
            I => \N__35162\
        );

    \I__7194\ : InMux
    port map (
            O => \N__35167\,
            I => \N__35162\
        );

    \I__7193\ : LocalMux
    port map (
            O => \N__35162\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__7192\ : InMux
    port map (
            O => \N__35159\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__7191\ : InMux
    port map (
            O => \N__35156\,
            I => \N__35150\
        );

    \I__7190\ : InMux
    port map (
            O => \N__35155\,
            I => \N__35150\
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__35150\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__7188\ : InMux
    port map (
            O => \N__35147\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__7187\ : InMux
    port map (
            O => \N__35144\,
            I => \N__35140\
        );

    \I__7186\ : InMux
    port map (
            O => \N__35143\,
            I => \N__35137\
        );

    \I__7185\ : LocalMux
    port map (
            O => \N__35140\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__7184\ : LocalMux
    port map (
            O => \N__35137\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__7183\ : InMux
    port map (
            O => \N__35132\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__7182\ : InMux
    port map (
            O => \N__35129\,
            I => \N__35125\
        );

    \I__7181\ : InMux
    port map (
            O => \N__35128\,
            I => \N__35121\
        );

    \I__7180\ : LocalMux
    port map (
            O => \N__35125\,
            I => \N__35118\
        );

    \I__7179\ : CascadeMux
    port map (
            O => \N__35124\,
            I => \N__35114\
        );

    \I__7178\ : LocalMux
    port map (
            O => \N__35121\,
            I => \N__35111\
        );

    \I__7177\ : Span4Mux_v
    port map (
            O => \N__35118\,
            I => \N__35108\
        );

    \I__7176\ : InMux
    port map (
            O => \N__35117\,
            I => \N__35105\
        );

    \I__7175\ : InMux
    port map (
            O => \N__35114\,
            I => \N__35102\
        );

    \I__7174\ : Span4Mux_v
    port map (
            O => \N__35111\,
            I => \N__35099\
        );

    \I__7173\ : Odrv4
    port map (
            O => \N__35108\,
            I => \delay_measurement_inst.delay_hc_reg3lto6\
        );

    \I__7172\ : LocalMux
    port map (
            O => \N__35105\,
            I => \delay_measurement_inst.delay_hc_reg3lto6\
        );

    \I__7171\ : LocalMux
    port map (
            O => \N__35102\,
            I => \delay_measurement_inst.delay_hc_reg3lto6\
        );

    \I__7170\ : Odrv4
    port map (
            O => \N__35099\,
            I => \delay_measurement_inst.delay_hc_reg3lto6\
        );

    \I__7169\ : InMux
    port map (
            O => \N__35090\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__7168\ : InMux
    port map (
            O => \N__35087\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__7167\ : InMux
    port map (
            O => \N__35084\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__7166\ : InMux
    port map (
            O => \N__35081\,
            I => \N__35077\
        );

    \I__7165\ : InMux
    port map (
            O => \N__35080\,
            I => \N__35072\
        );

    \I__7164\ : LocalMux
    port map (
            O => \N__35077\,
            I => \N__35069\
        );

    \I__7163\ : CascadeMux
    port map (
            O => \N__35076\,
            I => \N__35066\
        );

    \I__7162\ : InMux
    port map (
            O => \N__35075\,
            I => \N__35063\
        );

    \I__7161\ : LocalMux
    port map (
            O => \N__35072\,
            I => \N__35060\
        );

    \I__7160\ : Span4Mux_h
    port map (
            O => \N__35069\,
            I => \N__35057\
        );

    \I__7159\ : InMux
    port map (
            O => \N__35066\,
            I => \N__35054\
        );

    \I__7158\ : LocalMux
    port map (
            O => \N__35063\,
            I => \N__35049\
        );

    \I__7157\ : Span4Mux_h
    port map (
            O => \N__35060\,
            I => \N__35049\
        );

    \I__7156\ : Odrv4
    port map (
            O => \N__35057\,
            I => \delay_measurement_inst.delay_hc_reg3lto9\
        );

    \I__7155\ : LocalMux
    port map (
            O => \N__35054\,
            I => \delay_measurement_inst.delay_hc_reg3lto9\
        );

    \I__7154\ : Odrv4
    port map (
            O => \N__35049\,
            I => \delay_measurement_inst.delay_hc_reg3lto9\
        );

    \I__7153\ : InMux
    port map (
            O => \N__35042\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__7152\ : InMux
    port map (
            O => \N__35039\,
            I => \N__35035\
        );

    \I__7151\ : CascadeMux
    port map (
            O => \N__35038\,
            I => \N__35032\
        );

    \I__7150\ : LocalMux
    port map (
            O => \N__35035\,
            I => \N__35028\
        );

    \I__7149\ : InMux
    port map (
            O => \N__35032\,
            I => \N__35025\
        );

    \I__7148\ : InMux
    port map (
            O => \N__35031\,
            I => \N__35022\
        );

    \I__7147\ : Odrv4
    port map (
            O => \N__35028\,
            I => \delay_measurement_inst.elapsed_time_hc_10\
        );

    \I__7146\ : LocalMux
    port map (
            O => \N__35025\,
            I => \delay_measurement_inst.elapsed_time_hc_10\
        );

    \I__7145\ : LocalMux
    port map (
            O => \N__35022\,
            I => \delay_measurement_inst.elapsed_time_hc_10\
        );

    \I__7144\ : InMux
    port map (
            O => \N__35015\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__7143\ : CascadeMux
    port map (
            O => \N__35012\,
            I => \N__35008\
        );

    \I__7142\ : InMux
    port map (
            O => \N__35011\,
            I => \N__35003\
        );

    \I__7141\ : InMux
    port map (
            O => \N__35008\,
            I => \N__35003\
        );

    \I__7140\ : LocalMux
    port map (
            O => \N__35003\,
            I => \N__34999\
        );

    \I__7139\ : InMux
    port map (
            O => \N__35002\,
            I => \N__34996\
        );

    \I__7138\ : Span4Mux_v
    port map (
            O => \N__34999\,
            I => \N__34991\
        );

    \I__7137\ : LocalMux
    port map (
            O => \N__34996\,
            I => \N__34991\
        );

    \I__7136\ : Odrv4
    port map (
            O => \N__34991\,
            I => \delay_measurement_inst.elapsed_time_hc_11\
        );

    \I__7135\ : InMux
    port map (
            O => \N__34988\,
            I => \bfn_15_8_0_\
        );

    \I__7134\ : InMux
    port map (
            O => \N__34985\,
            I => \N__34978\
        );

    \I__7133\ : InMux
    port map (
            O => \N__34984\,
            I => \N__34978\
        );

    \I__7132\ : CascadeMux
    port map (
            O => \N__34983\,
            I => \N__34975\
        );

    \I__7131\ : LocalMux
    port map (
            O => \N__34978\,
            I => \N__34972\
        );

    \I__7130\ : InMux
    port map (
            O => \N__34975\,
            I => \N__34969\
        );

    \I__7129\ : Odrv4
    port map (
            O => \N__34972\,
            I => \delay_measurement_inst.elapsed_time_hc_12\
        );

    \I__7128\ : LocalMux
    port map (
            O => \N__34969\,
            I => \delay_measurement_inst.elapsed_time_hc_12\
        );

    \I__7127\ : InMux
    port map (
            O => \N__34964\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__7126\ : CascadeMux
    port map (
            O => \N__34961\,
            I => \N__34957\
        );

    \I__7125\ : InMux
    port map (
            O => \N__34960\,
            I => \N__34954\
        );

    \I__7124\ : InMux
    port map (
            O => \N__34957\,
            I => \N__34951\
        );

    \I__7123\ : LocalMux
    port map (
            O => \N__34954\,
            I => \N__34948\
        );

    \I__7122\ : LocalMux
    port map (
            O => \N__34951\,
            I => \N__34944\
        );

    \I__7121\ : Span4Mux_v
    port map (
            O => \N__34948\,
            I => \N__34941\
        );

    \I__7120\ : InMux
    port map (
            O => \N__34947\,
            I => \N__34938\
        );

    \I__7119\ : Span4Mux_h
    port map (
            O => \N__34944\,
            I => \N__34935\
        );

    \I__7118\ : Odrv4
    port map (
            O => \N__34941\,
            I => \delay_measurement_inst.elapsed_time_hc_13\
        );

    \I__7117\ : LocalMux
    port map (
            O => \N__34938\,
            I => \delay_measurement_inst.elapsed_time_hc_13\
        );

    \I__7116\ : Odrv4
    port map (
            O => \N__34935\,
            I => \delay_measurement_inst.elapsed_time_hc_13\
        );

    \I__7115\ : InMux
    port map (
            O => \N__34928\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__7114\ : InMux
    port map (
            O => \N__34925\,
            I => \N__34922\
        );

    \I__7113\ : LocalMux
    port map (
            O => \N__34922\,
            I => \N__34919\
        );

    \I__7112\ : Odrv12
    port map (
            O => \N__34919\,
            I => delay_tr_input_c
        );

    \I__7111\ : InMux
    port map (
            O => \N__34916\,
            I => \N__34913\
        );

    \I__7110\ : LocalMux
    port map (
            O => \N__34913\,
            I => delay_tr_d1
        );

    \I__7109\ : InMux
    port map (
            O => \N__34910\,
            I => \N__34907\
        );

    \I__7108\ : LocalMux
    port map (
            O => \N__34907\,
            I => \N__34901\
        );

    \I__7107\ : InMux
    port map (
            O => \N__34906\,
            I => \N__34894\
        );

    \I__7106\ : InMux
    port map (
            O => \N__34905\,
            I => \N__34894\
        );

    \I__7105\ : InMux
    port map (
            O => \N__34904\,
            I => \N__34894\
        );

    \I__7104\ : Span4Mux_v
    port map (
            O => \N__34901\,
            I => \N__34891\
        );

    \I__7103\ : LocalMux
    port map (
            O => \N__34894\,
            I => \N__34888\
        );

    \I__7102\ : Span4Mux_h
    port map (
            O => \N__34891\,
            I => \N__34885\
        );

    \I__7101\ : Span4Mux_v
    port map (
            O => \N__34888\,
            I => \N__34882\
        );

    \I__7100\ : Span4Mux_v
    port map (
            O => \N__34885\,
            I => \N__34879\
        );

    \I__7099\ : Span4Mux_v
    port map (
            O => \N__34882\,
            I => \N__34876\
        );

    \I__7098\ : Odrv4
    port map (
            O => \N__34879\,
            I => delay_tr_d2
        );

    \I__7097\ : Odrv4
    port map (
            O => \N__34876\,
            I => delay_tr_d2
        );

    \I__7096\ : InMux
    port map (
            O => \N__34871\,
            I => \N__34868\
        );

    \I__7095\ : LocalMux
    port map (
            O => \N__34868\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_4\
        );

    \I__7094\ : InMux
    port map (
            O => \N__34865\,
            I => \N__34862\
        );

    \I__7093\ : LocalMux
    port map (
            O => \N__34862\,
            I => \N__34859\
        );

    \I__7092\ : Span4Mux_v
    port map (
            O => \N__34859\,
            I => \N__34855\
        );

    \I__7091\ : InMux
    port map (
            O => \N__34858\,
            I => \N__34852\
        );

    \I__7090\ : Odrv4
    port map (
            O => \N__34855\,
            I => \delay_measurement_inst.elapsed_time_hc_1\
        );

    \I__7089\ : LocalMux
    port map (
            O => \N__34852\,
            I => \delay_measurement_inst.elapsed_time_hc_1\
        );

    \I__7088\ : InMux
    port map (
            O => \N__34847\,
            I => \N__34844\
        );

    \I__7087\ : LocalMux
    port map (
            O => \N__34844\,
            I => \N__34841\
        );

    \I__7086\ : Span4Mux_h
    port map (
            O => \N__34841\,
            I => \N__34836\
        );

    \I__7085\ : InMux
    port map (
            O => \N__34840\,
            I => \N__34833\
        );

    \I__7084\ : InMux
    port map (
            O => \N__34839\,
            I => \N__34830\
        );

    \I__7083\ : Odrv4
    port map (
            O => \N__34836\,
            I => \delay_measurement_inst.elapsed_time_hc_2\
        );

    \I__7082\ : LocalMux
    port map (
            O => \N__34833\,
            I => \delay_measurement_inst.elapsed_time_hc_2\
        );

    \I__7081\ : LocalMux
    port map (
            O => \N__34830\,
            I => \delay_measurement_inst.elapsed_time_hc_2\
        );

    \I__7080\ : InMux
    port map (
            O => \N__34823\,
            I => \N__34820\
        );

    \I__7079\ : LocalMux
    port map (
            O => \N__34820\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6\
        );

    \I__7078\ : InMux
    port map (
            O => \N__34817\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__7077\ : InMux
    port map (
            O => \N__34814\,
            I => \N__34810\
        );

    \I__7076\ : CascadeMux
    port map (
            O => \N__34813\,
            I => \N__34807\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__34810\,
            I => \N__34804\
        );

    \I__7074\ : InMux
    port map (
            O => \N__34807\,
            I => \N__34800\
        );

    \I__7073\ : Span4Mux_v
    port map (
            O => \N__34804\,
            I => \N__34797\
        );

    \I__7072\ : InMux
    port map (
            O => \N__34803\,
            I => \N__34794\
        );

    \I__7071\ : LocalMux
    port map (
            O => \N__34800\,
            I => \N__34791\
        );

    \I__7070\ : Odrv4
    port map (
            O => \N__34797\,
            I => \delay_measurement_inst.elapsed_time_hc_5\
        );

    \I__7069\ : LocalMux
    port map (
            O => \N__34794\,
            I => \delay_measurement_inst.elapsed_time_hc_5\
        );

    \I__7068\ : Odrv4
    port map (
            O => \N__34791\,
            I => \delay_measurement_inst.elapsed_time_hc_5\
        );

    \I__7067\ : InMux
    port map (
            O => \N__34784\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__7066\ : InMux
    port map (
            O => \N__34781\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12\
        );

    \I__7065\ : InMux
    port map (
            O => \N__34778\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13\
        );

    \I__7064\ : InMux
    port map (
            O => \N__34775\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14\
        );

    \I__7063\ : InMux
    port map (
            O => \N__34772\,
            I => \bfn_14_24_0_\
        );

    \I__7062\ : InMux
    port map (
            O => \N__34769\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16\
        );

    \I__7061\ : InMux
    port map (
            O => \N__34766\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17\
        );

    \I__7060\ : InMux
    port map (
            O => \N__34763\,
            I => \N__34760\
        );

    \I__7059\ : LocalMux
    port map (
            O => \N__34760\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13\
        );

    \I__7058\ : InMux
    port map (
            O => \N__34757\,
            I => \N__34754\
        );

    \I__7057\ : LocalMux
    port map (
            O => \N__34754\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17\
        );

    \I__7056\ : InMux
    port map (
            O => \N__34751\,
            I => \N__34748\
        );

    \I__7055\ : LocalMux
    port map (
            O => \N__34748\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18\
        );

    \I__7054\ : InMux
    port map (
            O => \N__34745\,
            I => \N__34742\
        );

    \I__7053\ : LocalMux
    port map (
            O => \N__34742\,
            I => \N__34739\
        );

    \I__7052\ : Span4Mux_v
    port map (
            O => \N__34739\,
            I => \N__34736\
        );

    \I__7051\ : Odrv4
    port map (
            O => \N__34736\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5\
        );

    \I__7050\ : InMux
    port map (
            O => \N__34733\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3\
        );

    \I__7049\ : InMux
    port map (
            O => \N__34730\,
            I => \N__34727\
        );

    \I__7048\ : LocalMux
    port map (
            O => \N__34727\,
            I => \N__34723\
        );

    \I__7047\ : InMux
    port map (
            O => \N__34726\,
            I => \N__34720\
        );

    \I__7046\ : Odrv4
    port map (
            O => \N__34723\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__7045\ : LocalMux
    port map (
            O => \N__34720\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__7044\ : InMux
    port map (
            O => \N__34715\,
            I => \N__34712\
        );

    \I__7043\ : LocalMux
    port map (
            O => \N__34712\,
            I => \N__34709\
        );

    \I__7042\ : Odrv4
    port map (
            O => \N__34709\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6\
        );

    \I__7041\ : InMux
    port map (
            O => \N__34706\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4\
        );

    \I__7040\ : InMux
    port map (
            O => \N__34703\,
            I => \N__34700\
        );

    \I__7039\ : LocalMux
    port map (
            O => \N__34700\,
            I => \N__34696\
        );

    \I__7038\ : InMux
    port map (
            O => \N__34699\,
            I => \N__34693\
        );

    \I__7037\ : Odrv4
    port map (
            O => \N__34696\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__7036\ : LocalMux
    port map (
            O => \N__34693\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__7035\ : InMux
    port map (
            O => \N__34688\,
            I => \N__34685\
        );

    \I__7034\ : LocalMux
    port map (
            O => \N__34685\,
            I => \N__34682\
        );

    \I__7033\ : Span4Mux_v
    port map (
            O => \N__34682\,
            I => \N__34679\
        );

    \I__7032\ : Span4Mux_h
    port map (
            O => \N__34679\,
            I => \N__34676\
        );

    \I__7031\ : Odrv4
    port map (
            O => \N__34676\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7\
        );

    \I__7030\ : InMux
    port map (
            O => \N__34673\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5\
        );

    \I__7029\ : InMux
    port map (
            O => \N__34670\,
            I => \N__34667\
        );

    \I__7028\ : LocalMux
    port map (
            O => \N__34667\,
            I => \N__34663\
        );

    \I__7027\ : InMux
    port map (
            O => \N__34666\,
            I => \N__34660\
        );

    \I__7026\ : Odrv4
    port map (
            O => \N__34663\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__7025\ : LocalMux
    port map (
            O => \N__34660\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__7024\ : CascadeMux
    port map (
            O => \N__34655\,
            I => \N__34652\
        );

    \I__7023\ : InMux
    port map (
            O => \N__34652\,
            I => \N__34649\
        );

    \I__7022\ : LocalMux
    port map (
            O => \N__34649\,
            I => \N__34646\
        );

    \I__7021\ : Odrv12
    port map (
            O => \N__34646\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8\
        );

    \I__7020\ : InMux
    port map (
            O => \N__34643\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6\
        );

    \I__7019\ : InMux
    port map (
            O => \N__34640\,
            I => \bfn_14_23_0_\
        );

    \I__7018\ : InMux
    port map (
            O => \N__34637\,
            I => \N__34633\
        );

    \I__7017\ : InMux
    port map (
            O => \N__34636\,
            I => \N__34630\
        );

    \I__7016\ : LocalMux
    port map (
            O => \N__34633\,
            I => \N__34627\
        );

    \I__7015\ : LocalMux
    port map (
            O => \N__34630\,
            I => \N__34624\
        );

    \I__7014\ : Odrv12
    port map (
            O => \N__34627\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__7013\ : Odrv4
    port map (
            O => \N__34624\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__7012\ : InMux
    port map (
            O => \N__34619\,
            I => \N__34616\
        );

    \I__7011\ : LocalMux
    port map (
            O => \N__34616\,
            I => \N__34613\
        );

    \I__7010\ : Odrv12
    port map (
            O => \N__34613\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10\
        );

    \I__7009\ : InMux
    port map (
            O => \N__34610\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8\
        );

    \I__7008\ : InMux
    port map (
            O => \N__34607\,
            I => \N__34603\
        );

    \I__7007\ : InMux
    port map (
            O => \N__34606\,
            I => \N__34600\
        );

    \I__7006\ : LocalMux
    port map (
            O => \N__34603\,
            I => \N__34597\
        );

    \I__7005\ : LocalMux
    port map (
            O => \N__34600\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__7004\ : Odrv4
    port map (
            O => \N__34597\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__7003\ : InMux
    port map (
            O => \N__34592\,
            I => \N__34589\
        );

    \I__7002\ : LocalMux
    port map (
            O => \N__34589\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11\
        );

    \I__7001\ : InMux
    port map (
            O => \N__34586\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9\
        );

    \I__7000\ : InMux
    port map (
            O => \N__34583\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10\
        );

    \I__6999\ : InMux
    port map (
            O => \N__34580\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11\
        );

    \I__6998\ : InMux
    port map (
            O => \N__34577\,
            I => \N__34574\
        );

    \I__6997\ : LocalMux
    port map (
            O => \N__34574\,
            I => \N__34571\
        );

    \I__6996\ : Odrv4
    port map (
            O => \N__34571\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0\
        );

    \I__6995\ : InMux
    port map (
            O => \N__34568\,
            I => \N__34565\
        );

    \I__6994\ : LocalMux
    port map (
            O => \N__34565\,
            I => \N__34561\
        );

    \I__6993\ : InMux
    port map (
            O => \N__34564\,
            I => \N__34558\
        );

    \I__6992\ : Span4Mux_s1_v
    port map (
            O => \N__34561\,
            I => \N__34552\
        );

    \I__6991\ : LocalMux
    port map (
            O => \N__34558\,
            I => \N__34552\
        );

    \I__6990\ : InMux
    port map (
            O => \N__34557\,
            I => \N__34549\
        );

    \I__6989\ : Span4Mux_v
    port map (
            O => \N__34552\,
            I => \N__34546\
        );

    \I__6988\ : LocalMux
    port map (
            O => \N__34549\,
            I => \N__34541\
        );

    \I__6987\ : Span4Mux_h
    port map (
            O => \N__34546\,
            I => \N__34538\
        );

    \I__6986\ : InMux
    port map (
            O => \N__34545\,
            I => \N__34531\
        );

    \I__6985\ : InMux
    port map (
            O => \N__34544\,
            I => \N__34531\
        );

    \I__6984\ : Span4Mux_v
    port map (
            O => \N__34541\,
            I => \N__34528\
        );

    \I__6983\ : Sp12to4
    port map (
            O => \N__34538\,
            I => \N__34525\
        );

    \I__6982\ : InMux
    port map (
            O => \N__34537\,
            I => \N__34522\
        );

    \I__6981\ : CascadeMux
    port map (
            O => \N__34536\,
            I => \N__34519\
        );

    \I__6980\ : LocalMux
    port map (
            O => \N__34531\,
            I => \N__34516\
        );

    \I__6979\ : Span4Mux_h
    port map (
            O => \N__34528\,
            I => \N__34513\
        );

    \I__6978\ : Span12Mux_s11_v
    port map (
            O => \N__34525\,
            I => \N__34510\
        );

    \I__6977\ : LocalMux
    port map (
            O => \N__34522\,
            I => \N__34507\
        );

    \I__6976\ : InMux
    port map (
            O => \N__34519\,
            I => \N__34504\
        );

    \I__6975\ : Span4Mux_v
    port map (
            O => \N__34516\,
            I => \N__34501\
        );

    \I__6974\ : Sp12to4
    port map (
            O => \N__34513\,
            I => \N__34498\
        );

    \I__6973\ : Span12Mux_v
    port map (
            O => \N__34510\,
            I => \N__34491\
        );

    \I__6972\ : Sp12to4
    port map (
            O => \N__34507\,
            I => \N__34491\
        );

    \I__6971\ : LocalMux
    port map (
            O => \N__34504\,
            I => \N__34491\
        );

    \I__6970\ : Span4Mux_h
    port map (
            O => \N__34501\,
            I => \N__34488\
        );

    \I__6969\ : Span12Mux_v
    port map (
            O => \N__34498\,
            I => \N__34483\
        );

    \I__6968\ : Span12Mux_h
    port map (
            O => \N__34491\,
            I => \N__34483\
        );

    \I__6967\ : Span4Mux_v
    port map (
            O => \N__34488\,
            I => \N__34480\
        );

    \I__6966\ : Odrv12
    port map (
            O => \N__34483\,
            I => start_stop_c
        );

    \I__6965\ : Odrv4
    port map (
            O => \N__34480\,
            I => start_stop_c
        );

    \I__6964\ : InMux
    port map (
            O => \N__34475\,
            I => \N__34471\
        );

    \I__6963\ : CascadeMux
    port map (
            O => \N__34474\,
            I => \N__34468\
        );

    \I__6962\ : LocalMux
    port map (
            O => \N__34471\,
            I => \N__34465\
        );

    \I__6961\ : InMux
    port map (
            O => \N__34468\,
            I => \N__34462\
        );

    \I__6960\ : Span12Mux_s10_v
    port map (
            O => \N__34465\,
            I => \N__34459\
        );

    \I__6959\ : LocalMux
    port map (
            O => \N__34462\,
            I => shift_flag_start
        );

    \I__6958\ : Odrv12
    port map (
            O => \N__34459\,
            I => shift_flag_start
        );

    \I__6957\ : InMux
    port map (
            O => \N__34454\,
            I => \N__34448\
        );

    \I__6956\ : InMux
    port map (
            O => \N__34453\,
            I => \N__34448\
        );

    \I__6955\ : LocalMux
    port map (
            O => \N__34448\,
            I => \N__34445\
        );

    \I__6954\ : Span4Mux_v
    port map (
            O => \N__34445\,
            I => \N__34442\
        );

    \I__6953\ : Odrv4
    port map (
            O => \N__34442\,
            I => \phase_controller_slave.un1_startZ0\
        );

    \I__6952\ : InMux
    port map (
            O => \N__34439\,
            I => \N__34436\
        );

    \I__6951\ : LocalMux
    port map (
            O => \N__34436\,
            I => \N__34433\
        );

    \I__6950\ : Span4Mux_h
    port map (
            O => \N__34433\,
            I => \N__34428\
        );

    \I__6949\ : InMux
    port map (
            O => \N__34432\,
            I => \N__34423\
        );

    \I__6948\ : InMux
    port map (
            O => \N__34431\,
            I => \N__34423\
        );

    \I__6947\ : Odrv4
    port map (
            O => \N__34428\,
            I => \phase_controller_slave.stoper_tr.time_passed11\
        );

    \I__6946\ : LocalMux
    port map (
            O => \N__34423\,
            I => \phase_controller_slave.stoper_tr.time_passed11\
        );

    \I__6945\ : InMux
    port map (
            O => \N__34418\,
            I => \N__34412\
        );

    \I__6944\ : InMux
    port map (
            O => \N__34417\,
            I => \N__34412\
        );

    \I__6943\ : LocalMux
    port map (
            O => \N__34412\,
            I => \N__34407\
        );

    \I__6942\ : InMux
    port map (
            O => \N__34411\,
            I => \N__34404\
        );

    \I__6941\ : InMux
    port map (
            O => \N__34410\,
            I => \N__34399\
        );

    \I__6940\ : Span4Mux_v
    port map (
            O => \N__34407\,
            I => \N__34396\
        );

    \I__6939\ : LocalMux
    port map (
            O => \N__34404\,
            I => \N__34393\
        );

    \I__6938\ : InMux
    port map (
            O => \N__34403\,
            I => \N__34388\
        );

    \I__6937\ : InMux
    port map (
            O => \N__34402\,
            I => \N__34388\
        );

    \I__6936\ : LocalMux
    port map (
            O => \N__34399\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__6935\ : Odrv4
    port map (
            O => \N__34396\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__6934\ : Odrv4
    port map (
            O => \N__34393\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__6933\ : LocalMux
    port map (
            O => \N__34388\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__6932\ : InMux
    port map (
            O => \N__34379\,
            I => \N__34376\
        );

    \I__6931\ : LocalMux
    port map (
            O => \N__34376\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2\
        );

    \I__6930\ : CascadeMux
    port map (
            O => \N__34373\,
            I => \N__34370\
        );

    \I__6929\ : InMux
    port map (
            O => \N__34370\,
            I => \N__34366\
        );

    \I__6928\ : InMux
    port map (
            O => \N__34369\,
            I => \N__34362\
        );

    \I__6927\ : LocalMux
    port map (
            O => \N__34366\,
            I => \N__34359\
        );

    \I__6926\ : InMux
    port map (
            O => \N__34365\,
            I => \N__34356\
        );

    \I__6925\ : LocalMux
    port map (
            O => \N__34362\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__6924\ : Odrv12
    port map (
            O => \N__34359\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__6923\ : LocalMux
    port map (
            O => \N__34356\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__6922\ : InMux
    port map (
            O => \N__34349\,
            I => \N__34346\
        );

    \I__6921\ : LocalMux
    port map (
            O => \N__34346\,
            I => \N__34342\
        );

    \I__6920\ : InMux
    port map (
            O => \N__34345\,
            I => \N__34339\
        );

    \I__6919\ : Odrv12
    port map (
            O => \N__34342\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__6918\ : LocalMux
    port map (
            O => \N__34339\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__6917\ : InMux
    port map (
            O => \N__34334\,
            I => \N__34331\
        );

    \I__6916\ : LocalMux
    port map (
            O => \N__34331\,
            I => \N__34328\
        );

    \I__6915\ : Odrv4
    port map (
            O => \N__34328\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2\
        );

    \I__6914\ : InMux
    port map (
            O => \N__34325\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0\
        );

    \I__6913\ : InMux
    port map (
            O => \N__34322\,
            I => \N__34319\
        );

    \I__6912\ : LocalMux
    port map (
            O => \N__34319\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6\
        );

    \I__6911\ : CascadeMux
    port map (
            O => \N__34316\,
            I => \N__34313\
        );

    \I__6910\ : InMux
    port map (
            O => \N__34313\,
            I => \N__34310\
        );

    \I__6909\ : LocalMux
    port map (
            O => \N__34310\,
            I => \N__34306\
        );

    \I__6908\ : InMux
    port map (
            O => \N__34309\,
            I => \N__34303\
        );

    \I__6907\ : Odrv12
    port map (
            O => \N__34306\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__6906\ : LocalMux
    port map (
            O => \N__34303\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__6905\ : InMux
    port map (
            O => \N__34298\,
            I => \N__34295\
        );

    \I__6904\ : LocalMux
    port map (
            O => \N__34295\,
            I => \N__34292\
        );

    \I__6903\ : Span4Mux_v
    port map (
            O => \N__34292\,
            I => \N__34289\
        );

    \I__6902\ : Odrv4
    port map (
            O => \N__34289\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3\
        );

    \I__6901\ : InMux
    port map (
            O => \N__34286\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1\
        );

    \I__6900\ : InMux
    port map (
            O => \N__34283\,
            I => \N__34280\
        );

    \I__6899\ : LocalMux
    port map (
            O => \N__34280\,
            I => \N__34276\
        );

    \I__6898\ : InMux
    port map (
            O => \N__34279\,
            I => \N__34273\
        );

    \I__6897\ : Odrv4
    port map (
            O => \N__34276\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__6896\ : LocalMux
    port map (
            O => \N__34273\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__6895\ : CascadeMux
    port map (
            O => \N__34268\,
            I => \N__34265\
        );

    \I__6894\ : InMux
    port map (
            O => \N__34265\,
            I => \N__34262\
        );

    \I__6893\ : LocalMux
    port map (
            O => \N__34262\,
            I => \N__34259\
        );

    \I__6892\ : Odrv4
    port map (
            O => \N__34259\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4\
        );

    \I__6891\ : InMux
    port map (
            O => \N__34256\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2\
        );

    \I__6890\ : InMux
    port map (
            O => \N__34253\,
            I => \N__34250\
        );

    \I__6889\ : LocalMux
    port map (
            O => \N__34250\,
            I => \N__34246\
        );

    \I__6888\ : InMux
    port map (
            O => \N__34249\,
            I => \N__34243\
        );

    \I__6887\ : Odrv4
    port map (
            O => \N__34246\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__6886\ : LocalMux
    port map (
            O => \N__34243\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__6885\ : InMux
    port map (
            O => \N__34238\,
            I => \N__34235\
        );

    \I__6884\ : LocalMux
    port map (
            O => \N__34235\,
            I => \N__34232\
        );

    \I__6883\ : Span4Mux_h
    port map (
            O => \N__34232\,
            I => \N__34229\
        );

    \I__6882\ : Odrv4
    port map (
            O => \N__34229\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3\
        );

    \I__6881\ : CascadeMux
    port map (
            O => \N__34226\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3Z0Z_3_cascade_\
        );

    \I__6880\ : InMux
    port map (
            O => \N__34223\,
            I => \N__34220\
        );

    \I__6879\ : LocalMux
    port map (
            O => \N__34220\,
            I => \N__34217\
        );

    \I__6878\ : Span4Mux_h
    port map (
            O => \N__34217\,
            I => \N__34214\
        );

    \I__6877\ : Odrv4
    port map (
            O => \N__34214\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_5Z0Z_3\
        );

    \I__6876\ : CascadeMux
    port map (
            O => \N__34211\,
            I => \phase_controller_slave.stoper_hc.time_passed11_cascade_\
        );

    \I__6875\ : InMux
    port map (
            O => \N__34208\,
            I => \N__34205\
        );

    \I__6874\ : LocalMux
    port map (
            O => \N__34205\,
            I => \N__34202\
        );

    \I__6873\ : Odrv4
    port map (
            O => \N__34202\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1\
        );

    \I__6872\ : InMux
    port map (
            O => \N__34199\,
            I => \N__34196\
        );

    \I__6871\ : LocalMux
    port map (
            O => \N__34196\,
            I => \N__34193\
        );

    \I__6870\ : Span4Mux_v
    port map (
            O => \N__34193\,
            I => \N__34190\
        );

    \I__6869\ : Odrv4
    port map (
            O => \N__34190\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8\
        );

    \I__6868\ : CascadeMux
    port map (
            O => \N__34187\,
            I => \N__34184\
        );

    \I__6867\ : InMux
    port map (
            O => \N__34184\,
            I => \N__34181\
        );

    \I__6866\ : LocalMux
    port map (
            O => \N__34181\,
            I => \N__34178\
        );

    \I__6865\ : Span4Mux_h
    port map (
            O => \N__34178\,
            I => \N__34175\
        );

    \I__6864\ : Odrv4
    port map (
            O => \N__34175\,
            I => \phase_controller_slave.stoper_hc.time_passed_1_sqmuxa\
        );

    \I__6863\ : CascadeMux
    port map (
            O => \N__34172\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\
        );

    \I__6862\ : InMux
    port map (
            O => \N__34169\,
            I => \N__34166\
        );

    \I__6861\ : LocalMux
    port map (
            O => \N__34166\,
            I => \N__34162\
        );

    \I__6860\ : InMux
    port map (
            O => \N__34165\,
            I => \N__34159\
        );

    \I__6859\ : Span4Mux_v
    port map (
            O => \N__34162\,
            I => \N__34155\
        );

    \I__6858\ : LocalMux
    port map (
            O => \N__34159\,
            I => \N__34152\
        );

    \I__6857\ : CascadeMux
    port map (
            O => \N__34158\,
            I => \N__34147\
        );

    \I__6856\ : Span4Mux_h
    port map (
            O => \N__34155\,
            I => \N__34144\
        );

    \I__6855\ : Span4Mux_v
    port map (
            O => \N__34152\,
            I => \N__34141\
        );

    \I__6854\ : InMux
    port map (
            O => \N__34151\,
            I => \N__34138\
        );

    \I__6853\ : InMux
    port map (
            O => \N__34150\,
            I => \N__34135\
        );

    \I__6852\ : InMux
    port map (
            O => \N__34147\,
            I => \N__34132\
        );

    \I__6851\ : Span4Mux_h
    port map (
            O => \N__34144\,
            I => \N__34125\
        );

    \I__6850\ : Span4Mux_v
    port map (
            O => \N__34141\,
            I => \N__34125\
        );

    \I__6849\ : LocalMux
    port map (
            O => \N__34138\,
            I => \N__34125\
        );

    \I__6848\ : LocalMux
    port map (
            O => \N__34135\,
            I => \N__34122\
        );

    \I__6847\ : LocalMux
    port map (
            O => \N__34132\,
            I => measured_delay_hc_6
        );

    \I__6846\ : Odrv4
    port map (
            O => \N__34125\,
            I => measured_delay_hc_6
        );

    \I__6845\ : Odrv4
    port map (
            O => \N__34122\,
            I => measured_delay_hc_6
        );

    \I__6844\ : InMux
    port map (
            O => \N__34115\,
            I => \N__34111\
        );

    \I__6843\ : CascadeMux
    port map (
            O => \N__34114\,
            I => \N__34108\
        );

    \I__6842\ : LocalMux
    port map (
            O => \N__34111\,
            I => \N__34103\
        );

    \I__6841\ : InMux
    port map (
            O => \N__34108\,
            I => \N__34100\
        );

    \I__6840\ : InMux
    port map (
            O => \N__34107\,
            I => \N__34096\
        );

    \I__6839\ : CascadeMux
    port map (
            O => \N__34106\,
            I => \N__34093\
        );

    \I__6838\ : Span4Mux_v
    port map (
            O => \N__34103\,
            I => \N__34090\
        );

    \I__6837\ : LocalMux
    port map (
            O => \N__34100\,
            I => \N__34087\
        );

    \I__6836\ : InMux
    port map (
            O => \N__34099\,
            I => \N__34084\
        );

    \I__6835\ : LocalMux
    port map (
            O => \N__34096\,
            I => \N__34081\
        );

    \I__6834\ : InMux
    port map (
            O => \N__34093\,
            I => \N__34078\
        );

    \I__6833\ : Span4Mux_v
    port map (
            O => \N__34090\,
            I => \N__34075\
        );

    \I__6832\ : Span12Mux_h
    port map (
            O => \N__34087\,
            I => \N__34072\
        );

    \I__6831\ : LocalMux
    port map (
            O => \N__34084\,
            I => \N__34069\
        );

    \I__6830\ : Span4Mux_v
    port map (
            O => \N__34081\,
            I => \N__34066\
        );

    \I__6829\ : LocalMux
    port map (
            O => \N__34078\,
            I => measured_delay_hc_2
        );

    \I__6828\ : Odrv4
    port map (
            O => \N__34075\,
            I => measured_delay_hc_2
        );

    \I__6827\ : Odrv12
    port map (
            O => \N__34072\,
            I => measured_delay_hc_2
        );

    \I__6826\ : Odrv4
    port map (
            O => \N__34069\,
            I => measured_delay_hc_2
        );

    \I__6825\ : Odrv4
    port map (
            O => \N__34066\,
            I => measured_delay_hc_2
        );

    \I__6824\ : CascadeMux
    port map (
            O => \N__34055\,
            I => \N__34052\
        );

    \I__6823\ : InMux
    port map (
            O => \N__34052\,
            I => \N__34049\
        );

    \I__6822\ : LocalMux
    port map (
            O => \N__34049\,
            I => \N__34043\
        );

    \I__6821\ : InMux
    port map (
            O => \N__34048\,
            I => \N__34040\
        );

    \I__6820\ : InMux
    port map (
            O => \N__34047\,
            I => \N__34037\
        );

    \I__6819\ : CascadeMux
    port map (
            O => \N__34046\,
            I => \N__34034\
        );

    \I__6818\ : Span4Mux_h
    port map (
            O => \N__34043\,
            I => \N__34031\
        );

    \I__6817\ : LocalMux
    port map (
            O => \N__34040\,
            I => \N__34024\
        );

    \I__6816\ : LocalMux
    port map (
            O => \N__34037\,
            I => \N__34024\
        );

    \I__6815\ : InMux
    port map (
            O => \N__34034\,
            I => \N__34021\
        );

    \I__6814\ : Span4Mux_v
    port map (
            O => \N__34031\,
            I => \N__34018\
        );

    \I__6813\ : InMux
    port map (
            O => \N__34030\,
            I => \N__34015\
        );

    \I__6812\ : InMux
    port map (
            O => \N__34029\,
            I => \N__34012\
        );

    \I__6811\ : Span4Mux_v
    port map (
            O => \N__34024\,
            I => \N__34009\
        );

    \I__6810\ : LocalMux
    port map (
            O => \N__34021\,
            I => measured_delay_hc_9
        );

    \I__6809\ : Odrv4
    port map (
            O => \N__34018\,
            I => measured_delay_hc_9
        );

    \I__6808\ : LocalMux
    port map (
            O => \N__34015\,
            I => measured_delay_hc_9
        );

    \I__6807\ : LocalMux
    port map (
            O => \N__34012\,
            I => measured_delay_hc_9
        );

    \I__6806\ : Odrv4
    port map (
            O => \N__34009\,
            I => measured_delay_hc_9
        );

    \I__6805\ : InMux
    port map (
            O => \N__33998\,
            I => \N__33995\
        );

    \I__6804\ : LocalMux
    port map (
            O => \N__33995\,
            I => \N__33992\
        );

    \I__6803\ : Span4Mux_v
    port map (
            O => \N__33992\,
            I => \N__33989\
        );

    \I__6802\ : Odrv4
    port map (
            O => \N__33989\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7\
        );

    \I__6801\ : InMux
    port map (
            O => \N__33986\,
            I => \N__33983\
        );

    \I__6800\ : LocalMux
    port map (
            O => \N__33983\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_9\
        );

    \I__6799\ : InMux
    port map (
            O => \N__33980\,
            I => \N__33977\
        );

    \I__6798\ : LocalMux
    port map (
            O => \N__33977\,
            I => \N__33974\
        );

    \I__6797\ : Span4Mux_v
    port map (
            O => \N__33974\,
            I => \N__33971\
        );

    \I__6796\ : Odrv4
    port map (
            O => \N__33971\,
            I => \current_shift_inst.un4_control_input_axb_9\
        );

    \I__6795\ : InMux
    port map (
            O => \N__33968\,
            I => \N__33965\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__33965\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_16\
        );

    \I__6793\ : InMux
    port map (
            O => \N__33962\,
            I => \N__33959\
        );

    \I__6792\ : LocalMux
    port map (
            O => \N__33959\,
            I => \N__33956\
        );

    \I__6791\ : Span4Mux_h
    port map (
            O => \N__33956\,
            I => \N__33953\
        );

    \I__6790\ : Odrv4
    port map (
            O => \N__33953\,
            I => \current_shift_inst.un4_control_input_axb_16\
        );

    \I__6789\ : InMux
    port map (
            O => \N__33950\,
            I => \N__33947\
        );

    \I__6788\ : LocalMux
    port map (
            O => \N__33947\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_17\
        );

    \I__6787\ : InMux
    port map (
            O => \N__33944\,
            I => \N__33941\
        );

    \I__6786\ : LocalMux
    port map (
            O => \N__33941\,
            I => \N__33938\
        );

    \I__6785\ : Span4Mux_h
    port map (
            O => \N__33938\,
            I => \N__33935\
        );

    \I__6784\ : Odrv4
    port map (
            O => \N__33935\,
            I => \current_shift_inst.un4_control_input_axb_17\
        );

    \I__6783\ : InMux
    port map (
            O => \N__33932\,
            I => \N__33929\
        );

    \I__6782\ : LocalMux
    port map (
            O => \N__33929\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_13\
        );

    \I__6781\ : InMux
    port map (
            O => \N__33926\,
            I => \N__33923\
        );

    \I__6780\ : LocalMux
    port map (
            O => \N__33923\,
            I => \N__33920\
        );

    \I__6779\ : Odrv4
    port map (
            O => \N__33920\,
            I => \current_shift_inst.un4_control_input_axb_13\
        );

    \I__6778\ : InMux
    port map (
            O => \N__33917\,
            I => \N__33913\
        );

    \I__6777\ : InMux
    port map (
            O => \N__33916\,
            I => \N__33910\
        );

    \I__6776\ : LocalMux
    port map (
            O => \N__33913\,
            I => \N__33907\
        );

    \I__6775\ : LocalMux
    port map (
            O => \N__33910\,
            I => \N__33904\
        );

    \I__6774\ : Span4Mux_v
    port map (
            O => \N__33907\,
            I => \N__33898\
        );

    \I__6773\ : Span4Mux_h
    port map (
            O => \N__33904\,
            I => \N__33895\
        );

    \I__6772\ : InMux
    port map (
            O => \N__33903\,
            I => \N__33892\
        );

    \I__6771\ : InMux
    port map (
            O => \N__33902\,
            I => \N__33887\
        );

    \I__6770\ : InMux
    port map (
            O => \N__33901\,
            I => \N__33887\
        );

    \I__6769\ : Odrv4
    port map (
            O => \N__33898\,
            I => measured_delay_hc_15
        );

    \I__6768\ : Odrv4
    port map (
            O => \N__33895\,
            I => measured_delay_hc_15
        );

    \I__6767\ : LocalMux
    port map (
            O => \N__33892\,
            I => measured_delay_hc_15
        );

    \I__6766\ : LocalMux
    port map (
            O => \N__33887\,
            I => measured_delay_hc_15
        );

    \I__6765\ : InMux
    port map (
            O => \N__33878\,
            I => \N__33873\
        );

    \I__6764\ : InMux
    port map (
            O => \N__33877\,
            I => \N__33870\
        );

    \I__6763\ : CascadeMux
    port map (
            O => \N__33876\,
            I => \N__33867\
        );

    \I__6762\ : LocalMux
    port map (
            O => \N__33873\,
            I => \N__33863\
        );

    \I__6761\ : LocalMux
    port map (
            O => \N__33870\,
            I => \N__33860\
        );

    \I__6760\ : InMux
    port map (
            O => \N__33867\,
            I => \N__33857\
        );

    \I__6759\ : CascadeMux
    port map (
            O => \N__33866\,
            I => \N__33854\
        );

    \I__6758\ : Span4Mux_v
    port map (
            O => \N__33863\,
            I => \N__33850\
        );

    \I__6757\ : Span4Mux_v
    port map (
            O => \N__33860\,
            I => \N__33845\
        );

    \I__6756\ : LocalMux
    port map (
            O => \N__33857\,
            I => \N__33845\
        );

    \I__6755\ : InMux
    port map (
            O => \N__33854\,
            I => \N__33840\
        );

    \I__6754\ : InMux
    port map (
            O => \N__33853\,
            I => \N__33840\
        );

    \I__6753\ : Odrv4
    port map (
            O => \N__33850\,
            I => measured_delay_hc_14
        );

    \I__6752\ : Odrv4
    port map (
            O => \N__33845\,
            I => measured_delay_hc_14
        );

    \I__6751\ : LocalMux
    port map (
            O => \N__33840\,
            I => measured_delay_hc_14
        );

    \I__6750\ : InMux
    port map (
            O => \N__33833\,
            I => \N__33827\
        );

    \I__6749\ : InMux
    port map (
            O => \N__33832\,
            I => \N__33827\
        );

    \I__6748\ : LocalMux
    port map (
            O => \N__33827\,
            I => \N__33823\
        );

    \I__6747\ : InMux
    port map (
            O => \N__33826\,
            I => \N__33820\
        );

    \I__6746\ : Span4Mux_h
    port map (
            O => \N__33823\,
            I => \N__33817\
        );

    \I__6745\ : LocalMux
    port map (
            O => \N__33820\,
            I => \delay_measurement_inst.tr_stateZ0Z_0\
        );

    \I__6744\ : Odrv4
    port map (
            O => \N__33817\,
            I => \delay_measurement_inst.tr_stateZ0Z_0\
        );

    \I__6743\ : InMux
    port map (
            O => \N__33812\,
            I => \N__33809\
        );

    \I__6742\ : LocalMux
    port map (
            O => \N__33809\,
            I => \N__33806\
        );

    \I__6741\ : Span4Mux_v
    port map (
            O => \N__33806\,
            I => \N__33801\
        );

    \I__6740\ : InMux
    port map (
            O => \N__33805\,
            I => \N__33796\
        );

    \I__6739\ : InMux
    port map (
            O => \N__33804\,
            I => \N__33796\
        );

    \I__6738\ : Odrv4
    port map (
            O => \N__33801\,
            I => \delay_measurement_inst.prev_tr_sigZ0\
        );

    \I__6737\ : LocalMux
    port map (
            O => \N__33796\,
            I => \delay_measurement_inst.prev_tr_sigZ0\
        );

    \I__6736\ : CascadeMux
    port map (
            O => \N__33791\,
            I => \delay_measurement_inst.tr_state_RNIMR6LZ0Z_0_cascade_\
        );

    \I__6735\ : InMux
    port map (
            O => \N__33788\,
            I => \N__33784\
        );

    \I__6734\ : CascadeMux
    port map (
            O => \N__33787\,
            I => \N__33780\
        );

    \I__6733\ : LocalMux
    port map (
            O => \N__33784\,
            I => \N__33777\
        );

    \I__6732\ : CascadeMux
    port map (
            O => \N__33783\,
            I => \N__33774\
        );

    \I__6731\ : InMux
    port map (
            O => \N__33780\,
            I => \N__33770\
        );

    \I__6730\ : Span4Mux_v
    port map (
            O => \N__33777\,
            I => \N__33767\
        );

    \I__6729\ : InMux
    port map (
            O => \N__33774\,
            I => \N__33762\
        );

    \I__6728\ : InMux
    port map (
            O => \N__33773\,
            I => \N__33762\
        );

    \I__6727\ : LocalMux
    port map (
            O => \N__33770\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__6726\ : Odrv4
    port map (
            O => \N__33767\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__6725\ : LocalMux
    port map (
            O => \N__33762\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__6724\ : InMux
    port map (
            O => \N__33755\,
            I => \N__33752\
        );

    \I__6723\ : LocalMux
    port map (
            O => \N__33752\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_8\
        );

    \I__6722\ : InMux
    port map (
            O => \N__33749\,
            I => \N__33746\
        );

    \I__6721\ : LocalMux
    port map (
            O => \N__33746\,
            I => \N__33743\
        );

    \I__6720\ : Odrv4
    port map (
            O => \N__33743\,
            I => \current_shift_inst.un4_control_input_axb_8\
        );

    \I__6719\ : InMux
    port map (
            O => \N__33740\,
            I => \N__33737\
        );

    \I__6718\ : LocalMux
    port map (
            O => \N__33737\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_23\
        );

    \I__6717\ : InMux
    port map (
            O => \N__33734\,
            I => \N__33731\
        );

    \I__6716\ : LocalMux
    port map (
            O => \N__33731\,
            I => \N__33728\
        );

    \I__6715\ : Span4Mux_h
    port map (
            O => \N__33728\,
            I => \N__33725\
        );

    \I__6714\ : Odrv4
    port map (
            O => \N__33725\,
            I => \current_shift_inst.un4_control_input_axb_23\
        );

    \I__6713\ : CascadeMux
    port map (
            O => \N__33722\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto13_3Z0Z_1_cascade_\
        );

    \I__6712\ : InMux
    port map (
            O => \N__33719\,
            I => \N__33716\
        );

    \I__6711\ : LocalMux
    port map (
            O => \N__33716\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto13\
        );

    \I__6710\ : InMux
    port map (
            O => \N__33713\,
            I => \N__33704\
        );

    \I__6709\ : InMux
    port map (
            O => \N__33712\,
            I => \N__33704\
        );

    \I__6708\ : InMux
    port map (
            O => \N__33711\,
            I => \N__33704\
        );

    \I__6707\ : LocalMux
    port map (
            O => \N__33704\,
            I => measured_delay_hc_20
        );

    \I__6706\ : CascadeMux
    port map (
            O => \N__33701\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto30_2_cascade_\
        );

    \I__6705\ : InMux
    port map (
            O => \N__33698\,
            I => \N__33695\
        );

    \I__6704\ : LocalMux
    port map (
            O => \N__33695\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt15\
        );

    \I__6703\ : InMux
    port map (
            O => \N__33692\,
            I => \N__33688\
        );

    \I__6702\ : InMux
    port map (
            O => \N__33691\,
            I => \N__33685\
        );

    \I__6701\ : LocalMux
    port map (
            O => \N__33688\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1\
        );

    \I__6700\ : LocalMux
    port map (
            O => \N__33685\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1\
        );

    \I__6699\ : InMux
    port map (
            O => \N__33680\,
            I => \N__33677\
        );

    \I__6698\ : LocalMux
    port map (
            O => \N__33677\,
            I => \N__33674\
        );

    \I__6697\ : Odrv4
    port map (
            O => \N__33674\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_2_tz\
        );

    \I__6696\ : CascadeMux
    port map (
            O => \N__33671\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a1_1_cascade_\
        );

    \I__6695\ : InMux
    port map (
            O => \N__33668\,
            I => \N__33665\
        );

    \I__6694\ : LocalMux
    port map (
            O => \N__33665\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_0\
        );

    \I__6693\ : CascadeMux
    port map (
            O => \N__33662\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_1_cascade_\
        );

    \I__6692\ : CascadeMux
    port map (
            O => \N__33659\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2_cascade_\
        );

    \I__6691\ : InMux
    port map (
            O => \N__33656\,
            I => \N__33653\
        );

    \I__6690\ : LocalMux
    port map (
            O => \N__33653\,
            I => \N__33650\
        );

    \I__6689\ : Odrv4
    port map (
            O => \N__33650\,
            I => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2\
        );

    \I__6688\ : InMux
    port map (
            O => \N__33647\,
            I => \N__33641\
        );

    \I__6687\ : InMux
    port map (
            O => \N__33646\,
            I => \N__33641\
        );

    \I__6686\ : LocalMux
    port map (
            O => \N__33641\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8\
        );

    \I__6685\ : CascadeMux
    port map (
            O => \N__33638\,
            I => \N__33635\
        );

    \I__6684\ : InMux
    port map (
            O => \N__33635\,
            I => \N__33632\
        );

    \I__6683\ : LocalMux
    port map (
            O => \N__33632\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_1\
        );

    \I__6682\ : InMux
    port map (
            O => \N__33629\,
            I => \N__33623\
        );

    \I__6681\ : InMux
    port map (
            O => \N__33628\,
            I => \N__33623\
        );

    \I__6680\ : LocalMux
    port map (
            O => \N__33623\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt30\
        );

    \I__6679\ : InMux
    port map (
            O => \N__33620\,
            I => \N__33617\
        );

    \I__6678\ : LocalMux
    port map (
            O => \N__33617\,
            I => \N__33614\
        );

    \I__6677\ : Odrv4
    port map (
            O => \N__33614\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9\
        );

    \I__6676\ : InMux
    port map (
            O => \N__33611\,
            I => \N__33608\
        );

    \I__6675\ : LocalMux
    port map (
            O => \N__33608\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0\
        );

    \I__6674\ : CascadeMux
    port map (
            O => \N__33605\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0_cascade_\
        );

    \I__6673\ : CascadeMux
    port map (
            O => \N__33602\,
            I => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1_cascade_\
        );

    \I__6672\ : InMux
    port map (
            O => \N__33599\,
            I => \N__33596\
        );

    \I__6671\ : LocalMux
    port map (
            O => \N__33596\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt30_0\
        );

    \I__6670\ : InMux
    port map (
            O => \N__33593\,
            I => \N__33586\
        );

    \I__6669\ : InMux
    port map (
            O => \N__33592\,
            I => \N__33586\
        );

    \I__6668\ : InMux
    port map (
            O => \N__33591\,
            I => \N__33582\
        );

    \I__6667\ : LocalMux
    port map (
            O => \N__33586\,
            I => \N__33579\
        );

    \I__6666\ : InMux
    port map (
            O => \N__33585\,
            I => \N__33576\
        );

    \I__6665\ : LocalMux
    port map (
            O => \N__33582\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__6664\ : Odrv12
    port map (
            O => \N__33579\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__6663\ : LocalMux
    port map (
            O => \N__33576\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__6662\ : InMux
    port map (
            O => \N__33569\,
            I => \N__33566\
        );

    \I__6661\ : LocalMux
    port map (
            O => \N__33566\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8\
        );

    \I__6660\ : CascadeMux
    port map (
            O => \N__33563\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_2_cascade_\
        );

    \I__6659\ : InMux
    port map (
            O => \N__33560\,
            I => \N__33557\
        );

    \I__6658\ : LocalMux
    port map (
            O => \N__33557\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_11\
        );

    \I__6657\ : InMux
    port map (
            O => \N__33554\,
            I => \N__33550\
        );

    \I__6656\ : InMux
    port map (
            O => \N__33553\,
            I => \N__33547\
        );

    \I__6655\ : LocalMux
    port map (
            O => \N__33550\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_1\
        );

    \I__6654\ : LocalMux
    port map (
            O => \N__33547\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_1\
        );

    \I__6653\ : InMux
    port map (
            O => \N__33542\,
            I => \N__33538\
        );

    \I__6652\ : InMux
    port map (
            O => \N__33541\,
            I => \N__33535\
        );

    \I__6651\ : LocalMux
    port map (
            O => \N__33538\,
            I => \N__33530\
        );

    \I__6650\ : LocalMux
    port map (
            O => \N__33535\,
            I => \N__33530\
        );

    \I__6649\ : Sp12to4
    port map (
            O => \N__33530\,
            I => \N__33526\
        );

    \I__6648\ : InMux
    port map (
            O => \N__33529\,
            I => \N__33523\
        );

    \I__6647\ : Span12Mux_v
    port map (
            O => \N__33526\,
            I => \N__33520\
        );

    \I__6646\ : LocalMux
    port map (
            O => \N__33523\,
            I => \current_shift_inst.start_timer_phaseZ0\
        );

    \I__6645\ : Odrv12
    port map (
            O => \N__33520\,
            I => \current_shift_inst.start_timer_phaseZ0\
        );

    \I__6644\ : InMux
    port map (
            O => \N__33515\,
            I => \N__33509\
        );

    \I__6643\ : InMux
    port map (
            O => \N__33514\,
            I => \N__33506\
        );

    \I__6642\ : InMux
    port map (
            O => \N__33513\,
            I => \N__33503\
        );

    \I__6641\ : InMux
    port map (
            O => \N__33512\,
            I => \N__33500\
        );

    \I__6640\ : LocalMux
    port map (
            O => \N__33509\,
            I => \current_shift_inst.timer_phase.runningZ0\
        );

    \I__6639\ : LocalMux
    port map (
            O => \N__33506\,
            I => \current_shift_inst.timer_phase.runningZ0\
        );

    \I__6638\ : LocalMux
    port map (
            O => \N__33503\,
            I => \current_shift_inst.timer_phase.runningZ0\
        );

    \I__6637\ : LocalMux
    port map (
            O => \N__33500\,
            I => \current_shift_inst.timer_phase.runningZ0\
        );

    \I__6636\ : InMux
    port map (
            O => \N__33491\,
            I => \N__33486\
        );

    \I__6635\ : InMux
    port map (
            O => \N__33490\,
            I => \N__33483\
        );

    \I__6634\ : InMux
    port map (
            O => \N__33489\,
            I => \N__33479\
        );

    \I__6633\ : LocalMux
    port map (
            O => \N__33486\,
            I => \N__33476\
        );

    \I__6632\ : LocalMux
    port map (
            O => \N__33483\,
            I => \N__33473\
        );

    \I__6631\ : CascadeMux
    port map (
            O => \N__33482\,
            I => \N__33470\
        );

    \I__6630\ : LocalMux
    port map (
            O => \N__33479\,
            I => \N__33463\
        );

    \I__6629\ : Sp12to4
    port map (
            O => \N__33476\,
            I => \N__33463\
        );

    \I__6628\ : Span12Mux_s4_v
    port map (
            O => \N__33473\,
            I => \N__33463\
        );

    \I__6627\ : InMux
    port map (
            O => \N__33470\,
            I => \N__33460\
        );

    \I__6626\ : Span12Mux_v
    port map (
            O => \N__33463\,
            I => \N__33457\
        );

    \I__6625\ : LocalMux
    port map (
            O => \N__33460\,
            I => \current_shift_inst.stop_timer_phaseZ0\
        );

    \I__6624\ : Odrv12
    port map (
            O => \N__33457\,
            I => \current_shift_inst.stop_timer_phaseZ0\
        );

    \I__6623\ : IoInMux
    port map (
            O => \N__33452\,
            I => \N__33449\
        );

    \I__6622\ : LocalMux
    port map (
            O => \N__33449\,
            I => \N__33446\
        );

    \I__6621\ : Odrv12
    port map (
            O => \N__33446\,
            I => \current_shift_inst.timer_phase.N_188_i\
        );

    \I__6620\ : IoInMux
    port map (
            O => \N__33443\,
            I => \N__33440\
        );

    \I__6619\ : LocalMux
    port map (
            O => \N__33440\,
            I => \N__33437\
        );

    \I__6618\ : Odrv4
    port map (
            O => \N__33437\,
            I => s2_phy_c
        );

    \I__6617\ : CascadeMux
    port map (
            O => \N__33434\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_3_cascade_\
        );

    \I__6616\ : InMux
    port map (
            O => \N__33431\,
            I => \N__33428\
        );

    \I__6615\ : LocalMux
    port map (
            O => \N__33428\,
            I => \N__33423\
        );

    \I__6614\ : InMux
    port map (
            O => \N__33427\,
            I => \N__33420\
        );

    \I__6613\ : InMux
    port map (
            O => \N__33426\,
            I => \N__33417\
        );

    \I__6612\ : Span4Mux_v
    port map (
            O => \N__33423\,
            I => \N__33412\
        );

    \I__6611\ : LocalMux
    port map (
            O => \N__33420\,
            I => \N__33412\
        );

    \I__6610\ : LocalMux
    port map (
            O => \N__33417\,
            I => \N__33409\
        );

    \I__6609\ : Odrv4
    port map (
            O => \N__33412\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__6608\ : Odrv12
    port map (
            O => \N__33409\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__6607\ : CascadeMux
    port map (
            O => \N__33404\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt14_cascade_\
        );

    \I__6606\ : InMux
    port map (
            O => \N__33401\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9\
        );

    \I__6605\ : InMux
    port map (
            O => \N__33398\,
            I => \N__33395\
        );

    \I__6604\ : LocalMux
    port map (
            O => \N__33395\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12\
        );

    \I__6603\ : InMux
    port map (
            O => \N__33392\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10\
        );

    \I__6602\ : InMux
    port map (
            O => \N__33389\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11\
        );

    \I__6601\ : InMux
    port map (
            O => \N__33386\,
            I => \N__33383\
        );

    \I__6600\ : LocalMux
    port map (
            O => \N__33383\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14\
        );

    \I__6599\ : InMux
    port map (
            O => \N__33380\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12\
        );

    \I__6598\ : InMux
    port map (
            O => \N__33377\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13\
        );

    \I__6597\ : InMux
    port map (
            O => \N__33374\,
            I => \N__33371\
        );

    \I__6596\ : LocalMux
    port map (
            O => \N__33371\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16\
        );

    \I__6595\ : InMux
    port map (
            O => \N__33368\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14\
        );

    \I__6594\ : InMux
    port map (
            O => \N__33365\,
            I => \bfn_13_25_0_\
        );

    \I__6593\ : InMux
    port map (
            O => \N__33362\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16\
        );

    \I__6592\ : InMux
    port map (
            O => \N__33359\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17\
        );

    \I__6591\ : InMux
    port map (
            O => \N__33356\,
            I => \N__33353\
        );

    \I__6590\ : LocalMux
    port map (
            O => \N__33353\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19\
        );

    \I__6589\ : InMux
    port map (
            O => \N__33350\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0\
        );

    \I__6588\ : InMux
    port map (
            O => \N__33347\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1\
        );

    \I__6587\ : InMux
    port map (
            O => \N__33344\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2\
        );

    \I__6586\ : InMux
    port map (
            O => \N__33341\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3\
        );

    \I__6585\ : InMux
    port map (
            O => \N__33338\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4\
        );

    \I__6584\ : InMux
    port map (
            O => \N__33335\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5\
        );

    \I__6583\ : InMux
    port map (
            O => \N__33332\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6\
        );

    \I__6582\ : InMux
    port map (
            O => \N__33329\,
            I => \bfn_13_24_0_\
        );

    \I__6581\ : InMux
    port map (
            O => \N__33326\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8\
        );

    \I__6580\ : CascadeMux
    port map (
            O => \N__33323\,
            I => \N__33320\
        );

    \I__6579\ : InMux
    port map (
            O => \N__33320\,
            I => \N__33317\
        );

    \I__6578\ : LocalMux
    port map (
            O => \N__33317\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_18\
        );

    \I__6577\ : CascadeMux
    port map (
            O => \N__33314\,
            I => \N__33311\
        );

    \I__6576\ : InMux
    port map (
            O => \N__33311\,
            I => \N__33308\
        );

    \I__6575\ : LocalMux
    port map (
            O => \N__33308\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_19\
        );

    \I__6574\ : InMux
    port map (
            O => \N__33305\,
            I => \N__33298\
        );

    \I__6573\ : InMux
    port map (
            O => \N__33304\,
            I => \N__33298\
        );

    \I__6572\ : InMux
    port map (
            O => \N__33303\,
            I => \N__33295\
        );

    \I__6571\ : LocalMux
    port map (
            O => \N__33298\,
            I => \phase_controller_slave.stateZ0Z_0\
        );

    \I__6570\ : LocalMux
    port map (
            O => \N__33295\,
            I => \phase_controller_slave.stateZ0Z_0\
        );

    \I__6569\ : CascadeMux
    port map (
            O => \N__33290\,
            I => \N__33284\
        );

    \I__6568\ : InMux
    port map (
            O => \N__33289\,
            I => \N__33281\
        );

    \I__6567\ : InMux
    port map (
            O => \N__33288\,
            I => \N__33278\
        );

    \I__6566\ : InMux
    port map (
            O => \N__33287\,
            I => \N__33273\
        );

    \I__6565\ : InMux
    port map (
            O => \N__33284\,
            I => \N__33273\
        );

    \I__6564\ : LocalMux
    port map (
            O => \N__33281\,
            I => \phase_controller_slave.stateZ0Z_4\
        );

    \I__6563\ : LocalMux
    port map (
            O => \N__33278\,
            I => \phase_controller_slave.stateZ0Z_4\
        );

    \I__6562\ : LocalMux
    port map (
            O => \N__33273\,
            I => \phase_controller_slave.stateZ0Z_4\
        );

    \I__6561\ : InMux
    port map (
            O => \N__33266\,
            I => \N__33263\
        );

    \I__6560\ : LocalMux
    port map (
            O => \N__33263\,
            I => \N__33260\
        );

    \I__6559\ : Span4Mux_v
    port map (
            O => \N__33260\,
            I => \N__33257\
        );

    \I__6558\ : Odrv4
    port map (
            O => \N__33257\,
            I => \phase_controller_slave.start_timer_tr_0_sqmuxa\
        );

    \I__6557\ : CascadeMux
    port map (
            O => \N__33254\,
            I => \phase_controller_slave.N_210_cascade_\
        );

    \I__6556\ : CascadeMux
    port map (
            O => \N__33251\,
            I => \phase_controller_slave.stoper_tr.time_passed11_cascade_\
        );

    \I__6555\ : CascadeMux
    port map (
            O => \N__33248\,
            I => \N__33244\
        );

    \I__6554\ : InMux
    port map (
            O => \N__33247\,
            I => \N__33239\
        );

    \I__6553\ : InMux
    port map (
            O => \N__33244\,
            I => \N__33236\
        );

    \I__6552\ : InMux
    port map (
            O => \N__33243\,
            I => \N__33231\
        );

    \I__6551\ : InMux
    port map (
            O => \N__33242\,
            I => \N__33231\
        );

    \I__6550\ : LocalMux
    port map (
            O => \N__33239\,
            I => \phase_controller_slave.tr_time_passed\
        );

    \I__6549\ : LocalMux
    port map (
            O => \N__33236\,
            I => \phase_controller_slave.tr_time_passed\
        );

    \I__6548\ : LocalMux
    port map (
            O => \N__33231\,
            I => \phase_controller_slave.tr_time_passed\
        );

    \I__6547\ : InMux
    port map (
            O => \N__33224\,
            I => \N__33221\
        );

    \I__6546\ : LocalMux
    port map (
            O => \N__33221\,
            I => \phase_controller_slave.stoper_tr.time_passed_1_sqmuxa\
        );

    \I__6545\ : CascadeMux
    port map (
            O => \N__33218\,
            I => \N__33215\
        );

    \I__6544\ : InMux
    port map (
            O => \N__33215\,
            I => \N__33212\
        );

    \I__6543\ : LocalMux
    port map (
            O => \N__33212\,
            I => \N__33209\
        );

    \I__6542\ : Span4Mux_h
    port map (
            O => \N__33209\,
            I => \N__33206\
        );

    \I__6541\ : Odrv4
    port map (
            O => \N__33206\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_14\
        );

    \I__6540\ : InMux
    port map (
            O => \N__33203\,
            I => \N__33200\
        );

    \I__6539\ : LocalMux
    port map (
            O => \N__33200\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_14\
        );

    \I__6538\ : CascadeMux
    port map (
            O => \N__33197\,
            I => \N__33194\
        );

    \I__6537\ : InMux
    port map (
            O => \N__33194\,
            I => \N__33191\
        );

    \I__6536\ : LocalMux
    port map (
            O => \N__33191\,
            I => \N__33188\
        );

    \I__6535\ : Span4Mux_v
    port map (
            O => \N__33188\,
            I => \N__33185\
        );

    \I__6534\ : Span4Mux_v
    port map (
            O => \N__33185\,
            I => \N__33182\
        );

    \I__6533\ : Odrv4
    port map (
            O => \N__33182\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_15\
        );

    \I__6532\ : InMux
    port map (
            O => \N__33179\,
            I => \N__33176\
        );

    \I__6531\ : LocalMux
    port map (
            O => \N__33176\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_15\
        );

    \I__6530\ : InMux
    port map (
            O => \N__33173\,
            I => \N__33170\
        );

    \I__6529\ : LocalMux
    port map (
            O => \N__33170\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_16\
        );

    \I__6528\ : InMux
    port map (
            O => \N__33167\,
            I => \N__33164\
        );

    \I__6527\ : LocalMux
    port map (
            O => \N__33164\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_17\
        );

    \I__6526\ : InMux
    port map (
            O => \N__33161\,
            I => \N__33158\
        );

    \I__6525\ : LocalMux
    port map (
            O => \N__33158\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_18\
        );

    \I__6524\ : InMux
    port map (
            O => \N__33155\,
            I => \N__33152\
        );

    \I__6523\ : LocalMux
    port map (
            O => \N__33152\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_19\
        );

    \I__6522\ : InMux
    port map (
            O => \N__33149\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__6521\ : CascadeMux
    port map (
            O => \N__33146\,
            I => \N__33143\
        );

    \I__6520\ : InMux
    port map (
            O => \N__33143\,
            I => \N__33140\
        );

    \I__6519\ : LocalMux
    port map (
            O => \N__33140\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_17\
        );

    \I__6518\ : CascadeMux
    port map (
            O => \N__33137\,
            I => \N__33134\
        );

    \I__6517\ : InMux
    port map (
            O => \N__33134\,
            I => \N__33131\
        );

    \I__6516\ : LocalMux
    port map (
            O => \N__33131\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_6\
        );

    \I__6515\ : InMux
    port map (
            O => \N__33128\,
            I => \N__33125\
        );

    \I__6514\ : LocalMux
    port map (
            O => \N__33125\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_6\
        );

    \I__6513\ : CascadeMux
    port map (
            O => \N__33122\,
            I => \N__33119\
        );

    \I__6512\ : InMux
    port map (
            O => \N__33119\,
            I => \N__33116\
        );

    \I__6511\ : LocalMux
    port map (
            O => \N__33116\,
            I => \N__33113\
        );

    \I__6510\ : Odrv4
    port map (
            O => \N__33113\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_7\
        );

    \I__6509\ : InMux
    port map (
            O => \N__33110\,
            I => \N__33107\
        );

    \I__6508\ : LocalMux
    port map (
            O => \N__33107\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_7\
        );

    \I__6507\ : CascadeMux
    port map (
            O => \N__33104\,
            I => \N__33101\
        );

    \I__6506\ : InMux
    port map (
            O => \N__33101\,
            I => \N__33098\
        );

    \I__6505\ : LocalMux
    port map (
            O => \N__33098\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_8\
        );

    \I__6504\ : InMux
    port map (
            O => \N__33095\,
            I => \N__33092\
        );

    \I__6503\ : LocalMux
    port map (
            O => \N__33092\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_8\
        );

    \I__6502\ : CascadeMux
    port map (
            O => \N__33089\,
            I => \N__33086\
        );

    \I__6501\ : InMux
    port map (
            O => \N__33086\,
            I => \N__33083\
        );

    \I__6500\ : LocalMux
    port map (
            O => \N__33083\,
            I => \N__33080\
        );

    \I__6499\ : Odrv4
    port map (
            O => \N__33080\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_9\
        );

    \I__6498\ : InMux
    port map (
            O => \N__33077\,
            I => \N__33074\
        );

    \I__6497\ : LocalMux
    port map (
            O => \N__33074\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_9\
        );

    \I__6496\ : CascadeMux
    port map (
            O => \N__33071\,
            I => \N__33068\
        );

    \I__6495\ : InMux
    port map (
            O => \N__33068\,
            I => \N__33065\
        );

    \I__6494\ : LocalMux
    port map (
            O => \N__33065\,
            I => \N__33062\
        );

    \I__6493\ : Span12Mux_h
    port map (
            O => \N__33062\,
            I => \N__33059\
        );

    \I__6492\ : Odrv12
    port map (
            O => \N__33059\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_10\
        );

    \I__6491\ : InMux
    port map (
            O => \N__33056\,
            I => \N__33053\
        );

    \I__6490\ : LocalMux
    port map (
            O => \N__33053\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_10\
        );

    \I__6489\ : CascadeMux
    port map (
            O => \N__33050\,
            I => \N__33047\
        );

    \I__6488\ : InMux
    port map (
            O => \N__33047\,
            I => \N__33044\
        );

    \I__6487\ : LocalMux
    port map (
            O => \N__33044\,
            I => \N__33041\
        );

    \I__6486\ : Span4Mux_v
    port map (
            O => \N__33041\,
            I => \N__33038\
        );

    \I__6485\ : Span4Mux_v
    port map (
            O => \N__33038\,
            I => \N__33035\
        );

    \I__6484\ : Odrv4
    port map (
            O => \N__33035\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_11\
        );

    \I__6483\ : InMux
    port map (
            O => \N__33032\,
            I => \N__33029\
        );

    \I__6482\ : LocalMux
    port map (
            O => \N__33029\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_11\
        );

    \I__6481\ : CascadeMux
    port map (
            O => \N__33026\,
            I => \N__33023\
        );

    \I__6480\ : InMux
    port map (
            O => \N__33023\,
            I => \N__33020\
        );

    \I__6479\ : LocalMux
    port map (
            O => \N__33020\,
            I => \N__33017\
        );

    \I__6478\ : Span4Mux_v
    port map (
            O => \N__33017\,
            I => \N__33014\
        );

    \I__6477\ : Span4Mux_v
    port map (
            O => \N__33014\,
            I => \N__33011\
        );

    \I__6476\ : Odrv4
    port map (
            O => \N__33011\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_12\
        );

    \I__6475\ : InMux
    port map (
            O => \N__33008\,
            I => \N__33005\
        );

    \I__6474\ : LocalMux
    port map (
            O => \N__33005\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_12\
        );

    \I__6473\ : CascadeMux
    port map (
            O => \N__33002\,
            I => \N__32999\
        );

    \I__6472\ : InMux
    port map (
            O => \N__32999\,
            I => \N__32996\
        );

    \I__6471\ : LocalMux
    port map (
            O => \N__32996\,
            I => \N__32993\
        );

    \I__6470\ : Span4Mux_v
    port map (
            O => \N__32993\,
            I => \N__32990\
        );

    \I__6469\ : Span4Mux_v
    port map (
            O => \N__32990\,
            I => \N__32987\
        );

    \I__6468\ : Odrv4
    port map (
            O => \N__32987\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_13\
        );

    \I__6467\ : InMux
    port map (
            O => \N__32984\,
            I => \N__32981\
        );

    \I__6466\ : LocalMux
    port map (
            O => \N__32981\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_13\
        );

    \I__6465\ : CascadeMux
    port map (
            O => \N__32978\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6_cascade_\
        );

    \I__6464\ : CascadeMux
    port map (
            O => \N__32975\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13_cascade_\
        );

    \I__6463\ : CascadeMux
    port map (
            O => \N__32972\,
            I => \N__32969\
        );

    \I__6462\ : InMux
    port map (
            O => \N__32969\,
            I => \N__32966\
        );

    \I__6461\ : LocalMux
    port map (
            O => \N__32966\,
            I => \N__32963\
        );

    \I__6460\ : Odrv4
    port map (
            O => \N__32963\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_1\
        );

    \I__6459\ : InMux
    port map (
            O => \N__32960\,
            I => \N__32957\
        );

    \I__6458\ : LocalMux
    port map (
            O => \N__32957\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_1\
        );

    \I__6457\ : CascadeMux
    port map (
            O => \N__32954\,
            I => \N__32951\
        );

    \I__6456\ : InMux
    port map (
            O => \N__32951\,
            I => \N__32948\
        );

    \I__6455\ : LocalMux
    port map (
            O => \N__32948\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_2\
        );

    \I__6454\ : InMux
    port map (
            O => \N__32945\,
            I => \N__32942\
        );

    \I__6453\ : LocalMux
    port map (
            O => \N__32942\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_2\
        );

    \I__6452\ : CascadeMux
    port map (
            O => \N__32939\,
            I => \N__32936\
        );

    \I__6451\ : InMux
    port map (
            O => \N__32936\,
            I => \N__32933\
        );

    \I__6450\ : LocalMux
    port map (
            O => \N__32933\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_3\
        );

    \I__6449\ : InMux
    port map (
            O => \N__32930\,
            I => \N__32927\
        );

    \I__6448\ : LocalMux
    port map (
            O => \N__32927\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_3\
        );

    \I__6447\ : CascadeMux
    port map (
            O => \N__32924\,
            I => \N__32921\
        );

    \I__6446\ : InMux
    port map (
            O => \N__32921\,
            I => \N__32918\
        );

    \I__6445\ : LocalMux
    port map (
            O => \N__32918\,
            I => \N__32915\
        );

    \I__6444\ : Odrv4
    port map (
            O => \N__32915\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_4\
        );

    \I__6443\ : InMux
    port map (
            O => \N__32912\,
            I => \N__32909\
        );

    \I__6442\ : LocalMux
    port map (
            O => \N__32909\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_4\
        );

    \I__6441\ : CascadeMux
    port map (
            O => \N__32906\,
            I => \N__32903\
        );

    \I__6440\ : InMux
    port map (
            O => \N__32903\,
            I => \N__32900\
        );

    \I__6439\ : LocalMux
    port map (
            O => \N__32900\,
            I => \N__32897\
        );

    \I__6438\ : Odrv12
    port map (
            O => \N__32897\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_5\
        );

    \I__6437\ : InMux
    port map (
            O => \N__32894\,
            I => \N__32891\
        );

    \I__6436\ : LocalMux
    port map (
            O => \N__32891\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_5\
        );

    \I__6435\ : IoInMux
    port map (
            O => \N__32888\,
            I => \N__32885\
        );

    \I__6434\ : LocalMux
    port map (
            O => \N__32885\,
            I => \N__32882\
        );

    \I__6433\ : IoSpan4Mux
    port map (
            O => \N__32882\,
            I => \N__32879\
        );

    \I__6432\ : Span4Mux_s3_v
    port map (
            O => \N__32879\,
            I => \N__32876\
        );

    \I__6431\ : Span4Mux_v
    port map (
            O => \N__32876\,
            I => \N__32872\
        );

    \I__6430\ : InMux
    port map (
            O => \N__32875\,
            I => \N__32869\
        );

    \I__6429\ : Span4Mux_v
    port map (
            O => \N__32872\,
            I => \N__32866\
        );

    \I__6428\ : LocalMux
    port map (
            O => \N__32869\,
            I => \N__32863\
        );

    \I__6427\ : Span4Mux_v
    port map (
            O => \N__32866\,
            I => \N__32858\
        );

    \I__6426\ : Span4Mux_v
    port map (
            O => \N__32863\,
            I => \N__32858\
        );

    \I__6425\ : Odrv4
    port map (
            O => \N__32858\,
            I => s1_phy_c
        );

    \I__6424\ : InMux
    port map (
            O => \N__32855\,
            I => \N__32852\
        );

    \I__6423\ : LocalMux
    port map (
            O => \N__32852\,
            I => \current_shift_inst.S1_syncZ0Z0\
        );

    \I__6422\ : InMux
    port map (
            O => \N__32849\,
            I => \N__32846\
        );

    \I__6421\ : LocalMux
    port map (
            O => \N__32846\,
            I => \current_shift_inst.S3_sync_prevZ0\
        );

    \I__6420\ : InMux
    port map (
            O => \N__32843\,
            I => \N__32839\
        );

    \I__6419\ : CascadeMux
    port map (
            O => \N__32842\,
            I => \N__32835\
        );

    \I__6418\ : LocalMux
    port map (
            O => \N__32839\,
            I => \N__32832\
        );

    \I__6417\ : InMux
    port map (
            O => \N__32838\,
            I => \N__32827\
        );

    \I__6416\ : InMux
    port map (
            O => \N__32835\,
            I => \N__32827\
        );

    \I__6415\ : Span4Mux_h
    port map (
            O => \N__32832\,
            I => \N__32822\
        );

    \I__6414\ : LocalMux
    port map (
            O => \N__32827\,
            I => \N__32822\
        );

    \I__6413\ : Sp12to4
    port map (
            O => \N__32822\,
            I => \N__32819\
        );

    \I__6412\ : Odrv12
    port map (
            O => \N__32819\,
            I => \current_shift_inst.S3_riseZ0\
        );

    \I__6411\ : InMux
    port map (
            O => \N__32816\,
            I => \N__32810\
        );

    \I__6410\ : InMux
    port map (
            O => \N__32815\,
            I => \N__32810\
        );

    \I__6409\ : LocalMux
    port map (
            O => \N__32810\,
            I => \current_shift_inst.S1_syncZ0Z1\
        );

    \I__6408\ : InMux
    port map (
            O => \N__32807\,
            I => \N__32804\
        );

    \I__6407\ : LocalMux
    port map (
            O => \N__32804\,
            I => \current_shift_inst.S1_sync_prevZ0\
        );

    \I__6406\ : InMux
    port map (
            O => \N__32801\,
            I => \N__32798\
        );

    \I__6405\ : LocalMux
    port map (
            O => \N__32798\,
            I => \current_shift_inst.S3_syncZ0Z0\
        );

    \I__6404\ : InMux
    port map (
            O => \N__32795\,
            I => \N__32789\
        );

    \I__6403\ : InMux
    port map (
            O => \N__32794\,
            I => \N__32789\
        );

    \I__6402\ : LocalMux
    port map (
            O => \N__32789\,
            I => \current_shift_inst.S3_syncZ0Z1\
        );

    \I__6401\ : InMux
    port map (
            O => \N__32786\,
            I => \N__32783\
        );

    \I__6400\ : LocalMux
    port map (
            O => \N__32783\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_26\
        );

    \I__6399\ : InMux
    port map (
            O => \N__32780\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\
        );

    \I__6398\ : InMux
    port map (
            O => \N__32777\,
            I => \N__32774\
        );

    \I__6397\ : LocalMux
    port map (
            O => \N__32774\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_27\
        );

    \I__6396\ : InMux
    port map (
            O => \N__32771\,
            I => \bfn_13_16_0_\
        );

    \I__6395\ : InMux
    port map (
            O => \N__32768\,
            I => \N__32765\
        );

    \I__6394\ : LocalMux
    port map (
            O => \N__32765\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_28\
        );

    \I__6393\ : InMux
    port map (
            O => \N__32762\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\
        );

    \I__6392\ : InMux
    port map (
            O => \N__32759\,
            I => \N__32756\
        );

    \I__6391\ : LocalMux
    port map (
            O => \N__32756\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_29\
        );

    \I__6390\ : InMux
    port map (
            O => \N__32753\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\
        );

    \I__6389\ : InMux
    port map (
            O => \N__32750\,
            I => \N__32747\
        );

    \I__6388\ : LocalMux
    port map (
            O => \N__32747\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_30\
        );

    \I__6387\ : InMux
    port map (
            O => \N__32744\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\
        );

    \I__6386\ : CEMux
    port map (
            O => \N__32741\,
            I => \N__32726\
        );

    \I__6385\ : CEMux
    port map (
            O => \N__32740\,
            I => \N__32726\
        );

    \I__6384\ : CEMux
    port map (
            O => \N__32739\,
            I => \N__32726\
        );

    \I__6383\ : CEMux
    port map (
            O => \N__32738\,
            I => \N__32726\
        );

    \I__6382\ : CEMux
    port map (
            O => \N__32737\,
            I => \N__32726\
        );

    \I__6381\ : GlobalMux
    port map (
            O => \N__32726\,
            I => \N__32723\
        );

    \I__6380\ : gio2CtrlBuf
    port map (
            O => \N__32723\,
            I => \current_shift_inst.timer_s1.N_187_i_g\
        );

    \I__6379\ : InMux
    port map (
            O => \N__32720\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\
        );

    \I__6378\ : InMux
    port map (
            O => \N__32717\,
            I => \N__32711\
        );

    \I__6377\ : InMux
    port map (
            O => \N__32716\,
            I => \N__32711\
        );

    \I__6376\ : LocalMux
    port map (
            O => \N__32711\,
            I => \N__32708\
        );

    \I__6375\ : Span4Mux_v
    port map (
            O => \N__32708\,
            I => \N__32705\
        );

    \I__6374\ : Odrv4
    port map (
            O => \N__32705\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__6373\ : InMux
    port map (
            O => \N__32702\,
            I => \N__32691\
        );

    \I__6372\ : InMux
    port map (
            O => \N__32701\,
            I => \N__32691\
        );

    \I__6371\ : InMux
    port map (
            O => \N__32700\,
            I => \N__32680\
        );

    \I__6370\ : InMux
    port map (
            O => \N__32699\,
            I => \N__32680\
        );

    \I__6369\ : InMux
    port map (
            O => \N__32698\,
            I => \N__32680\
        );

    \I__6368\ : InMux
    port map (
            O => \N__32697\,
            I => \N__32680\
        );

    \I__6367\ : InMux
    port map (
            O => \N__32696\,
            I => \N__32680\
        );

    \I__6366\ : LocalMux
    port map (
            O => \N__32691\,
            I => \N__32675\
        );

    \I__6365\ : LocalMux
    port map (
            O => \N__32680\,
            I => \N__32675\
        );

    \I__6364\ : Odrv12
    port map (
            O => \N__32675\,
            I => \current_shift_inst.S1_riseZ0\
        );

    \I__6363\ : InMux
    port map (
            O => \N__32672\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\
        );

    \I__6362\ : InMux
    port map (
            O => \N__32669\,
            I => \N__32666\
        );

    \I__6361\ : LocalMux
    port map (
            O => \N__32666\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_18\
        );

    \I__6360\ : InMux
    port map (
            O => \N__32663\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\
        );

    \I__6359\ : InMux
    port map (
            O => \N__32660\,
            I => \N__32657\
        );

    \I__6358\ : LocalMux
    port map (
            O => \N__32657\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_19\
        );

    \I__6357\ : InMux
    port map (
            O => \N__32654\,
            I => \bfn_13_15_0_\
        );

    \I__6356\ : InMux
    port map (
            O => \N__32651\,
            I => \N__32648\
        );

    \I__6355\ : LocalMux
    port map (
            O => \N__32648\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_20\
        );

    \I__6354\ : InMux
    port map (
            O => \N__32645\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\
        );

    \I__6353\ : InMux
    port map (
            O => \N__32642\,
            I => \N__32639\
        );

    \I__6352\ : LocalMux
    port map (
            O => \N__32639\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_21\
        );

    \I__6351\ : InMux
    port map (
            O => \N__32636\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\
        );

    \I__6350\ : InMux
    port map (
            O => \N__32633\,
            I => \N__32630\
        );

    \I__6349\ : LocalMux
    port map (
            O => \N__32630\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_22\
        );

    \I__6348\ : InMux
    port map (
            O => \N__32627\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\
        );

    \I__6347\ : InMux
    port map (
            O => \N__32624\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\
        );

    \I__6346\ : InMux
    port map (
            O => \N__32621\,
            I => \N__32618\
        );

    \I__6345\ : LocalMux
    port map (
            O => \N__32618\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_24\
        );

    \I__6344\ : InMux
    port map (
            O => \N__32615\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\
        );

    \I__6343\ : InMux
    port map (
            O => \N__32612\,
            I => \N__32609\
        );

    \I__6342\ : LocalMux
    port map (
            O => \N__32609\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_25\
        );

    \I__6341\ : InMux
    port map (
            O => \N__32606\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\
        );

    \I__6340\ : InMux
    port map (
            O => \N__32603\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\
        );

    \I__6339\ : InMux
    port map (
            O => \N__32600\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\
        );

    \I__6338\ : InMux
    port map (
            O => \N__32597\,
            I => \N__32594\
        );

    \I__6337\ : LocalMux
    port map (
            O => \N__32594\,
            I => \N__32591\
        );

    \I__6336\ : Odrv4
    port map (
            O => \N__32591\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_10\
        );

    \I__6335\ : InMux
    port map (
            O => \N__32588\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\
        );

    \I__6334\ : InMux
    port map (
            O => \N__32585\,
            I => \N__32582\
        );

    \I__6333\ : LocalMux
    port map (
            O => \N__32582\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_11\
        );

    \I__6332\ : InMux
    port map (
            O => \N__32579\,
            I => \bfn_13_14_0_\
        );

    \I__6331\ : InMux
    port map (
            O => \N__32576\,
            I => \N__32573\
        );

    \I__6330\ : LocalMux
    port map (
            O => \N__32573\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_12\
        );

    \I__6329\ : InMux
    port map (
            O => \N__32570\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\
        );

    \I__6328\ : InMux
    port map (
            O => \N__32567\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\
        );

    \I__6327\ : InMux
    port map (
            O => \N__32564\,
            I => \N__32561\
        );

    \I__6326\ : LocalMux
    port map (
            O => \N__32561\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_14\
        );

    \I__6325\ : InMux
    port map (
            O => \N__32558\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\
        );

    \I__6324\ : InMux
    port map (
            O => \N__32555\,
            I => \N__32552\
        );

    \I__6323\ : LocalMux
    port map (
            O => \N__32552\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_15\
        );

    \I__6322\ : InMux
    port map (
            O => \N__32549\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\
        );

    \I__6321\ : InMux
    port map (
            O => \N__32546\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\
        );

    \I__6320\ : InMux
    port map (
            O => \N__32543\,
            I => \N__32540\
        );

    \I__6319\ : LocalMux
    port map (
            O => \N__32540\,
            I => \N__32535\
        );

    \I__6318\ : InMux
    port map (
            O => \N__32539\,
            I => \N__32532\
        );

    \I__6317\ : InMux
    port map (
            O => \N__32538\,
            I => \N__32529\
        );

    \I__6316\ : Span4Mux_v
    port map (
            O => \N__32535\,
            I => \N__32526\
        );

    \I__6315\ : LocalMux
    port map (
            O => \N__32532\,
            I => \N__32521\
        );

    \I__6314\ : LocalMux
    port map (
            O => \N__32529\,
            I => \N__32521\
        );

    \I__6313\ : Span4Mux_h
    port map (
            O => \N__32526\,
            I => \N__32518\
        );

    \I__6312\ : Span4Mux_v
    port map (
            O => \N__32521\,
            I => \N__32515\
        );

    \I__6311\ : Odrv4
    port map (
            O => \N__32518\,
            I => \il_max_comp1_D2\
        );

    \I__6310\ : Odrv4
    port map (
            O => \N__32515\,
            I => \il_max_comp1_D2\
        );

    \I__6309\ : CascadeMux
    port map (
            O => \N__32510\,
            I => \phase_controller_inst1.N_86_cascade_\
        );

    \I__6308\ : InMux
    port map (
            O => \N__32507\,
            I => \N__32499\
        );

    \I__6307\ : InMux
    port map (
            O => \N__32506\,
            I => \N__32499\
        );

    \I__6306\ : InMux
    port map (
            O => \N__32505\,
            I => \N__32496\
        );

    \I__6305\ : InMux
    port map (
            O => \N__32504\,
            I => \N__32493\
        );

    \I__6304\ : LocalMux
    port map (
            O => \N__32499\,
            I => \phase_controller_inst1.stateZ0Z_3\
        );

    \I__6303\ : LocalMux
    port map (
            O => \N__32496\,
            I => \phase_controller_inst1.stateZ0Z_3\
        );

    \I__6302\ : LocalMux
    port map (
            O => \N__32493\,
            I => \phase_controller_inst1.stateZ0Z_3\
        );

    \I__6301\ : InMux
    port map (
            O => \N__32486\,
            I => \N__32483\
        );

    \I__6300\ : LocalMux
    port map (
            O => \N__32483\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_3\
        );

    \I__6299\ : InMux
    port map (
            O => \N__32480\,
            I => \N__32477\
        );

    \I__6298\ : LocalMux
    port map (
            O => \N__32477\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_4\
        );

    \I__6297\ : InMux
    port map (
            O => \N__32474\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\
        );

    \I__6296\ : InMux
    port map (
            O => \N__32471\,
            I => \N__32468\
        );

    \I__6295\ : LocalMux
    port map (
            O => \N__32468\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_5\
        );

    \I__6294\ : InMux
    port map (
            O => \N__32465\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\
        );

    \I__6293\ : InMux
    port map (
            O => \N__32462\,
            I => \N__32459\
        );

    \I__6292\ : LocalMux
    port map (
            O => \N__32459\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_6\
        );

    \I__6291\ : InMux
    port map (
            O => \N__32456\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\
        );

    \I__6290\ : InMux
    port map (
            O => \N__32453\,
            I => \N__32450\
        );

    \I__6289\ : LocalMux
    port map (
            O => \N__32450\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_7\
        );

    \I__6288\ : InMux
    port map (
            O => \N__32447\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\
        );

    \I__6287\ : InMux
    port map (
            O => \N__32444\,
            I => \N__32441\
        );

    \I__6286\ : LocalMux
    port map (
            O => \N__32441\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt8\
        );

    \I__6285\ : CascadeMux
    port map (
            O => \N__32438\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8_cascade_\
        );

    \I__6284\ : InMux
    port map (
            O => \N__32435\,
            I => \N__32432\
        );

    \I__6283\ : LocalMux
    port map (
            O => \N__32432\,
            I => \N__32429\
        );

    \I__6282\ : Odrv4
    port map (
            O => \N__32429\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_10\
        );

    \I__6281\ : InMux
    port map (
            O => \N__32426\,
            I => \N__32423\
        );

    \I__6280\ : LocalMux
    port map (
            O => \N__32423\,
            I => \N__32420\
        );

    \I__6279\ : Span4Mux_v
    port map (
            O => \N__32420\,
            I => \N__32417\
        );

    \I__6278\ : Odrv4
    port map (
            O => \N__32417\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_13\
        );

    \I__6277\ : IoInMux
    port map (
            O => \N__32414\,
            I => \N__32411\
        );

    \I__6276\ : LocalMux
    port map (
            O => \N__32411\,
            I => \N__32408\
        );

    \I__6275\ : Span4Mux_s0_v
    port map (
            O => \N__32408\,
            I => \N__32405\
        );

    \I__6274\ : Sp12to4
    port map (
            O => \N__32405\,
            I => \N__32402\
        );

    \I__6273\ : Span12Mux_h
    port map (
            O => \N__32402\,
            I => \N__32399\
        );

    \I__6272\ : Span12Mux_v
    port map (
            O => \N__32399\,
            I => \N__32396\
        );

    \I__6271\ : Odrv12
    port map (
            O => \N__32396\,
            I => \current_shift_inst.timer_s1.N_187_i\
        );

    \I__6270\ : InMux
    port map (
            O => \N__32393\,
            I => \N__32389\
        );

    \I__6269\ : CascadeMux
    port map (
            O => \N__32392\,
            I => \N__32386\
        );

    \I__6268\ : LocalMux
    port map (
            O => \N__32389\,
            I => \N__32382\
        );

    \I__6267\ : InMux
    port map (
            O => \N__32386\,
            I => \N__32375\
        );

    \I__6266\ : InMux
    port map (
            O => \N__32385\,
            I => \N__32375\
        );

    \I__6265\ : Span4Mux_h
    port map (
            O => \N__32382\,
            I => \N__32372\
        );

    \I__6264\ : InMux
    port map (
            O => \N__32381\,
            I => \N__32367\
        );

    \I__6263\ : InMux
    port map (
            O => \N__32380\,
            I => \N__32367\
        );

    \I__6262\ : LocalMux
    port map (
            O => \N__32375\,
            I => \N__32362\
        );

    \I__6261\ : Span4Mux_h
    port map (
            O => \N__32372\,
            I => \N__32362\
        );

    \I__6260\ : LocalMux
    port map (
            O => \N__32367\,
            I => \current_shift_inst.phase_validZ0\
        );

    \I__6259\ : Odrv4
    port map (
            O => \N__32362\,
            I => \current_shift_inst.phase_validZ0\
        );

    \I__6258\ : CascadeMux
    port map (
            O => \N__32357\,
            I => \N__32353\
        );

    \I__6257\ : CascadeMux
    port map (
            O => \N__32356\,
            I => \N__32347\
        );

    \I__6256\ : InMux
    port map (
            O => \N__32353\,
            I => \N__32342\
        );

    \I__6255\ : InMux
    port map (
            O => \N__32352\,
            I => \N__32342\
        );

    \I__6254\ : InMux
    port map (
            O => \N__32351\,
            I => \N__32335\
        );

    \I__6253\ : InMux
    port map (
            O => \N__32350\,
            I => \N__32335\
        );

    \I__6252\ : InMux
    port map (
            O => \N__32347\,
            I => \N__32335\
        );

    \I__6251\ : LocalMux
    port map (
            O => \N__32342\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__6250\ : LocalMux
    port map (
            O => \N__32335\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__6249\ : InMux
    port map (
            O => \N__32330\,
            I => \N__32324\
        );

    \I__6248\ : InMux
    port map (
            O => \N__32329\,
            I => \N__32321\
        );

    \I__6247\ : InMux
    port map (
            O => \N__32328\,
            I => \N__32316\
        );

    \I__6246\ : InMux
    port map (
            O => \N__32327\,
            I => \N__32316\
        );

    \I__6245\ : LocalMux
    port map (
            O => \N__32324\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__6244\ : LocalMux
    port map (
            O => \N__32321\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__6243\ : LocalMux
    port map (
            O => \N__32316\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__6242\ : CascadeMux
    port map (
            O => \N__32309\,
            I => \N__32301\
        );

    \I__6241\ : InMux
    port map (
            O => \N__32308\,
            I => \N__32293\
        );

    \I__6240\ : InMux
    port map (
            O => \N__32307\,
            I => \N__32293\
        );

    \I__6239\ : InMux
    port map (
            O => \N__32306\,
            I => \N__32293\
        );

    \I__6238\ : InMux
    port map (
            O => \N__32305\,
            I => \N__32288\
        );

    \I__6237\ : InMux
    port map (
            O => \N__32304\,
            I => \N__32288\
        );

    \I__6236\ : InMux
    port map (
            O => \N__32301\,
            I => \N__32283\
        );

    \I__6235\ : InMux
    port map (
            O => \N__32300\,
            I => \N__32283\
        );

    \I__6234\ : LocalMux
    port map (
            O => \N__32293\,
            I => \current_shift_inst.meas_stateZ0Z_0\
        );

    \I__6233\ : LocalMux
    port map (
            O => \N__32288\,
            I => \current_shift_inst.meas_stateZ0Z_0\
        );

    \I__6232\ : LocalMux
    port map (
            O => \N__32283\,
            I => \current_shift_inst.meas_stateZ0Z_0\
        );

    \I__6231\ : CascadeMux
    port map (
            O => \N__32276\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto5Z0Z_3_cascade_\
        );

    \I__6230\ : IoInMux
    port map (
            O => \N__32273\,
            I => \N__32270\
        );

    \I__6229\ : LocalMux
    port map (
            O => \N__32270\,
            I => \N__32267\
        );

    \I__6228\ : Span4Mux_s0_v
    port map (
            O => \N__32267\,
            I => \N__32264\
        );

    \I__6227\ : Span4Mux_v
    port map (
            O => \N__32264\,
            I => \N__32261\
        );

    \I__6226\ : Odrv4
    port map (
            O => \N__32261\,
            I => \delay_measurement_inst.delay_hc_timer.N_321_i\
        );

    \I__6225\ : CascadeMux
    port map (
            O => \N__32258\,
            I => \current_shift_inst.N_199_cascade_\
        );

    \I__6224\ : InMux
    port map (
            O => \N__32255\,
            I => \N__32252\
        );

    \I__6223\ : LocalMux
    port map (
            O => \N__32252\,
            I => \N__32247\
        );

    \I__6222\ : CascadeMux
    port map (
            O => \N__32251\,
            I => \N__32243\
        );

    \I__6221\ : InMux
    port map (
            O => \N__32250\,
            I => \N__32240\
        );

    \I__6220\ : Span4Mux_v
    port map (
            O => \N__32247\,
            I => \N__32237\
        );

    \I__6219\ : InMux
    port map (
            O => \N__32246\,
            I => \N__32234\
        );

    \I__6218\ : InMux
    port map (
            O => \N__32243\,
            I => \N__32231\
        );

    \I__6217\ : LocalMux
    port map (
            O => \N__32240\,
            I => \N__32228\
        );

    \I__6216\ : Odrv4
    port map (
            O => \N__32237\,
            I => \phase_controller_slave.stateZ0Z_1\
        );

    \I__6215\ : LocalMux
    port map (
            O => \N__32234\,
            I => \phase_controller_slave.stateZ0Z_1\
        );

    \I__6214\ : LocalMux
    port map (
            O => \N__32231\,
            I => \phase_controller_slave.stateZ0Z_1\
        );

    \I__6213\ : Odrv4
    port map (
            O => \N__32228\,
            I => \phase_controller_slave.stateZ0Z_1\
        );

    \I__6212\ : InMux
    port map (
            O => \N__32219\,
            I => \N__32214\
        );

    \I__6211\ : InMux
    port map (
            O => \N__32218\,
            I => \N__32211\
        );

    \I__6210\ : InMux
    port map (
            O => \N__32217\,
            I => \N__32208\
        );

    \I__6209\ : LocalMux
    port map (
            O => \N__32214\,
            I => \N__32203\
        );

    \I__6208\ : LocalMux
    port map (
            O => \N__32211\,
            I => \N__32203\
        );

    \I__6207\ : LocalMux
    port map (
            O => \N__32208\,
            I => \N__32200\
        );

    \I__6206\ : Span4Mux_h
    port map (
            O => \N__32203\,
            I => \N__32197\
        );

    \I__6205\ : Span4Mux_h
    port map (
            O => \N__32200\,
            I => \N__32194\
        );

    \I__6204\ : Span4Mux_v
    port map (
            O => \N__32197\,
            I => \N__32191\
        );

    \I__6203\ : Span4Mux_v
    port map (
            O => \N__32194\,
            I => \N__32188\
        );

    \I__6202\ : Sp12to4
    port map (
            O => \N__32191\,
            I => \N__32185\
        );

    \I__6201\ : Span4Mux_v
    port map (
            O => \N__32188\,
            I => \N__32182\
        );

    \I__6200\ : Span12Mux_v
    port map (
            O => \N__32185\,
            I => \N__32179\
        );

    \I__6199\ : Span4Mux_v
    port map (
            O => \N__32182\,
            I => \N__32176\
        );

    \I__6198\ : Odrv12
    port map (
            O => \N__32179\,
            I => \il_min_comp2_D2\
        );

    \I__6197\ : Odrv4
    port map (
            O => \N__32176\,
            I => \il_min_comp2_D2\
        );

    \I__6196\ : CascadeMux
    port map (
            O => \N__32171\,
            I => \N__32168\
        );

    \I__6195\ : InMux
    port map (
            O => \N__32168\,
            I => \N__32163\
        );

    \I__6194\ : InMux
    port map (
            O => \N__32167\,
            I => \N__32158\
        );

    \I__6193\ : InMux
    port map (
            O => \N__32166\,
            I => \N__32158\
        );

    \I__6192\ : LocalMux
    port map (
            O => \N__32163\,
            I => \il_max_comp2_D2\
        );

    \I__6191\ : LocalMux
    port map (
            O => \N__32158\,
            I => \il_max_comp2_D2\
        );

    \I__6190\ : InMux
    port map (
            O => \N__32153\,
            I => \N__32145\
        );

    \I__6189\ : InMux
    port map (
            O => \N__32152\,
            I => \N__32145\
        );

    \I__6188\ : InMux
    port map (
            O => \N__32151\,
            I => \N__32140\
        );

    \I__6187\ : InMux
    port map (
            O => \N__32150\,
            I => \N__32140\
        );

    \I__6186\ : LocalMux
    port map (
            O => \N__32145\,
            I => \phase_controller_slave.stateZ0Z_3\
        );

    \I__6185\ : LocalMux
    port map (
            O => \N__32140\,
            I => \phase_controller_slave.stateZ0Z_3\
        );

    \I__6184\ : CEMux
    port map (
            O => \N__32135\,
            I => \N__32130\
        );

    \I__6183\ : CEMux
    port map (
            O => \N__32134\,
            I => \N__32127\
        );

    \I__6182\ : CEMux
    port map (
            O => \N__32133\,
            I => \N__32123\
        );

    \I__6181\ : LocalMux
    port map (
            O => \N__32130\,
            I => \N__32120\
        );

    \I__6180\ : LocalMux
    port map (
            O => \N__32127\,
            I => \N__32117\
        );

    \I__6179\ : CEMux
    port map (
            O => \N__32126\,
            I => \N__32114\
        );

    \I__6178\ : LocalMux
    port map (
            O => \N__32123\,
            I => \N__32111\
        );

    \I__6177\ : Span4Mux_v
    port map (
            O => \N__32120\,
            I => \N__32106\
        );

    \I__6176\ : Span4Mux_v
    port map (
            O => \N__32117\,
            I => \N__32106\
        );

    \I__6175\ : LocalMux
    port map (
            O => \N__32114\,
            I => \N__32103\
        );

    \I__6174\ : Span4Mux_v
    port map (
            O => \N__32111\,
            I => \N__32098\
        );

    \I__6173\ : Span4Mux_h
    port map (
            O => \N__32106\,
            I => \N__32098\
        );

    \I__6172\ : Span4Mux_h
    port map (
            O => \N__32103\,
            I => \N__32095\
        );

    \I__6171\ : Odrv4
    port map (
            O => \N__32098\,
            I => \current_shift_inst.timer_phase.N_192_i\
        );

    \I__6170\ : Odrv4
    port map (
            O => \N__32095\,
            I => \current_shift_inst.timer_phase.N_192_i\
        );

    \I__6169\ : InMux
    port map (
            O => \N__32090\,
            I => \N__32056\
        );

    \I__6168\ : InMux
    port map (
            O => \N__32089\,
            I => \N__32056\
        );

    \I__6167\ : InMux
    port map (
            O => \N__32088\,
            I => \N__32047\
        );

    \I__6166\ : InMux
    port map (
            O => \N__32087\,
            I => \N__32047\
        );

    \I__6165\ : InMux
    port map (
            O => \N__32086\,
            I => \N__32047\
        );

    \I__6164\ : InMux
    port map (
            O => \N__32085\,
            I => \N__32047\
        );

    \I__6163\ : InMux
    port map (
            O => \N__32084\,
            I => \N__32038\
        );

    \I__6162\ : InMux
    port map (
            O => \N__32083\,
            I => \N__32038\
        );

    \I__6161\ : InMux
    port map (
            O => \N__32082\,
            I => \N__32038\
        );

    \I__6160\ : InMux
    port map (
            O => \N__32081\,
            I => \N__32038\
        );

    \I__6159\ : InMux
    port map (
            O => \N__32080\,
            I => \N__32029\
        );

    \I__6158\ : InMux
    port map (
            O => \N__32079\,
            I => \N__32029\
        );

    \I__6157\ : InMux
    port map (
            O => \N__32078\,
            I => \N__32029\
        );

    \I__6156\ : InMux
    port map (
            O => \N__32077\,
            I => \N__32029\
        );

    \I__6155\ : InMux
    port map (
            O => \N__32076\,
            I => \N__32020\
        );

    \I__6154\ : InMux
    port map (
            O => \N__32075\,
            I => \N__32020\
        );

    \I__6153\ : InMux
    port map (
            O => \N__32074\,
            I => \N__32020\
        );

    \I__6152\ : InMux
    port map (
            O => \N__32073\,
            I => \N__32020\
        );

    \I__6151\ : InMux
    port map (
            O => \N__32072\,
            I => \N__32011\
        );

    \I__6150\ : InMux
    port map (
            O => \N__32071\,
            I => \N__32011\
        );

    \I__6149\ : InMux
    port map (
            O => \N__32070\,
            I => \N__32011\
        );

    \I__6148\ : InMux
    port map (
            O => \N__32069\,
            I => \N__32011\
        );

    \I__6147\ : InMux
    port map (
            O => \N__32068\,
            I => \N__32002\
        );

    \I__6146\ : InMux
    port map (
            O => \N__32067\,
            I => \N__32002\
        );

    \I__6145\ : InMux
    port map (
            O => \N__32066\,
            I => \N__32002\
        );

    \I__6144\ : InMux
    port map (
            O => \N__32065\,
            I => \N__32002\
        );

    \I__6143\ : InMux
    port map (
            O => \N__32064\,
            I => \N__31993\
        );

    \I__6142\ : InMux
    port map (
            O => \N__32063\,
            I => \N__31993\
        );

    \I__6141\ : InMux
    port map (
            O => \N__32062\,
            I => \N__31993\
        );

    \I__6140\ : InMux
    port map (
            O => \N__32061\,
            I => \N__31993\
        );

    \I__6139\ : LocalMux
    port map (
            O => \N__32056\,
            I => \N__31988\
        );

    \I__6138\ : LocalMux
    port map (
            O => \N__32047\,
            I => \N__31988\
        );

    \I__6137\ : LocalMux
    port map (
            O => \N__32038\,
            I => \N__31983\
        );

    \I__6136\ : LocalMux
    port map (
            O => \N__32029\,
            I => \N__31983\
        );

    \I__6135\ : LocalMux
    port map (
            O => \N__32020\,
            I => \N__31978\
        );

    \I__6134\ : LocalMux
    port map (
            O => \N__32011\,
            I => \N__31978\
        );

    \I__6133\ : LocalMux
    port map (
            O => \N__32002\,
            I => \N__31973\
        );

    \I__6132\ : LocalMux
    port map (
            O => \N__31993\,
            I => \N__31973\
        );

    \I__6131\ : Span4Mux_h
    port map (
            O => \N__31988\,
            I => \N__31970\
        );

    \I__6130\ : Span4Mux_h
    port map (
            O => \N__31983\,
            I => \N__31967\
        );

    \I__6129\ : Span4Mux_h
    port map (
            O => \N__31978\,
            I => \N__31964\
        );

    \I__6128\ : Odrv4
    port map (
            O => \N__31973\,
            I => \current_shift_inst.timer_phase.running_i\
        );

    \I__6127\ : Odrv4
    port map (
            O => \N__31970\,
            I => \current_shift_inst.timer_phase.running_i\
        );

    \I__6126\ : Odrv4
    port map (
            O => \N__31967\,
            I => \current_shift_inst.timer_phase.running_i\
        );

    \I__6125\ : Odrv4
    port map (
            O => \N__31964\,
            I => \current_shift_inst.timer_phase.running_i\
        );

    \I__6124\ : InMux
    port map (
            O => \N__31955\,
            I => \N__31952\
        );

    \I__6123\ : LocalMux
    port map (
            O => \N__31952\,
            I => \N__31949\
        );

    \I__6122\ : Glb2LocalMux
    port map (
            O => \N__31949\,
            I => \N__31946\
        );

    \I__6121\ : GlobalMux
    port map (
            O => \N__31946\,
            I => clk_12mhz
        );

    \I__6120\ : IoInMux
    port map (
            O => \N__31943\,
            I => \N__31940\
        );

    \I__6119\ : LocalMux
    port map (
            O => \N__31940\,
            I => \N__31937\
        );

    \I__6118\ : Span12Mux_s0_v
    port map (
            O => \N__31937\,
            I => \N__31934\
        );

    \I__6117\ : Odrv12
    port map (
            O => \N__31934\,
            I => \GB_BUFFER_clk_12mhz_THRU_CO\
        );

    \I__6116\ : CascadeMux
    port map (
            O => \N__31931\,
            I => \N__31928\
        );

    \I__6115\ : InMux
    port map (
            O => \N__31928\,
            I => \N__31925\
        );

    \I__6114\ : LocalMux
    port map (
            O => \N__31925\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1Z0Z_6\
        );

    \I__6113\ : CascadeMux
    port map (
            O => \N__31922\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1Z0Z_6_cascade_\
        );

    \I__6112\ : CascadeMux
    port map (
            O => \N__31919\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6_cascade_\
        );

    \I__6111\ : CascadeMux
    port map (
            O => \N__31916\,
            I => \phase_controller_slave.start_timer_hc_0_sqmuxa_cascade_\
        );

    \I__6110\ : IoInMux
    port map (
            O => \N__31913\,
            I => \N__31910\
        );

    \I__6109\ : LocalMux
    port map (
            O => \N__31910\,
            I => \N__31907\
        );

    \I__6108\ : IoSpan4Mux
    port map (
            O => \N__31907\,
            I => \N__31904\
        );

    \I__6107\ : Span4Mux_s3_v
    port map (
            O => \N__31904\,
            I => \N__31900\
        );

    \I__6106\ : InMux
    port map (
            O => \N__31903\,
            I => \N__31897\
        );

    \I__6105\ : Span4Mux_v
    port map (
            O => \N__31900\,
            I => \N__31894\
        );

    \I__6104\ : LocalMux
    port map (
            O => \N__31897\,
            I => \N__31891\
        );

    \I__6103\ : Odrv4
    port map (
            O => \N__31894\,
            I => s3_phy_c
        );

    \I__6102\ : Odrv12
    port map (
            O => \N__31891\,
            I => s3_phy_c
        );

    \I__6101\ : CascadeMux
    port map (
            O => \N__31886\,
            I => \N__31883\
        );

    \I__6100\ : InMux
    port map (
            O => \N__31883\,
            I => \N__31880\
        );

    \I__6099\ : LocalMux
    port map (
            O => \N__31880\,
            I => \N__31877\
        );

    \I__6098\ : Span4Mux_h
    port map (
            O => \N__31877\,
            I => \N__31874\
        );

    \I__6097\ : Odrv4
    port map (
            O => \N__31874\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI1C4K_24\
        );

    \I__6096\ : CascadeMux
    port map (
            O => \N__31871\,
            I => \N__31868\
        );

    \I__6095\ : InMux
    port map (
            O => \N__31868\,
            I => \N__31863\
        );

    \I__6094\ : InMux
    port map (
            O => \N__31867\,
            I => \N__31860\
        );

    \I__6093\ : InMux
    port map (
            O => \N__31866\,
            I => \N__31856\
        );

    \I__6092\ : LocalMux
    port map (
            O => \N__31863\,
            I => \N__31853\
        );

    \I__6091\ : LocalMux
    port map (
            O => \N__31860\,
            I => \N__31850\
        );

    \I__6090\ : InMux
    port map (
            O => \N__31859\,
            I => \N__31847\
        );

    \I__6089\ : LocalMux
    port map (
            O => \N__31856\,
            I => \N__31842\
        );

    \I__6088\ : Span12Mux_h
    port map (
            O => \N__31853\,
            I => \N__31842\
        );

    \I__6087\ : Span4Mux_h
    port map (
            O => \N__31850\,
            I => \N__31837\
        );

    \I__6086\ : LocalMux
    port map (
            O => \N__31847\,
            I => \N__31837\
        );

    \I__6085\ : Odrv12
    port map (
            O => \N__31842\,
            I => \current_shift_inst.elapsed_time_ns_phase_26\
        );

    \I__6084\ : Odrv4
    port map (
            O => \N__31837\,
            I => \current_shift_inst.elapsed_time_ns_phase_26\
        );

    \I__6083\ : CascadeMux
    port map (
            O => \N__31832\,
            I => \N__31829\
        );

    \I__6082\ : InMux
    port map (
            O => \N__31829\,
            I => \N__31826\
        );

    \I__6081\ : LocalMux
    port map (
            O => \N__31826\,
            I => \N__31820\
        );

    \I__6080\ : InMux
    port map (
            O => \N__31825\,
            I => \N__31817\
        );

    \I__6079\ : CascadeMux
    port map (
            O => \N__31824\,
            I => \N__31814\
        );

    \I__6078\ : InMux
    port map (
            O => \N__31823\,
            I => \N__31811\
        );

    \I__6077\ : Span4Mux_h
    port map (
            O => \N__31820\,
            I => \N__31806\
        );

    \I__6076\ : LocalMux
    port map (
            O => \N__31817\,
            I => \N__31806\
        );

    \I__6075\ : InMux
    port map (
            O => \N__31814\,
            I => \N__31803\
        );

    \I__6074\ : LocalMux
    port map (
            O => \N__31811\,
            I => \current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0\
        );

    \I__6073\ : Odrv4
    port map (
            O => \N__31806\,
            I => \current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__31803\,
            I => \current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0\
        );

    \I__6071\ : InMux
    port map (
            O => \N__31796\,
            I => \N__31793\
        );

    \I__6070\ : LocalMux
    port map (
            O => \N__31793\,
            I => \N__31790\
        );

    \I__6069\ : Span4Mux_h
    port map (
            O => \N__31790\,
            I => \N__31787\
        );

    \I__6068\ : Odrv4
    port map (
            O => \N__31787\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIB4C81_25\
        );

    \I__6067\ : InMux
    port map (
            O => \N__31784\,
            I => \N__31779\
        );

    \I__6066\ : InMux
    port map (
            O => \N__31783\,
            I => \N__31774\
        );

    \I__6065\ : InMux
    port map (
            O => \N__31782\,
            I => \N__31774\
        );

    \I__6064\ : LocalMux
    port map (
            O => \N__31779\,
            I => \N__31769\
        );

    \I__6063\ : LocalMux
    port map (
            O => \N__31774\,
            I => \N__31769\
        );

    \I__6062\ : Span4Mux_h
    port map (
            O => \N__31769\,
            I => \N__31765\
        );

    \I__6061\ : InMux
    port map (
            O => \N__31768\,
            I => \N__31762\
        );

    \I__6060\ : Span4Mux_v
    port map (
            O => \N__31765\,
            I => \N__31759\
        );

    \I__6059\ : LocalMux
    port map (
            O => \N__31762\,
            I => \N__31756\
        );

    \I__6058\ : Odrv4
    port map (
            O => \N__31759\,
            I => \current_shift_inst.elapsed_time_ns_phase_25\
        );

    \I__6057\ : Odrv4
    port map (
            O => \N__31756\,
            I => \current_shift_inst.elapsed_time_ns_phase_25\
        );

    \I__6056\ : InMux
    port map (
            O => \N__31751\,
            I => \N__31743\
        );

    \I__6055\ : InMux
    port map (
            O => \N__31750\,
            I => \N__31743\
        );

    \I__6054\ : InMux
    port map (
            O => \N__31749\,
            I => \N__31740\
        );

    \I__6053\ : InMux
    port map (
            O => \N__31748\,
            I => \N__31737\
        );

    \I__6052\ : LocalMux
    port map (
            O => \N__31743\,
            I => \current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0\
        );

    \I__6051\ : LocalMux
    port map (
            O => \N__31740\,
            I => \current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0\
        );

    \I__6050\ : LocalMux
    port map (
            O => \N__31737\,
            I => \current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0\
        );

    \I__6049\ : CascadeMux
    port map (
            O => \N__31730\,
            I => \N__31727\
        );

    \I__6048\ : InMux
    port map (
            O => \N__31727\,
            I => \N__31724\
        );

    \I__6047\ : LocalMux
    port map (
            O => \N__31724\,
            I => \N__31721\
        );

    \I__6046\ : Span4Mux_v
    port map (
            O => \N__31721\,
            I => \N__31718\
        );

    \I__6045\ : Span4Mux_h
    port map (
            O => \N__31718\,
            I => \N__31715\
        );

    \I__6044\ : Odrv4
    port map (
            O => \N__31715\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI4G5K_25\
        );

    \I__6043\ : InMux
    port map (
            O => \N__31712\,
            I => \N__31709\
        );

    \I__6042\ : LocalMux
    port map (
            O => \N__31709\,
            I => \N__31706\
        );

    \I__6041\ : Span4Mux_v
    port map (
            O => \N__31706\,
            I => \N__31701\
        );

    \I__6040\ : InMux
    port map (
            O => \N__31705\,
            I => \N__31698\
        );

    \I__6039\ : InMux
    port map (
            O => \N__31704\,
            I => \N__31695\
        );

    \I__6038\ : Span4Mux_h
    port map (
            O => \N__31701\,
            I => \N__31692\
        );

    \I__6037\ : LocalMux
    port map (
            O => \N__31698\,
            I => \N__31689\
        );

    \I__6036\ : LocalMux
    port map (
            O => \N__31695\,
            I => \N__31686\
        );

    \I__6035\ : Odrv4
    port map (
            O => \N__31692\,
            I => \current_shift_inst.elapsed_time_ns_phase_29\
        );

    \I__6034\ : Odrv12
    port map (
            O => \N__31689\,
            I => \current_shift_inst.elapsed_time_ns_phase_29\
        );

    \I__6033\ : Odrv4
    port map (
            O => \N__31686\,
            I => \current_shift_inst.elapsed_time_ns_phase_29\
        );

    \I__6032\ : InMux
    port map (
            O => \N__31679\,
            I => \N__31676\
        );

    \I__6031\ : LocalMux
    port map (
            O => \N__31676\,
            I => \N__31672\
        );

    \I__6030\ : InMux
    port map (
            O => \N__31675\,
            I => \N__31668\
        );

    \I__6029\ : Span4Mux_h
    port map (
            O => \N__31672\,
            I => \N__31665\
        );

    \I__6028\ : InMux
    port map (
            O => \N__31671\,
            I => \N__31662\
        );

    \I__6027\ : LocalMux
    port map (
            O => \N__31668\,
            I => \current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0\
        );

    \I__6026\ : Odrv4
    port map (
            O => \N__31665\,
            I => \current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0\
        );

    \I__6025\ : LocalMux
    port map (
            O => \N__31662\,
            I => \current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0\
        );

    \I__6024\ : InMux
    port map (
            O => \N__31655\,
            I => \N__31651\
        );

    \I__6023\ : CascadeMux
    port map (
            O => \N__31654\,
            I => \N__31648\
        );

    \I__6022\ : LocalMux
    port map (
            O => \N__31651\,
            I => \N__31645\
        );

    \I__6021\ : InMux
    port map (
            O => \N__31648\,
            I => \N__31642\
        );

    \I__6020\ : Span4Mux_v
    port map (
            O => \N__31645\,
            I => \N__31639\
        );

    \I__6019\ : LocalMux
    port map (
            O => \N__31642\,
            I => \N__31636\
        );

    \I__6018\ : Span4Mux_h
    port map (
            O => \N__31639\,
            I => \N__31631\
        );

    \I__6017\ : Span4Mux_v
    port map (
            O => \N__31636\,
            I => \N__31631\
        );

    \I__6016\ : Odrv4
    port map (
            O => \N__31631\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI7OAK_29\
        );

    \I__6015\ : InMux
    port map (
            O => \N__31628\,
            I => \N__31623\
        );

    \I__6014\ : InMux
    port map (
            O => \N__31627\,
            I => \N__31617\
        );

    \I__6013\ : InMux
    port map (
            O => \N__31626\,
            I => \N__31617\
        );

    \I__6012\ : LocalMux
    port map (
            O => \N__31623\,
            I => \N__31614\
        );

    \I__6011\ : InMux
    port map (
            O => \N__31622\,
            I => \N__31611\
        );

    \I__6010\ : LocalMux
    port map (
            O => \N__31617\,
            I => \N__31608\
        );

    \I__6009\ : Span4Mux_v
    port map (
            O => \N__31614\,
            I => \N__31603\
        );

    \I__6008\ : LocalMux
    port map (
            O => \N__31611\,
            I => \N__31603\
        );

    \I__6007\ : Span12Mux_v
    port map (
            O => \N__31608\,
            I => \N__31600\
        );

    \I__6006\ : Span4Mux_v
    port map (
            O => \N__31603\,
            I => \N__31597\
        );

    \I__6005\ : Odrv12
    port map (
            O => \N__31600\,
            I => \current_shift_inst.elapsed_time_ns_phase_24\
        );

    \I__6004\ : Odrv4
    port map (
            O => \N__31597\,
            I => \current_shift_inst.elapsed_time_ns_phase_24\
        );

    \I__6003\ : InMux
    port map (
            O => \N__31592\,
            I => \N__31589\
        );

    \I__6002\ : LocalMux
    port map (
            O => \N__31589\,
            I => \N__31584\
        );

    \I__6001\ : InMux
    port map (
            O => \N__31588\,
            I => \N__31581\
        );

    \I__6000\ : InMux
    port map (
            O => \N__31587\,
            I => \N__31578\
        );

    \I__5999\ : Span4Mux_h
    port map (
            O => \N__31584\,
            I => \N__31573\
        );

    \I__5998\ : LocalMux
    port map (
            O => \N__31581\,
            I => \N__31573\
        );

    \I__5997\ : LocalMux
    port map (
            O => \N__31578\,
            I => \N__31569\
        );

    \I__5996\ : Span4Mux_v
    port map (
            O => \N__31573\,
            I => \N__31566\
        );

    \I__5995\ : InMux
    port map (
            O => \N__31572\,
            I => \N__31563\
        );

    \I__5994\ : Odrv4
    port map (
            O => \N__31569\,
            I => \current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0\
        );

    \I__5993\ : Odrv4
    port map (
            O => \N__31566\,
            I => \current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0\
        );

    \I__5992\ : LocalMux
    port map (
            O => \N__31563\,
            I => \current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0\
        );

    \I__5991\ : CascadeMux
    port map (
            O => \N__31556\,
            I => \N__31553\
        );

    \I__5990\ : InMux
    port map (
            O => \N__31553\,
            I => \N__31550\
        );

    \I__5989\ : LocalMux
    port map (
            O => \N__31550\,
            I => \N__31545\
        );

    \I__5988\ : InMux
    port map (
            O => \N__31549\,
            I => \N__31541\
        );

    \I__5987\ : InMux
    port map (
            O => \N__31548\,
            I => \N__31538\
        );

    \I__5986\ : Span4Mux_v
    port map (
            O => \N__31545\,
            I => \N__31535\
        );

    \I__5985\ : InMux
    port map (
            O => \N__31544\,
            I => \N__31532\
        );

    \I__5984\ : LocalMux
    port map (
            O => \N__31541\,
            I => \N__31529\
        );

    \I__5983\ : LocalMux
    port map (
            O => \N__31538\,
            I => \N__31526\
        );

    \I__5982\ : Span4Mux_h
    port map (
            O => \N__31535\,
            I => \N__31521\
        );

    \I__5981\ : LocalMux
    port map (
            O => \N__31532\,
            I => \N__31521\
        );

    \I__5980\ : Span4Mux_v
    port map (
            O => \N__31529\,
            I => \N__31518\
        );

    \I__5979\ : Span4Mux_v
    port map (
            O => \N__31526\,
            I => \N__31515\
        );

    \I__5978\ : Odrv4
    port map (
            O => \N__31521\,
            I => \current_shift_inst.elapsed_time_ns_phase_23\
        );

    \I__5977\ : Odrv4
    port map (
            O => \N__31518\,
            I => \current_shift_inst.elapsed_time_ns_phase_23\
        );

    \I__5976\ : Odrv4
    port map (
            O => \N__31515\,
            I => \current_shift_inst.elapsed_time_ns_phase_23\
        );

    \I__5975\ : CascadeMux
    port map (
            O => \N__31508\,
            I => \N__31504\
        );

    \I__5974\ : CascadeMux
    port map (
            O => \N__31507\,
            I => \N__31499\
        );

    \I__5973\ : InMux
    port map (
            O => \N__31504\,
            I => \N__31496\
        );

    \I__5972\ : InMux
    port map (
            O => \N__31503\,
            I => \N__31491\
        );

    \I__5971\ : InMux
    port map (
            O => \N__31502\,
            I => \N__31491\
        );

    \I__5970\ : InMux
    port map (
            O => \N__31499\,
            I => \N__31488\
        );

    \I__5969\ : LocalMux
    port map (
            O => \N__31496\,
            I => \current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0\
        );

    \I__5968\ : LocalMux
    port map (
            O => \N__31491\,
            I => \current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0\
        );

    \I__5967\ : LocalMux
    port map (
            O => \N__31488\,
            I => \current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0\
        );

    \I__5966\ : InMux
    port map (
            O => \N__31481\,
            I => \N__31478\
        );

    \I__5965\ : LocalMux
    port map (
            O => \N__31478\,
            I => \N__31475\
        );

    \I__5964\ : Span4Mux_h
    port map (
            O => \N__31475\,
            I => \N__31472\
        );

    \I__5963\ : Odrv4
    port map (
            O => \N__31472\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIVJ781_23\
        );

    \I__5962\ : CascadeMux
    port map (
            O => \N__31469\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3_cascade_\
        );

    \I__5961\ : InMux
    port map (
            O => \N__31466\,
            I => \N__31463\
        );

    \I__5960\ : LocalMux
    port map (
            O => \N__31463\,
            I => \current_shift_inst.un4_control_input_axb_27\
        );

    \I__5959\ : InMux
    port map (
            O => \N__31460\,
            I => \N__31457\
        );

    \I__5958\ : LocalMux
    port map (
            O => \N__31457\,
            I => \current_shift_inst.un4_control_input_axb_30\
        );

    \I__5957\ : InMux
    port map (
            O => \N__31454\,
            I => \N__31451\
        );

    \I__5956\ : LocalMux
    port map (
            O => \N__31451\,
            I => \current_shift_inst.un4_control_input_axb_21\
        );

    \I__5955\ : InMux
    port map (
            O => \N__31448\,
            I => \N__31445\
        );

    \I__5954\ : LocalMux
    port map (
            O => \N__31445\,
            I => \current_shift_inst.un4_control_input_axb_25\
        );

    \I__5953\ : InMux
    port map (
            O => \N__31442\,
            I => \N__31439\
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__31439\,
            I => \current_shift_inst.un4_control_input_axb_20\
        );

    \I__5951\ : InMux
    port map (
            O => \N__31436\,
            I => \N__31432\
        );

    \I__5950\ : InMux
    port map (
            O => \N__31435\,
            I => \N__31429\
        );

    \I__5949\ : LocalMux
    port map (
            O => \N__31432\,
            I => \N__31426\
        );

    \I__5948\ : LocalMux
    port map (
            O => \N__31429\,
            I => \N__31423\
        );

    \I__5947\ : Odrv4
    port map (
            O => \N__31426\,
            I => \current_shift_inst.z_31\
        );

    \I__5946\ : Odrv4
    port map (
            O => \N__31423\,
            I => \current_shift_inst.z_31\
        );

    \I__5945\ : InMux
    port map (
            O => \N__31418\,
            I => \N__31414\
        );

    \I__5944\ : CascadeMux
    port map (
            O => \N__31417\,
            I => \N__31411\
        );

    \I__5943\ : LocalMux
    port map (
            O => \N__31414\,
            I => \N__31408\
        );

    \I__5942\ : InMux
    port map (
            O => \N__31411\,
            I => \N__31405\
        );

    \I__5941\ : Sp12to4
    port map (
            O => \N__31408\,
            I => \N__31400\
        );

    \I__5940\ : LocalMux
    port map (
            O => \N__31405\,
            I => \N__31400\
        );

    \I__5939\ : Odrv12
    port map (
            O => \N__31400\,
            I => \current_shift_inst.z_i_31\
        );

    \I__5938\ : InMux
    port map (
            O => \N__31397\,
            I => \N__31394\
        );

    \I__5937\ : LocalMux
    port map (
            O => \N__31394\,
            I => \current_shift_inst.un4_control_input_axb_28\
        );

    \I__5936\ : InMux
    port map (
            O => \N__31391\,
            I => \N__31388\
        );

    \I__5935\ : LocalMux
    port map (
            O => \N__31388\,
            I => \current_shift_inst.un4_control_input_axb_11\
        );

    \I__5934\ : CascadeMux
    port map (
            O => \N__31385\,
            I => \N__31382\
        );

    \I__5933\ : InMux
    port map (
            O => \N__31382\,
            I => \N__31379\
        );

    \I__5932\ : LocalMux
    port map (
            O => \N__31379\,
            I => \current_shift_inst.un4_control_input_axb_19\
        );

    \I__5931\ : InMux
    port map (
            O => \N__31376\,
            I => \N__31373\
        );

    \I__5930\ : LocalMux
    port map (
            O => \N__31373\,
            I => \current_shift_inst.un4_control_input_axb_10\
        );

    \I__5929\ : InMux
    port map (
            O => \N__31370\,
            I => \N__31367\
        );

    \I__5928\ : LocalMux
    port map (
            O => \N__31367\,
            I => \current_shift_inst.un4_control_input_axb_12\
        );

    \I__5927\ : InMux
    port map (
            O => \N__31364\,
            I => \N__31361\
        );

    \I__5926\ : LocalMux
    port map (
            O => \N__31361\,
            I => \current_shift_inst.un4_control_input_axb_14\
        );

    \I__5925\ : InMux
    port map (
            O => \N__31358\,
            I => \N__31355\
        );

    \I__5924\ : LocalMux
    port map (
            O => \N__31355\,
            I => \current_shift_inst.un4_control_input_axb_18\
        );

    \I__5923\ : InMux
    port map (
            O => \N__31352\,
            I => \N__31349\
        );

    \I__5922\ : LocalMux
    port map (
            O => \N__31349\,
            I => \current_shift_inst.un4_control_input_axb_29\
        );

    \I__5921\ : InMux
    port map (
            O => \N__31346\,
            I => \N__31343\
        );

    \I__5920\ : LocalMux
    port map (
            O => \N__31343\,
            I => \current_shift_inst.un4_control_input_axb_22\
        );

    \I__5919\ : InMux
    port map (
            O => \N__31340\,
            I => \N__31337\
        );

    \I__5918\ : LocalMux
    port map (
            O => \N__31337\,
            I => \current_shift_inst.un4_control_input_axb_26\
        );

    \I__5917\ : InMux
    port map (
            O => \N__31334\,
            I => \N__31331\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__31331\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_1\
        );

    \I__5915\ : InMux
    port map (
            O => \N__31328\,
            I => \N__31325\
        );

    \I__5914\ : LocalMux
    port map (
            O => \N__31325\,
            I => \current_shift_inst.un4_control_input_axb_1\
        );

    \I__5913\ : InMux
    port map (
            O => \N__31322\,
            I => \N__31319\
        );

    \I__5912\ : LocalMux
    port map (
            O => \N__31319\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_2\
        );

    \I__5911\ : InMux
    port map (
            O => \N__31316\,
            I => \N__31313\
        );

    \I__5910\ : LocalMux
    port map (
            O => \N__31313\,
            I => \current_shift_inst.un4_control_input_axb_2\
        );

    \I__5909\ : InMux
    port map (
            O => \N__31310\,
            I => \N__31307\
        );

    \I__5908\ : LocalMux
    port map (
            O => \N__31307\,
            I => \current_shift_inst.un4_control_input_axb_24\
        );

    \I__5907\ : InMux
    port map (
            O => \N__31304\,
            I => \N__31301\
        );

    \I__5906\ : LocalMux
    port map (
            O => \N__31301\,
            I => \current_shift_inst.un4_control_input_axb_15\
        );

    \I__5905\ : InMux
    port map (
            O => \N__31298\,
            I => \N__31295\
        );

    \I__5904\ : LocalMux
    port map (
            O => \N__31295\,
            I => \N__31292\
        );

    \I__5903\ : Odrv4
    port map (
            O => \N__31292\,
            I => \current_shift_inst.un4_control_input_axb_5\
        );

    \I__5902\ : CascadeMux
    port map (
            O => \N__31289\,
            I => \N__31286\
        );

    \I__5901\ : InMux
    port map (
            O => \N__31286\,
            I => \N__31283\
        );

    \I__5900\ : LocalMux
    port map (
            O => \N__31283\,
            I => \N__31280\
        );

    \I__5899\ : Odrv4
    port map (
            O => \N__31280\,
            I => \current_shift_inst.un4_control_input_axb_6\
        );

    \I__5898\ : InMux
    port map (
            O => \N__31277\,
            I => \N__31274\
        );

    \I__5897\ : LocalMux
    port map (
            O => \N__31274\,
            I => \N__31271\
        );

    \I__5896\ : Odrv4
    port map (
            O => \N__31271\,
            I => \current_shift_inst.un4_control_input_axb_7\
        );

    \I__5895\ : CascadeMux
    port map (
            O => \N__31268\,
            I => \N__31265\
        );

    \I__5894\ : InMux
    port map (
            O => \N__31265\,
            I => \N__31262\
        );

    \I__5893\ : LocalMux
    port map (
            O => \N__31262\,
            I => \N__31259\
        );

    \I__5892\ : Odrv12
    port map (
            O => \N__31259\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\
        );

    \I__5891\ : CascadeMux
    port map (
            O => \N__31256\,
            I => \N__31253\
        );

    \I__5890\ : InMux
    port map (
            O => \N__31253\,
            I => \N__31250\
        );

    \I__5889\ : LocalMux
    port map (
            O => \N__31250\,
            I => \N__31247\
        );

    \I__5888\ : Odrv12
    port map (
            O => \N__31247\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\
        );

    \I__5887\ : CascadeMux
    port map (
            O => \N__31244\,
            I => \N__31241\
        );

    \I__5886\ : InMux
    port map (
            O => \N__31241\,
            I => \N__31238\
        );

    \I__5885\ : LocalMux
    port map (
            O => \N__31238\,
            I => \N__31235\
        );

    \I__5884\ : Span4Mux_h
    port map (
            O => \N__31235\,
            I => \N__31232\
        );

    \I__5883\ : Odrv4
    port map (
            O => \N__31232\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\
        );

    \I__5882\ : CEMux
    port map (
            O => \N__31229\,
            I => \N__31221\
        );

    \I__5881\ : CEMux
    port map (
            O => \N__31228\,
            I => \N__31218\
        );

    \I__5880\ : CEMux
    port map (
            O => \N__31227\,
            I => \N__31215\
        );

    \I__5879\ : CEMux
    port map (
            O => \N__31226\,
            I => \N__31212\
        );

    \I__5878\ : CEMux
    port map (
            O => \N__31225\,
            I => \N__31209\
        );

    \I__5877\ : CEMux
    port map (
            O => \N__31224\,
            I => \N__31206\
        );

    \I__5876\ : LocalMux
    port map (
            O => \N__31221\,
            I => \N__31203\
        );

    \I__5875\ : LocalMux
    port map (
            O => \N__31218\,
            I => \N__31200\
        );

    \I__5874\ : LocalMux
    port map (
            O => \N__31215\,
            I => \N__31197\
        );

    \I__5873\ : LocalMux
    port map (
            O => \N__31212\,
            I => \N__31194\
        );

    \I__5872\ : LocalMux
    port map (
            O => \N__31209\,
            I => \N__31191\
        );

    \I__5871\ : LocalMux
    port map (
            O => \N__31206\,
            I => \N__31188\
        );

    \I__5870\ : Span4Mux_h
    port map (
            O => \N__31203\,
            I => \N__31185\
        );

    \I__5869\ : Span4Mux_h
    port map (
            O => \N__31200\,
            I => \N__31180\
        );

    \I__5868\ : Span4Mux_v
    port map (
            O => \N__31197\,
            I => \N__31180\
        );

    \I__5867\ : Span4Mux_h
    port map (
            O => \N__31194\,
            I => \N__31177\
        );

    \I__5866\ : Span4Mux_h
    port map (
            O => \N__31191\,
            I => \N__31174\
        );

    \I__5865\ : Odrv12
    port map (
            O => \N__31188\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__5864\ : Odrv4
    port map (
            O => \N__31185\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__5863\ : Odrv4
    port map (
            O => \N__31180\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__5862\ : Odrv4
    port map (
            O => \N__31177\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__5861\ : Odrv4
    port map (
            O => \N__31174\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__5860\ : CascadeMux
    port map (
            O => \N__31163\,
            I => \N__31160\
        );

    \I__5859\ : InMux
    port map (
            O => \N__31160\,
            I => \N__31157\
        );

    \I__5858\ : LocalMux
    port map (
            O => \N__31157\,
            I => \current_shift_inst.un4_control_input_axb_3\
        );

    \I__5857\ : InMux
    port map (
            O => \N__31154\,
            I => \N__31151\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__31151\,
            I => \current_shift_inst.un4_control_input_axb_4\
        );

    \I__5855\ : InMux
    port map (
            O => \N__31148\,
            I => \N__31145\
        );

    \I__5854\ : LocalMux
    port map (
            O => \N__31145\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9\
        );

    \I__5853\ : InMux
    port map (
            O => \N__31142\,
            I => \N__31139\
        );

    \I__5852\ : LocalMux
    port map (
            O => \N__31139\,
            I => \N__31135\
        );

    \I__5851\ : InMux
    port map (
            O => \N__31138\,
            I => \N__31132\
        );

    \I__5850\ : Span4Mux_v
    port map (
            O => \N__31135\,
            I => \N__31129\
        );

    \I__5849\ : LocalMux
    port map (
            O => \N__31132\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__5848\ : Odrv4
    port map (
            O => \N__31129\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__5847\ : CascadeMux
    port map (
            O => \N__31124\,
            I => \phase_controller_inst1.start_timer_hc_0_sqmuxa_cascade_\
        );

    \I__5846\ : InMux
    port map (
            O => \N__31121\,
            I => \N__31118\
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__31118\,
            I => \phase_controller_inst1.N_88\
        );

    \I__5844\ : InMux
    port map (
            O => \N__31115\,
            I => \N__31112\
        );

    \I__5843\ : LocalMux
    port map (
            O => \N__31112\,
            I => \N__31107\
        );

    \I__5842\ : InMux
    port map (
            O => \N__31111\,
            I => \N__31101\
        );

    \I__5841\ : InMux
    port map (
            O => \N__31110\,
            I => \N__31101\
        );

    \I__5840\ : Span4Mux_h
    port map (
            O => \N__31107\,
            I => \N__31098\
        );

    \I__5839\ : InMux
    port map (
            O => \N__31106\,
            I => \N__31095\
        );

    \I__5838\ : LocalMux
    port map (
            O => \N__31101\,
            I => \N__31092\
        );

    \I__5837\ : Odrv4
    port map (
            O => \N__31098\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__5836\ : LocalMux
    port map (
            O => \N__31095\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__5835\ : Odrv4
    port map (
            O => \N__31092\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__5834\ : InMux
    port map (
            O => \N__31085\,
            I => \N__31082\
        );

    \I__5833\ : LocalMux
    port map (
            O => \N__31082\,
            I => \N__31079\
        );

    \I__5832\ : Odrv4
    port map (
            O => \N__31079\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIDR081_20\
        );

    \I__5831\ : CascadeMux
    port map (
            O => \N__31076\,
            I => \N__31073\
        );

    \I__5830\ : InMux
    port map (
            O => \N__31073\,
            I => \N__31067\
        );

    \I__5829\ : InMux
    port map (
            O => \N__31072\,
            I => \N__31062\
        );

    \I__5828\ : InMux
    port map (
            O => \N__31071\,
            I => \N__31062\
        );

    \I__5827\ : CascadeMux
    port map (
            O => \N__31070\,
            I => \N__31059\
        );

    \I__5826\ : LocalMux
    port map (
            O => \N__31067\,
            I => \N__31054\
        );

    \I__5825\ : LocalMux
    port map (
            O => \N__31062\,
            I => \N__31054\
        );

    \I__5824\ : InMux
    port map (
            O => \N__31059\,
            I => \N__31051\
        );

    \I__5823\ : Odrv4
    port map (
            O => \N__31054\,
            I => \current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0\
        );

    \I__5822\ : LocalMux
    port map (
            O => \N__31051\,
            I => \current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0\
        );

    \I__5821\ : CascadeMux
    port map (
            O => \N__31046\,
            I => \N__31042\
        );

    \I__5820\ : InMux
    port map (
            O => \N__31045\,
            I => \N__31034\
        );

    \I__5819\ : InMux
    port map (
            O => \N__31042\,
            I => \N__31034\
        );

    \I__5818\ : InMux
    port map (
            O => \N__31041\,
            I => \N__31034\
        );

    \I__5817\ : LocalMux
    port map (
            O => \N__31034\,
            I => \N__31030\
        );

    \I__5816\ : InMux
    port map (
            O => \N__31033\,
            I => \N__31027\
        );

    \I__5815\ : Span4Mux_h
    port map (
            O => \N__31030\,
            I => \N__31022\
        );

    \I__5814\ : LocalMux
    port map (
            O => \N__31027\,
            I => \N__31022\
        );

    \I__5813\ : Odrv4
    port map (
            O => \N__31022\,
            I => \current_shift_inst.elapsed_time_ns_phase_20\
        );

    \I__5812\ : CascadeMux
    port map (
            O => \N__31019\,
            I => \N__31016\
        );

    \I__5811\ : InMux
    port map (
            O => \N__31016\,
            I => \N__31013\
        );

    \I__5810\ : LocalMux
    port map (
            O => \N__31013\,
            I => \N__31010\
        );

    \I__5809\ : Odrv4
    port map (
            O => \N__31010\,
            I => \current_shift_inst.elapsed_time_ns_1_RNILRVJ_20\
        );

    \I__5808\ : CascadeMux
    port map (
            O => \N__31007\,
            I => \N__31004\
        );

    \I__5807\ : InMux
    port map (
            O => \N__31004\,
            I => \N__30999\
        );

    \I__5806\ : InMux
    port map (
            O => \N__31003\,
            I => \N__30996\
        );

    \I__5805\ : InMux
    port map (
            O => \N__31002\,
            I => \N__30993\
        );

    \I__5804\ : LocalMux
    port map (
            O => \N__30999\,
            I => \N__30989\
        );

    \I__5803\ : LocalMux
    port map (
            O => \N__30996\,
            I => \N__30984\
        );

    \I__5802\ : LocalMux
    port map (
            O => \N__30993\,
            I => \N__30984\
        );

    \I__5801\ : InMux
    port map (
            O => \N__30992\,
            I => \N__30981\
        );

    \I__5800\ : Span4Mux_v
    port map (
            O => \N__30989\,
            I => \N__30978\
        );

    \I__5799\ : Span4Mux_h
    port map (
            O => \N__30984\,
            I => \N__30973\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__30981\,
            I => \N__30973\
        );

    \I__5797\ : Odrv4
    port map (
            O => \N__30978\,
            I => \current_shift_inst.elapsed_time_ns_phase_21\
        );

    \I__5796\ : Odrv4
    port map (
            O => \N__30973\,
            I => \current_shift_inst.elapsed_time_ns_phase_21\
        );

    \I__5795\ : InMux
    port map (
            O => \N__30968\,
            I => \N__30965\
        );

    \I__5794\ : LocalMux
    port map (
            O => \N__30965\,
            I => \N__30960\
        );

    \I__5793\ : InMux
    port map (
            O => \N__30964\,
            I => \N__30955\
        );

    \I__5792\ : InMux
    port map (
            O => \N__30963\,
            I => \N__30955\
        );

    \I__5791\ : Span4Mux_v
    port map (
            O => \N__30960\,
            I => \N__30951\
        );

    \I__5790\ : LocalMux
    port map (
            O => \N__30955\,
            I => \N__30948\
        );

    \I__5789\ : InMux
    port map (
            O => \N__30954\,
            I => \N__30945\
        );

    \I__5788\ : Odrv4
    port map (
            O => \N__30951\,
            I => \current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0\
        );

    \I__5787\ : Odrv4
    port map (
            O => \N__30948\,
            I => \current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0\
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__30945\,
            I => \current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0\
        );

    \I__5785\ : CascadeMux
    port map (
            O => \N__30938\,
            I => \N__30935\
        );

    \I__5784\ : InMux
    port map (
            O => \N__30935\,
            I => \N__30932\
        );

    \I__5783\ : LocalMux
    port map (
            O => \N__30932\,
            I => \N__30929\
        );

    \I__5782\ : Span4Mux_h
    port map (
            O => \N__30929\,
            I => \N__30926\
        );

    \I__5781\ : Odrv4
    port map (
            O => \N__30926\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIOV0K_21\
        );

    \I__5780\ : CascadeMux
    port map (
            O => \N__30923\,
            I => \N__30920\
        );

    \I__5779\ : InMux
    port map (
            O => \N__30920\,
            I => \N__30917\
        );

    \I__5778\ : LocalMux
    port map (
            O => \N__30917\,
            I => \N__30914\
        );

    \I__5777\ : Odrv12
    port map (
            O => \N__30914\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIU73K_23\
        );

    \I__5776\ : CascadeMux
    port map (
            O => \N__30911\,
            I => \N__30908\
        );

    \I__5775\ : InMux
    port map (
            O => \N__30908\,
            I => \N__30905\
        );

    \I__5774\ : LocalMux
    port map (
            O => \N__30905\,
            I => \N__30902\
        );

    \I__5773\ : Odrv12
    port map (
            O => \N__30902\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI7K6K_26\
        );

    \I__5772\ : InMux
    port map (
            O => \N__30899\,
            I => \N__30896\
        );

    \I__5771\ : LocalMux
    port map (
            O => \N__30896\,
            I => \N__30893\
        );

    \I__5770\ : Span12Mux_v
    port map (
            O => \N__30893\,
            I => \N__30890\
        );

    \I__5769\ : Span12Mux_v
    port map (
            O => \N__30890\,
            I => \N__30887\
        );

    \I__5768\ : Odrv12
    port map (
            O => \N__30887\,
            I => \il_max_comp2_D1\
        );

    \I__5767\ : InMux
    port map (
            O => \N__30884\,
            I => \N__30880\
        );

    \I__5766\ : InMux
    port map (
            O => \N__30883\,
            I => \N__30876\
        );

    \I__5765\ : LocalMux
    port map (
            O => \N__30880\,
            I => \N__30873\
        );

    \I__5764\ : InMux
    port map (
            O => \N__30879\,
            I => \N__30870\
        );

    \I__5763\ : LocalMux
    port map (
            O => \N__30876\,
            I => \N__30864\
        );

    \I__5762\ : Span4Mux_h
    port map (
            O => \N__30873\,
            I => \N__30864\
        );

    \I__5761\ : LocalMux
    port map (
            O => \N__30870\,
            I => \N__30861\
        );

    \I__5760\ : InMux
    port map (
            O => \N__30869\,
            I => \N__30858\
        );

    \I__5759\ : Span4Mux_v
    port map (
            O => \N__30864\,
            I => \N__30855\
        );

    \I__5758\ : Span4Mux_v
    port map (
            O => \N__30861\,
            I => \N__30852\
        );

    \I__5757\ : LocalMux
    port map (
            O => \N__30858\,
            I => \N__30849\
        );

    \I__5756\ : Odrv4
    port map (
            O => \N__30855\,
            I => \current_shift_inst.elapsed_time_ns_phase_28\
        );

    \I__5755\ : Odrv4
    port map (
            O => \N__30852\,
            I => \current_shift_inst.elapsed_time_ns_phase_28\
        );

    \I__5754\ : Odrv4
    port map (
            O => \N__30849\,
            I => \current_shift_inst.elapsed_time_ns_phase_28\
        );

    \I__5753\ : CascadeMux
    port map (
            O => \N__30842\,
            I => \N__30839\
        );

    \I__5752\ : InMux
    port map (
            O => \N__30839\,
            I => \N__30835\
        );

    \I__5751\ : InMux
    port map (
            O => \N__30838\,
            I => \N__30832\
        );

    \I__5750\ : LocalMux
    port map (
            O => \N__30835\,
            I => \N__30828\
        );

    \I__5749\ : LocalMux
    port map (
            O => \N__30832\,
            I => \N__30824\
        );

    \I__5748\ : CascadeMux
    port map (
            O => \N__30831\,
            I => \N__30821\
        );

    \I__5747\ : Span4Mux_v
    port map (
            O => \N__30828\,
            I => \N__30818\
        );

    \I__5746\ : InMux
    port map (
            O => \N__30827\,
            I => \N__30815\
        );

    \I__5745\ : Span4Mux_h
    port map (
            O => \N__30824\,
            I => \N__30812\
        );

    \I__5744\ : InMux
    port map (
            O => \N__30821\,
            I => \N__30809\
        );

    \I__5743\ : Odrv4
    port map (
            O => \N__30818\,
            I => \current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0\
        );

    \I__5742\ : LocalMux
    port map (
            O => \N__30815\,
            I => \current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0\
        );

    \I__5741\ : Odrv4
    port map (
            O => \N__30812\,
            I => \current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0\
        );

    \I__5740\ : LocalMux
    port map (
            O => \N__30809\,
            I => \current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0\
        );

    \I__5739\ : CascadeMux
    port map (
            O => \N__30800\,
            I => \N__30797\
        );

    \I__5738\ : InMux
    port map (
            O => \N__30797\,
            I => \N__30794\
        );

    \I__5737\ : LocalMux
    port map (
            O => \N__30794\,
            I => \N__30791\
        );

    \I__5736\ : Span4Mux_v
    port map (
            O => \N__30791\,
            I => \N__30788\
        );

    \I__5735\ : Odrv4
    port map (
            O => \N__30788\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIDS8K_28\
        );

    \I__5734\ : InMux
    port map (
            O => \N__30785\,
            I => \N__30782\
        );

    \I__5733\ : LocalMux
    port map (
            O => \N__30782\,
            I => \N__30779\
        );

    \I__5732\ : Span4Mux_h
    port map (
            O => \N__30779\,
            I => \N__30776\
        );

    \I__5731\ : Odrv4
    port map (
            O => \N__30776\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5S981_24\
        );

    \I__5730\ : CascadeMux
    port map (
            O => \N__30773\,
            I => \N__30768\
        );

    \I__5729\ : InMux
    port map (
            O => \N__30772\,
            I => \N__30763\
        );

    \I__5728\ : InMux
    port map (
            O => \N__30771\,
            I => \N__30763\
        );

    \I__5727\ : InMux
    port map (
            O => \N__30768\,
            I => \N__30759\
        );

    \I__5726\ : LocalMux
    port map (
            O => \N__30763\,
            I => \N__30756\
        );

    \I__5725\ : InMux
    port map (
            O => \N__30762\,
            I => \N__30753\
        );

    \I__5724\ : LocalMux
    port map (
            O => \N__30759\,
            I => \N__30750\
        );

    \I__5723\ : Span4Mux_h
    port map (
            O => \N__30756\,
            I => \N__30745\
        );

    \I__5722\ : LocalMux
    port map (
            O => \N__30753\,
            I => \N__30745\
        );

    \I__5721\ : Odrv12
    port map (
            O => \N__30750\,
            I => \current_shift_inst.elapsed_time_ns_phase_11\
        );

    \I__5720\ : Odrv4
    port map (
            O => \N__30745\,
            I => \current_shift_inst.elapsed_time_ns_phase_11\
        );

    \I__5719\ : InMux
    port map (
            O => \N__30740\,
            I => \N__30730\
        );

    \I__5718\ : InMux
    port map (
            O => \N__30739\,
            I => \N__30730\
        );

    \I__5717\ : InMux
    port map (
            O => \N__30738\,
            I => \N__30730\
        );

    \I__5716\ : CascadeMux
    port map (
            O => \N__30737\,
            I => \N__30727\
        );

    \I__5715\ : LocalMux
    port map (
            O => \N__30730\,
            I => \N__30724\
        );

    \I__5714\ : InMux
    port map (
            O => \N__30727\,
            I => \N__30721\
        );

    \I__5713\ : Odrv4
    port map (
            O => \N__30724\,
            I => \current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0\
        );

    \I__5712\ : LocalMux
    port map (
            O => \N__30721\,
            I => \current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0\
        );

    \I__5711\ : CascadeMux
    port map (
            O => \N__30716\,
            I => \N__30712\
        );

    \I__5710\ : InMux
    port map (
            O => \N__30715\,
            I => \N__30709\
        );

    \I__5709\ : InMux
    port map (
            O => \N__30712\,
            I => \N__30704\
        );

    \I__5708\ : LocalMux
    port map (
            O => \N__30709\,
            I => \N__30701\
        );

    \I__5707\ : InMux
    port map (
            O => \N__30708\,
            I => \N__30698\
        );

    \I__5706\ : CascadeMux
    port map (
            O => \N__30707\,
            I => \N__30695\
        );

    \I__5705\ : LocalMux
    port map (
            O => \N__30704\,
            I => \N__30688\
        );

    \I__5704\ : Span4Mux_h
    port map (
            O => \N__30701\,
            I => \N__30688\
        );

    \I__5703\ : LocalMux
    port map (
            O => \N__30698\,
            I => \N__30688\
        );

    \I__5702\ : InMux
    port map (
            O => \N__30695\,
            I => \N__30685\
        );

    \I__5701\ : Odrv4
    port map (
            O => \N__30688\,
            I => \current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0\
        );

    \I__5700\ : LocalMux
    port map (
            O => \N__30685\,
            I => \current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0\
        );

    \I__5699\ : CascadeMux
    port map (
            O => \N__30680\,
            I => \N__30676\
        );

    \I__5698\ : CascadeMux
    port map (
            O => \N__30679\,
            I => \N__30673\
        );

    \I__5697\ : InMux
    port map (
            O => \N__30676\,
            I => \N__30669\
        );

    \I__5696\ : InMux
    port map (
            O => \N__30673\,
            I => \N__30664\
        );

    \I__5695\ : InMux
    port map (
            O => \N__30672\,
            I => \N__30664\
        );

    \I__5694\ : LocalMux
    port map (
            O => \N__30669\,
            I => \N__30658\
        );

    \I__5693\ : LocalMux
    port map (
            O => \N__30664\,
            I => \N__30658\
        );

    \I__5692\ : InMux
    port map (
            O => \N__30663\,
            I => \N__30655\
        );

    \I__5691\ : Span4Mux_h
    port map (
            O => \N__30658\,
            I => \N__30650\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__30655\,
            I => \N__30650\
        );

    \I__5689\ : Odrv4
    port map (
            O => \N__30650\,
            I => \current_shift_inst.elapsed_time_ns_phase_12\
        );

    \I__5688\ : InMux
    port map (
            O => \N__30647\,
            I => \N__30644\
        );

    \I__5687\ : LocalMux
    port map (
            O => \N__30644\,
            I => \N__30641\
        );

    \I__5686\ : Odrv4
    port map (
            O => \N__30641\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIDLO51_11\
        );

    \I__5685\ : InMux
    port map (
            O => \N__30638\,
            I => \N__30635\
        );

    \I__5684\ : LocalMux
    port map (
            O => \N__30635\,
            I => \N__30632\
        );

    \I__5683\ : Span4Mux_v
    port map (
            O => \N__30632\,
            I => \N__30627\
        );

    \I__5682\ : InMux
    port map (
            O => \N__30631\,
            I => \N__30624\
        );

    \I__5681\ : InMux
    port map (
            O => \N__30630\,
            I => \N__30621\
        );

    \I__5680\ : Span4Mux_v
    port map (
            O => \N__30627\,
            I => \N__30618\
        );

    \I__5679\ : LocalMux
    port map (
            O => \N__30624\,
            I => \N__30615\
        );

    \I__5678\ : LocalMux
    port map (
            O => \N__30621\,
            I => \N__30612\
        );

    \I__5677\ : Odrv4
    port map (
            O => \N__30618\,
            I => \current_shift_inst.elapsed_time_ns_phase_30\
        );

    \I__5676\ : Odrv12
    port map (
            O => \N__30615\,
            I => \current_shift_inst.elapsed_time_ns_phase_30\
        );

    \I__5675\ : Odrv4
    port map (
            O => \N__30612\,
            I => \current_shift_inst.elapsed_time_ns_phase_30\
        );

    \I__5674\ : CascadeMux
    port map (
            O => \N__30605\,
            I => \N__30600\
        );

    \I__5673\ : CascadeMux
    port map (
            O => \N__30604\,
            I => \N__30595\
        );

    \I__5672\ : CascadeMux
    port map (
            O => \N__30603\,
            I => \N__30591\
        );

    \I__5671\ : InMux
    port map (
            O => \N__30600\,
            I => \N__30587\
        );

    \I__5670\ : InMux
    port map (
            O => \N__30599\,
            I => \N__30584\
        );

    \I__5669\ : InMux
    port map (
            O => \N__30598\,
            I => \N__30575\
        );

    \I__5668\ : InMux
    port map (
            O => \N__30595\,
            I => \N__30575\
        );

    \I__5667\ : InMux
    port map (
            O => \N__30594\,
            I => \N__30575\
        );

    \I__5666\ : InMux
    port map (
            O => \N__30591\,
            I => \N__30575\
        );

    \I__5665\ : InMux
    port map (
            O => \N__30590\,
            I => \N__30571\
        );

    \I__5664\ : LocalMux
    port map (
            O => \N__30587\,
            I => \N__30564\
        );

    \I__5663\ : LocalMux
    port map (
            O => \N__30584\,
            I => \N__30564\
        );

    \I__5662\ : LocalMux
    port map (
            O => \N__30575\,
            I => \N__30564\
        );

    \I__5661\ : InMux
    port map (
            O => \N__30574\,
            I => \N__30561\
        );

    \I__5660\ : LocalMux
    port map (
            O => \N__30571\,
            I => \N__30557\
        );

    \I__5659\ : Span4Mux_h
    port map (
            O => \N__30564\,
            I => \N__30554\
        );

    \I__5658\ : LocalMux
    port map (
            O => \N__30561\,
            I => \N__30551\
        );

    \I__5657\ : InMux
    port map (
            O => \N__30560\,
            I => \N__30548\
        );

    \I__5656\ : Span4Mux_v
    port map (
            O => \N__30557\,
            I => \N__30539\
        );

    \I__5655\ : Span4Mux_h
    port map (
            O => \N__30554\,
            I => \N__30539\
        );

    \I__5654\ : Span4Mux_h
    port map (
            O => \N__30551\,
            I => \N__30539\
        );

    \I__5653\ : LocalMux
    port map (
            O => \N__30548\,
            I => \N__30539\
        );

    \I__5652\ : Span4Mux_v
    port map (
            O => \N__30539\,
            I => \N__30536\
        );

    \I__5651\ : Odrv4
    port map (
            O => \N__30536\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__5650\ : CascadeMux
    port map (
            O => \N__30533\,
            I => \N__30530\
        );

    \I__5649\ : InMux
    port map (
            O => \N__30530\,
            I => \N__30526\
        );

    \I__5648\ : CascadeMux
    port map (
            O => \N__30529\,
            I => \N__30523\
        );

    \I__5647\ : LocalMux
    port map (
            O => \N__30526\,
            I => \N__30520\
        );

    \I__5646\ : InMux
    port map (
            O => \N__30523\,
            I => \N__30517\
        );

    \I__5645\ : Span4Mux_h
    port map (
            O => \N__30520\,
            I => \N__30514\
        );

    \I__5644\ : LocalMux
    port map (
            O => \N__30517\,
            I => \N__30511\
        );

    \I__5643\ : Span4Mux_v
    port map (
            O => \N__30514\,
            I => \N__30508\
        );

    \I__5642\ : Span4Mux_v
    port map (
            O => \N__30511\,
            I => \N__30505\
        );

    \I__5641\ : Odrv4
    port map (
            O => \N__30508\,
            I => \current_shift_inst.elapsed_time_ns_phase_31\
        );

    \I__5640\ : Odrv4
    port map (
            O => \N__30505\,
            I => \current_shift_inst.elapsed_time_ns_phase_31\
        );

    \I__5639\ : InMux
    port map (
            O => \N__30500\,
            I => \N__30496\
        );

    \I__5638\ : InMux
    port map (
            O => \N__30499\,
            I => \N__30493\
        );

    \I__5637\ : LocalMux
    port map (
            O => \N__30496\,
            I => \N__30490\
        );

    \I__5636\ : LocalMux
    port map (
            O => \N__30493\,
            I => \N__30484\
        );

    \I__5635\ : Span4Mux_h
    port map (
            O => \N__30490\,
            I => \N__30484\
        );

    \I__5634\ : InMux
    port map (
            O => \N__30489\,
            I => \N__30481\
        );

    \I__5633\ : Odrv4
    port map (
            O => \N__30484\,
            I => \current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0\
        );

    \I__5632\ : LocalMux
    port map (
            O => \N__30481\,
            I => \current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0\
        );

    \I__5631\ : InMux
    port map (
            O => \N__30476\,
            I => \N__30473\
        );

    \I__5630\ : LocalMux
    port map (
            O => \N__30473\,
            I => \N__30470\
        );

    \I__5629\ : Span4Mux_h
    port map (
            O => \N__30470\,
            I => \N__30467\
        );

    \I__5628\ : Odrv4
    port map (
            O => \N__30467\,
            I => \current_shift_inst.un38_control_input_0_axb_31\
        );

    \I__5627\ : InMux
    port map (
            O => \N__30464\,
            I => \N__30459\
        );

    \I__5626\ : InMux
    port map (
            O => \N__30463\,
            I => \N__30456\
        );

    \I__5625\ : InMux
    port map (
            O => \N__30462\,
            I => \N__30453\
        );

    \I__5624\ : LocalMux
    port map (
            O => \N__30459\,
            I => \N__30449\
        );

    \I__5623\ : LocalMux
    port map (
            O => \N__30456\,
            I => \N__30446\
        );

    \I__5622\ : LocalMux
    port map (
            O => \N__30453\,
            I => \N__30443\
        );

    \I__5621\ : InMux
    port map (
            O => \N__30452\,
            I => \N__30440\
        );

    \I__5620\ : Span4Mux_h
    port map (
            O => \N__30449\,
            I => \N__30435\
        );

    \I__5619\ : Span4Mux_v
    port map (
            O => \N__30446\,
            I => \N__30435\
        );

    \I__5618\ : Span4Mux_v
    port map (
            O => \N__30443\,
            I => \N__30430\
        );

    \I__5617\ : LocalMux
    port map (
            O => \N__30440\,
            I => \N__30430\
        );

    \I__5616\ : Odrv4
    port map (
            O => \N__30435\,
            I => \current_shift_inst.elapsed_time_ns_phase_19\
        );

    \I__5615\ : Odrv4
    port map (
            O => \N__30430\,
            I => \current_shift_inst.elapsed_time_ns_phase_19\
        );

    \I__5614\ : CascadeMux
    port map (
            O => \N__30425\,
            I => \N__30421\
        );

    \I__5613\ : InMux
    port map (
            O => \N__30424\,
            I => \N__30418\
        );

    \I__5612\ : InMux
    port map (
            O => \N__30421\,
            I => \N__30413\
        );

    \I__5611\ : LocalMux
    port map (
            O => \N__30418\,
            I => \N__30410\
        );

    \I__5610\ : InMux
    port map (
            O => \N__30417\,
            I => \N__30407\
        );

    \I__5609\ : CascadeMux
    port map (
            O => \N__30416\,
            I => \N__30404\
        );

    \I__5608\ : LocalMux
    port map (
            O => \N__30413\,
            I => \N__30401\
        );

    \I__5607\ : Span4Mux_v
    port map (
            O => \N__30410\,
            I => \N__30398\
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__30407\,
            I => \N__30395\
        );

    \I__5605\ : InMux
    port map (
            O => \N__30404\,
            I => \N__30392\
        );

    \I__5604\ : Odrv12
    port map (
            O => \N__30401\,
            I => \current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0\
        );

    \I__5603\ : Odrv4
    port map (
            O => \N__30398\,
            I => \current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0\
        );

    \I__5602\ : Odrv4
    port map (
            O => \N__30395\,
            I => \current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0\
        );

    \I__5601\ : LocalMux
    port map (
            O => \N__30392\,
            I => \current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0\
        );

    \I__5600\ : InMux
    port map (
            O => \N__30383\,
            I => \N__30380\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__30380\,
            I => \N__30377\
        );

    \I__5598\ : Odrv12
    port map (
            O => \N__30377\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPC571_19\
        );

    \I__5597\ : CascadeMux
    port map (
            O => \N__30374\,
            I => \N__30371\
        );

    \I__5596\ : InMux
    port map (
            O => \N__30371\,
            I => \N__30368\
        );

    \I__5595\ : LocalMux
    port map (
            O => \N__30368\,
            I => \N__30365\
        );

    \I__5594\ : Span4Mux_h
    port map (
            O => \N__30365\,
            I => \N__30362\
        );

    \I__5593\ : Odrv4
    port map (
            O => \N__30362\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI190J_15\
        );

    \I__5592\ : InMux
    port map (
            O => \N__30359\,
            I => \N__30354\
        );

    \I__5591\ : CascadeMux
    port map (
            O => \N__30358\,
            I => \N__30351\
        );

    \I__5590\ : CascadeMux
    port map (
            O => \N__30357\,
            I => \N__30347\
        );

    \I__5589\ : LocalMux
    port map (
            O => \N__30354\,
            I => \N__30344\
        );

    \I__5588\ : InMux
    port map (
            O => \N__30351\,
            I => \N__30341\
        );

    \I__5587\ : InMux
    port map (
            O => \N__30350\,
            I => \N__30338\
        );

    \I__5586\ : InMux
    port map (
            O => \N__30347\,
            I => \N__30335\
        );

    \I__5585\ : Span4Mux_v
    port map (
            O => \N__30344\,
            I => \N__30332\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__30341\,
            I => \N__30325\
        );

    \I__5583\ : LocalMux
    port map (
            O => \N__30338\,
            I => \N__30325\
        );

    \I__5582\ : LocalMux
    port map (
            O => \N__30335\,
            I => \N__30325\
        );

    \I__5581\ : Odrv4
    port map (
            O => \N__30332\,
            I => \current_shift_inst.elapsed_time_ns_phase_16\
        );

    \I__5580\ : Odrv4
    port map (
            O => \N__30325\,
            I => \current_shift_inst.elapsed_time_ns_phase_16\
        );

    \I__5579\ : InMux
    port map (
            O => \N__30320\,
            I => \N__30316\
        );

    \I__5578\ : InMux
    port map (
            O => \N__30319\,
            I => \N__30313\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__30316\,
            I => \N__30307\
        );

    \I__5576\ : LocalMux
    port map (
            O => \N__30313\,
            I => \N__30307\
        );

    \I__5575\ : InMux
    port map (
            O => \N__30312\,
            I => \N__30304\
        );

    \I__5574\ : Span4Mux_v
    port map (
            O => \N__30307\,
            I => \N__30300\
        );

    \I__5573\ : LocalMux
    port map (
            O => \N__30304\,
            I => \N__30297\
        );

    \I__5572\ : InMux
    port map (
            O => \N__30303\,
            I => \N__30294\
        );

    \I__5571\ : Odrv4
    port map (
            O => \N__30300\,
            I => \current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0\
        );

    \I__5570\ : Odrv12
    port map (
            O => \N__30297\,
            I => \current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0\
        );

    \I__5569\ : LocalMux
    port map (
            O => \N__30294\,
            I => \current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0\
        );

    \I__5568\ : InMux
    port map (
            O => \N__30287\,
            I => \N__30284\
        );

    \I__5567\ : LocalMux
    port map (
            O => \N__30284\,
            I => \N__30281\
        );

    \I__5566\ : Odrv4
    port map (
            O => \N__30281\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5M161_15\
        );

    \I__5565\ : InMux
    port map (
            O => \N__30278\,
            I => \N__30275\
        );

    \I__5564\ : LocalMux
    port map (
            O => \N__30275\,
            I => \N__30272\
        );

    \I__5563\ : Span4Mux_h
    port map (
            O => \N__30272\,
            I => \N__30266\
        );

    \I__5562\ : InMux
    port map (
            O => \N__30271\,
            I => \N__30263\
        );

    \I__5561\ : InMux
    port map (
            O => \N__30270\,
            I => \N__30260\
        );

    \I__5560\ : InMux
    port map (
            O => \N__30269\,
            I => \N__30257\
        );

    \I__5559\ : Span4Mux_h
    port map (
            O => \N__30266\,
            I => \N__30254\
        );

    \I__5558\ : LocalMux
    port map (
            O => \N__30263\,
            I => \N__30251\
        );

    \I__5557\ : LocalMux
    port map (
            O => \N__30260\,
            I => \N__30246\
        );

    \I__5556\ : LocalMux
    port map (
            O => \N__30257\,
            I => \N__30246\
        );

    \I__5555\ : Odrv4
    port map (
            O => \N__30254\,
            I => \current_shift_inst.elapsed_time_ns_phase_14\
        );

    \I__5554\ : Odrv12
    port map (
            O => \N__30251\,
            I => \current_shift_inst.elapsed_time_ns_phase_14\
        );

    \I__5553\ : Odrv4
    port map (
            O => \N__30246\,
            I => \current_shift_inst.elapsed_time_ns_phase_14\
        );

    \I__5552\ : CascadeMux
    port map (
            O => \N__30239\,
            I => \N__30236\
        );

    \I__5551\ : InMux
    port map (
            O => \N__30236\,
            I => \N__30226\
        );

    \I__5550\ : InMux
    port map (
            O => \N__30235\,
            I => \N__30226\
        );

    \I__5549\ : InMux
    port map (
            O => \N__30234\,
            I => \N__30226\
        );

    \I__5548\ : CascadeMux
    port map (
            O => \N__30233\,
            I => \N__30223\
        );

    \I__5547\ : LocalMux
    port map (
            O => \N__30226\,
            I => \N__30220\
        );

    \I__5546\ : InMux
    port map (
            O => \N__30223\,
            I => \N__30217\
        );

    \I__5545\ : Odrv12
    port map (
            O => \N__30220\,
            I => \current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0\
        );

    \I__5544\ : LocalMux
    port map (
            O => \N__30217\,
            I => \current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0\
        );

    \I__5543\ : CascadeMux
    port map (
            O => \N__30212\,
            I => \N__30208\
        );

    \I__5542\ : InMux
    port map (
            O => \N__30211\,
            I => \N__30204\
        );

    \I__5541\ : InMux
    port map (
            O => \N__30208\,
            I => \N__30201\
        );

    \I__5540\ : InMux
    port map (
            O => \N__30207\,
            I => \N__30198\
        );

    \I__5539\ : LocalMux
    port map (
            O => \N__30204\,
            I => \N__30194\
        );

    \I__5538\ : LocalMux
    port map (
            O => \N__30201\,
            I => \N__30191\
        );

    \I__5537\ : LocalMux
    port map (
            O => \N__30198\,
            I => \N__30188\
        );

    \I__5536\ : CascadeMux
    port map (
            O => \N__30197\,
            I => \N__30185\
        );

    \I__5535\ : Span4Mux_v
    port map (
            O => \N__30194\,
            I => \N__30182\
        );

    \I__5534\ : Span4Mux_v
    port map (
            O => \N__30191\,
            I => \N__30177\
        );

    \I__5533\ : Span4Mux_h
    port map (
            O => \N__30188\,
            I => \N__30177\
        );

    \I__5532\ : InMux
    port map (
            O => \N__30185\,
            I => \N__30174\
        );

    \I__5531\ : Odrv4
    port map (
            O => \N__30182\,
            I => \current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0\
        );

    \I__5530\ : Odrv4
    port map (
            O => \N__30177\,
            I => \current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0\
        );

    \I__5529\ : LocalMux
    port map (
            O => \N__30174\,
            I => \current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0\
        );

    \I__5528\ : InMux
    port map (
            O => \N__30167\,
            I => \N__30157\
        );

    \I__5527\ : InMux
    port map (
            O => \N__30166\,
            I => \N__30157\
        );

    \I__5526\ : InMux
    port map (
            O => \N__30165\,
            I => \N__30157\
        );

    \I__5525\ : InMux
    port map (
            O => \N__30164\,
            I => \N__30154\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__30157\,
            I => \N__30151\
        );

    \I__5523\ : LocalMux
    port map (
            O => \N__30154\,
            I => \N__30148\
        );

    \I__5522\ : Span4Mux_v
    port map (
            O => \N__30151\,
            I => \N__30145\
        );

    \I__5521\ : Span4Mux_v
    port map (
            O => \N__30148\,
            I => \N__30142\
        );

    \I__5520\ : Odrv4
    port map (
            O => \N__30145\,
            I => \current_shift_inst.elapsed_time_ns_phase_15\
        );

    \I__5519\ : Odrv4
    port map (
            O => \N__30142\,
            I => \current_shift_inst.elapsed_time_ns_phase_15\
        );

    \I__5518\ : InMux
    port map (
            O => \N__30137\,
            I => \N__30134\
        );

    \I__5517\ : LocalMux
    port map (
            O => \N__30134\,
            I => \N__30131\
        );

    \I__5516\ : Odrv4
    port map (
            O => \N__30131\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIVDV51_14\
        );

    \I__5515\ : CascadeMux
    port map (
            O => \N__30128\,
            I => \N__30125\
        );

    \I__5514\ : InMux
    port map (
            O => \N__30125\,
            I => \N__30122\
        );

    \I__5513\ : LocalMux
    port map (
            O => \N__30122\,
            I => \N__30117\
        );

    \I__5512\ : InMux
    port map (
            O => \N__30121\,
            I => \N__30112\
        );

    \I__5511\ : InMux
    port map (
            O => \N__30120\,
            I => \N__30112\
        );

    \I__5510\ : Span4Mux_h
    port map (
            O => \N__30117\,
            I => \N__30108\
        );

    \I__5509\ : LocalMux
    port map (
            O => \N__30112\,
            I => \N__30105\
        );

    \I__5508\ : CascadeMux
    port map (
            O => \N__30111\,
            I => \N__30102\
        );

    \I__5507\ : Sp12to4
    port map (
            O => \N__30108\,
            I => \N__30099\
        );

    \I__5506\ : Span4Mux_h
    port map (
            O => \N__30105\,
            I => \N__30096\
        );

    \I__5505\ : InMux
    port map (
            O => \N__30102\,
            I => \N__30093\
        );

    \I__5504\ : Odrv12
    port map (
            O => \N__30099\,
            I => \current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0\
        );

    \I__5503\ : Odrv4
    port map (
            O => \N__30096\,
            I => \current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0\
        );

    \I__5502\ : LocalMux
    port map (
            O => \N__30093\,
            I => \current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0\
        );

    \I__5501\ : InMux
    port map (
            O => \N__30086\,
            I => \current_shift_inst.un4_control_input_cry_27\
        );

    \I__5500\ : InMux
    port map (
            O => \N__30083\,
            I => \current_shift_inst.un4_control_input_cry_28\
        );

    \I__5499\ : InMux
    port map (
            O => \N__30080\,
            I => \current_shift_inst.un4_control_input_cry_29\
        );

    \I__5498\ : InMux
    port map (
            O => \N__30077\,
            I => \current_shift_inst.un4_control_input_cry_30\
        );

    \I__5497\ : InMux
    port map (
            O => \N__30074\,
            I => \N__30070\
        );

    \I__5496\ : InMux
    port map (
            O => \N__30073\,
            I => \N__30066\
        );

    \I__5495\ : LocalMux
    port map (
            O => \N__30070\,
            I => \N__30062\
        );

    \I__5494\ : InMux
    port map (
            O => \N__30069\,
            I => \N__30059\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__30066\,
            I => \N__30056\
        );

    \I__5492\ : InMux
    port map (
            O => \N__30065\,
            I => \N__30053\
        );

    \I__5491\ : Span4Mux_h
    port map (
            O => \N__30062\,
            I => \N__30044\
        );

    \I__5490\ : LocalMux
    port map (
            O => \N__30059\,
            I => \N__30044\
        );

    \I__5489\ : Span4Mux_h
    port map (
            O => \N__30056\,
            I => \N__30044\
        );

    \I__5488\ : LocalMux
    port map (
            O => \N__30053\,
            I => \N__30044\
        );

    \I__5487\ : Odrv4
    port map (
            O => \N__30044\,
            I => \current_shift_inst.elapsed_time_ns_phase_9\
        );

    \I__5486\ : CascadeMux
    port map (
            O => \N__30041\,
            I => \N__30038\
        );

    \I__5485\ : InMux
    port map (
            O => \N__30038\,
            I => \N__30034\
        );

    \I__5484\ : InMux
    port map (
            O => \N__30037\,
            I => \N__30031\
        );

    \I__5483\ : LocalMux
    port map (
            O => \N__30034\,
            I => \N__30024\
        );

    \I__5482\ : LocalMux
    port map (
            O => \N__30031\,
            I => \N__30024\
        );

    \I__5481\ : InMux
    port map (
            O => \N__30030\,
            I => \N__30021\
        );

    \I__5480\ : CascadeMux
    port map (
            O => \N__30029\,
            I => \N__30018\
        );

    \I__5479\ : Span4Mux_v
    port map (
            O => \N__30024\,
            I => \N__30015\
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__30021\,
            I => \N__30012\
        );

    \I__5477\ : InMux
    port map (
            O => \N__30018\,
            I => \N__30009\
        );

    \I__5476\ : Odrv4
    port map (
            O => \N__30015\,
            I => \current_shift_inst.un4_control_input_cry_9_c_RNIALDJZ0\
        );

    \I__5475\ : Odrv12
    port map (
            O => \N__30012\,
            I => \current_shift_inst.un4_control_input_cry_9_c_RNIALDJZ0\
        );

    \I__5474\ : LocalMux
    port map (
            O => \N__30009\,
            I => \current_shift_inst.un4_control_input_cry_9_c_RNIALDJZ0\
        );

    \I__5473\ : InMux
    port map (
            O => \N__30002\,
            I => \N__29999\
        );

    \I__5472\ : LocalMux
    port map (
            O => \N__29999\,
            I => \N__29996\
        );

    \I__5471\ : Odrv12
    port map (
            O => \N__29996\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIO0U12_8\
        );

    \I__5470\ : CascadeMux
    port map (
            O => \N__29993\,
            I => \N__29990\
        );

    \I__5469\ : InMux
    port map (
            O => \N__29990\,
            I => \N__29987\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__29987\,
            I => \N__29984\
        );

    \I__5467\ : Odrv12
    port map (
            O => \N__29984\,
            I => \current_shift_inst.elapsed_time_ns_1_RNILORI_11\
        );

    \I__5466\ : CascadeMux
    port map (
            O => \N__29981\,
            I => \N__29978\
        );

    \I__5465\ : InMux
    port map (
            O => \N__29978\,
            I => \N__29975\
        );

    \I__5464\ : LocalMux
    port map (
            O => \N__29975\,
            I => \N__29972\
        );

    \I__5463\ : Odrv4
    port map (
            O => \N__29972\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIOSSI_12\
        );

    \I__5462\ : InMux
    port map (
            O => \N__29969\,
            I => \N__29964\
        );

    \I__5461\ : InMux
    port map (
            O => \N__29968\,
            I => \N__29961\
        );

    \I__5460\ : InMux
    port map (
            O => \N__29967\,
            I => \N__29958\
        );

    \I__5459\ : LocalMux
    port map (
            O => \N__29964\,
            I => \N__29952\
        );

    \I__5458\ : LocalMux
    port map (
            O => \N__29961\,
            I => \N__29952\
        );

    \I__5457\ : LocalMux
    port map (
            O => \N__29958\,
            I => \N__29949\
        );

    \I__5456\ : InMux
    port map (
            O => \N__29957\,
            I => \N__29946\
        );

    \I__5455\ : Span4Mux_v
    port map (
            O => \N__29952\,
            I => \N__29943\
        );

    \I__5454\ : Span4Mux_h
    port map (
            O => \N__29949\,
            I => \N__29938\
        );

    \I__5453\ : LocalMux
    port map (
            O => \N__29946\,
            I => \N__29938\
        );

    \I__5452\ : Odrv4
    port map (
            O => \N__29943\,
            I => \current_shift_inst.elapsed_time_ns_phase_13\
        );

    \I__5451\ : Odrv4
    port map (
            O => \N__29938\,
            I => \current_shift_inst.elapsed_time_ns_phase_13\
        );

    \I__5450\ : CascadeMux
    port map (
            O => \N__29933\,
            I => \N__29930\
        );

    \I__5449\ : InMux
    port map (
            O => \N__29930\,
            I => \N__29926\
        );

    \I__5448\ : InMux
    port map (
            O => \N__29929\,
            I => \N__29922\
        );

    \I__5447\ : LocalMux
    port map (
            O => \N__29926\,
            I => \N__29918\
        );

    \I__5446\ : InMux
    port map (
            O => \N__29925\,
            I => \N__29915\
        );

    \I__5445\ : LocalMux
    port map (
            O => \N__29922\,
            I => \N__29912\
        );

    \I__5444\ : CascadeMux
    port map (
            O => \N__29921\,
            I => \N__29909\
        );

    \I__5443\ : Span4Mux_h
    port map (
            O => \N__29918\,
            I => \N__29904\
        );

    \I__5442\ : LocalMux
    port map (
            O => \N__29915\,
            I => \N__29904\
        );

    \I__5441\ : Span4Mux_v
    port map (
            O => \N__29912\,
            I => \N__29901\
        );

    \I__5440\ : InMux
    port map (
            O => \N__29909\,
            I => \N__29898\
        );

    \I__5439\ : Odrv4
    port map (
            O => \N__29904\,
            I => \current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0\
        );

    \I__5438\ : Odrv4
    port map (
            O => \N__29901\,
            I => \current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__29898\,
            I => \current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0\
        );

    \I__5436\ : InMux
    port map (
            O => \N__29891\,
            I => \N__29888\
        );

    \I__5435\ : LocalMux
    port map (
            O => \N__29888\,
            I => \N__29885\
        );

    \I__5434\ : Odrv12
    port map (
            O => \N__29885\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJTQ51_12\
        );

    \I__5433\ : InMux
    port map (
            O => \N__29882\,
            I => \N__29877\
        );

    \I__5432\ : InMux
    port map (
            O => \N__29881\,
            I => \N__29874\
        );

    \I__5431\ : InMux
    port map (
            O => \N__29880\,
            I => \N__29870\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__29877\,
            I => \N__29865\
        );

    \I__5429\ : LocalMux
    port map (
            O => \N__29874\,
            I => \N__29865\
        );

    \I__5428\ : InMux
    port map (
            O => \N__29873\,
            I => \N__29862\
        );

    \I__5427\ : LocalMux
    port map (
            O => \N__29870\,
            I => \N__29859\
        );

    \I__5426\ : Span4Mux_v
    port map (
            O => \N__29865\,
            I => \N__29856\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__29862\,
            I => \N__29853\
        );

    \I__5424\ : Odrv4
    port map (
            O => \N__29859\,
            I => \current_shift_inst.elapsed_time_ns_phase_8\
        );

    \I__5423\ : Odrv4
    port map (
            O => \N__29856\,
            I => \current_shift_inst.elapsed_time_ns_phase_8\
        );

    \I__5422\ : Odrv4
    port map (
            O => \N__29853\,
            I => \current_shift_inst.elapsed_time_ns_phase_8\
        );

    \I__5421\ : InMux
    port map (
            O => \N__29846\,
            I => \N__29842\
        );

    \I__5420\ : CascadeMux
    port map (
            O => \N__29845\,
            I => \N__29839\
        );

    \I__5419\ : LocalMux
    port map (
            O => \N__29842\,
            I => \N__29834\
        );

    \I__5418\ : InMux
    port map (
            O => \N__29839\,
            I => \N__29831\
        );

    \I__5417\ : InMux
    port map (
            O => \N__29838\,
            I => \N__29828\
        );

    \I__5416\ : CascadeMux
    port map (
            O => \N__29837\,
            I => \N__29825\
        );

    \I__5415\ : Span4Mux_v
    port map (
            O => \N__29834\,
            I => \N__29822\
        );

    \I__5414\ : LocalMux
    port map (
            O => \N__29831\,
            I => \N__29817\
        );

    \I__5413\ : LocalMux
    port map (
            O => \N__29828\,
            I => \N__29817\
        );

    \I__5412\ : InMux
    port map (
            O => \N__29825\,
            I => \N__29814\
        );

    \I__5411\ : Odrv4
    port map (
            O => \N__29822\,
            I => \current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0\
        );

    \I__5410\ : Odrv12
    port map (
            O => \N__29817\,
            I => \current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0\
        );

    \I__5409\ : LocalMux
    port map (
            O => \N__29814\,
            I => \current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0\
        );

    \I__5408\ : CascadeMux
    port map (
            O => \N__29807\,
            I => \N__29804\
        );

    \I__5407\ : InMux
    port map (
            O => \N__29804\,
            I => \N__29801\
        );

    \I__5406\ : LocalMux
    port map (
            O => \N__29801\,
            I => \N__29798\
        );

    \I__5405\ : Odrv4
    port map (
            O => \N__29798\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIN7DV_8\
        );

    \I__5404\ : InMux
    port map (
            O => \N__29795\,
            I => \current_shift_inst.un4_control_input_cry_18\
        );

    \I__5403\ : InMux
    port map (
            O => \N__29792\,
            I => \current_shift_inst.un4_control_input_cry_19\
        );

    \I__5402\ : InMux
    port map (
            O => \N__29789\,
            I => \current_shift_inst.un4_control_input_cry_20\
        );

    \I__5401\ : InMux
    port map (
            O => \N__29786\,
            I => \current_shift_inst.un4_control_input_cry_21\
        );

    \I__5400\ : CascadeMux
    port map (
            O => \N__29783\,
            I => \N__29780\
        );

    \I__5399\ : InMux
    port map (
            O => \N__29780\,
            I => \N__29771\
        );

    \I__5398\ : InMux
    port map (
            O => \N__29779\,
            I => \N__29771\
        );

    \I__5397\ : InMux
    port map (
            O => \N__29778\,
            I => \N__29771\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__29771\,
            I => \N__29767\
        );

    \I__5395\ : CascadeMux
    port map (
            O => \N__29770\,
            I => \N__29764\
        );

    \I__5394\ : Span4Mux_v
    port map (
            O => \N__29767\,
            I => \N__29761\
        );

    \I__5393\ : InMux
    port map (
            O => \N__29764\,
            I => \N__29758\
        );

    \I__5392\ : Odrv4
    port map (
            O => \N__29761\,
            I => \current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0\
        );

    \I__5391\ : LocalMux
    port map (
            O => \N__29758\,
            I => \current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0\
        );

    \I__5390\ : InMux
    port map (
            O => \N__29753\,
            I => \current_shift_inst.un4_control_input_cry_22\
        );

    \I__5389\ : InMux
    port map (
            O => \N__29750\,
            I => \current_shift_inst.un4_control_input_cry_23\
        );

    \I__5388\ : InMux
    port map (
            O => \N__29747\,
            I => \bfn_11_17_0_\
        );

    \I__5387\ : InMux
    port map (
            O => \N__29744\,
            I => \current_shift_inst.un4_control_input_cry_25\
        );

    \I__5386\ : InMux
    port map (
            O => \N__29741\,
            I => \current_shift_inst.un4_control_input_cry_26\
        );

    \I__5385\ : InMux
    port map (
            O => \N__29738\,
            I => \N__29733\
        );

    \I__5384\ : InMux
    port map (
            O => \N__29737\,
            I => \N__29728\
        );

    \I__5383\ : InMux
    port map (
            O => \N__29736\,
            I => \N__29728\
        );

    \I__5382\ : LocalMux
    port map (
            O => \N__29733\,
            I => \N__29725\
        );

    \I__5381\ : LocalMux
    port map (
            O => \N__29728\,
            I => \N__29722\
        );

    \I__5380\ : Span4Mux_v
    port map (
            O => \N__29725\,
            I => \N__29718\
        );

    \I__5379\ : Span4Mux_h
    port map (
            O => \N__29722\,
            I => \N__29715\
        );

    \I__5378\ : InMux
    port map (
            O => \N__29721\,
            I => \N__29712\
        );

    \I__5377\ : Odrv4
    port map (
            O => \N__29718\,
            I => \current_shift_inst.un4_control_input_cry_10_c_RNIJLTGZ0\
        );

    \I__5376\ : Odrv4
    port map (
            O => \N__29715\,
            I => \current_shift_inst.un4_control_input_cry_10_c_RNIJLTGZ0\
        );

    \I__5375\ : LocalMux
    port map (
            O => \N__29712\,
            I => \current_shift_inst.un4_control_input_cry_10_c_RNIJLTGZ0\
        );

    \I__5374\ : InMux
    port map (
            O => \N__29705\,
            I => \current_shift_inst.un4_control_input_cry_10\
        );

    \I__5373\ : InMux
    port map (
            O => \N__29702\,
            I => \current_shift_inst.un4_control_input_cry_11\
        );

    \I__5372\ : InMux
    port map (
            O => \N__29699\,
            I => \current_shift_inst.un4_control_input_cry_12\
        );

    \I__5371\ : InMux
    port map (
            O => \N__29696\,
            I => \current_shift_inst.un4_control_input_cry_13\
        );

    \I__5370\ : InMux
    port map (
            O => \N__29693\,
            I => \current_shift_inst.un4_control_input_cry_14\
        );

    \I__5369\ : InMux
    port map (
            O => \N__29690\,
            I => \current_shift_inst.un4_control_input_cry_15\
        );

    \I__5368\ : InMux
    port map (
            O => \N__29687\,
            I => \bfn_11_16_0_\
        );

    \I__5367\ : CascadeMux
    port map (
            O => \N__29684\,
            I => \N__29681\
        );

    \I__5366\ : InMux
    port map (
            O => \N__29681\,
            I => \N__29676\
        );

    \I__5365\ : InMux
    port map (
            O => \N__29680\,
            I => \N__29671\
        );

    \I__5364\ : InMux
    port map (
            O => \N__29679\,
            I => \N__29671\
        );

    \I__5363\ : LocalMux
    port map (
            O => \N__29676\,
            I => \N__29667\
        );

    \I__5362\ : LocalMux
    port map (
            O => \N__29671\,
            I => \N__29664\
        );

    \I__5361\ : CascadeMux
    port map (
            O => \N__29670\,
            I => \N__29661\
        );

    \I__5360\ : Span4Mux_h
    port map (
            O => \N__29667\,
            I => \N__29656\
        );

    \I__5359\ : Span4Mux_v
    port map (
            O => \N__29664\,
            I => \N__29656\
        );

    \I__5358\ : InMux
    port map (
            O => \N__29661\,
            I => \N__29653\
        );

    \I__5357\ : Odrv4
    port map (
            O => \N__29656\,
            I => \current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0\
        );

    \I__5356\ : LocalMux
    port map (
            O => \N__29653\,
            I => \current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0\
        );

    \I__5355\ : InMux
    port map (
            O => \N__29648\,
            I => \current_shift_inst.un4_control_input_cry_17\
        );

    \I__5354\ : InMux
    port map (
            O => \N__29645\,
            I => \N__29642\
        );

    \I__5353\ : LocalMux
    port map (
            O => \N__29642\,
            I => \N__29637\
        );

    \I__5352\ : InMux
    port map (
            O => \N__29641\,
            I => \N__29632\
        );

    \I__5351\ : InMux
    port map (
            O => \N__29640\,
            I => \N__29632\
        );

    \I__5350\ : Span4Mux_v
    port map (
            O => \N__29637\,
            I => \N__29628\
        );

    \I__5349\ : LocalMux
    port map (
            O => \N__29632\,
            I => \N__29625\
        );

    \I__5348\ : InMux
    port map (
            O => \N__29631\,
            I => \N__29622\
        );

    \I__5347\ : Odrv4
    port map (
            O => \N__29628\,
            I => \current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0\
        );

    \I__5346\ : Odrv4
    port map (
            O => \N__29625\,
            I => \current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0\
        );

    \I__5345\ : LocalMux
    port map (
            O => \N__29622\,
            I => \current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0\
        );

    \I__5344\ : CascadeMux
    port map (
            O => \N__29615\,
            I => \N__29611\
        );

    \I__5343\ : InMux
    port map (
            O => \N__29614\,
            I => \N__29608\
        );

    \I__5342\ : InMux
    port map (
            O => \N__29611\,
            I => \N__29605\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__29608\,
            I => \N__29599\
        );

    \I__5340\ : LocalMux
    port map (
            O => \N__29605\,
            I => \N__29599\
        );

    \I__5339\ : CascadeMux
    port map (
            O => \N__29604\,
            I => \N__29596\
        );

    \I__5338\ : Span4Mux_v
    port map (
            O => \N__29599\,
            I => \N__29593\
        );

    \I__5337\ : InMux
    port map (
            O => \N__29596\,
            I => \N__29590\
        );

    \I__5336\ : Odrv4
    port map (
            O => \N__29593\,
            I => \current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0\
        );

    \I__5335\ : LocalMux
    port map (
            O => \N__29590\,
            I => \current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0\
        );

    \I__5334\ : InMux
    port map (
            O => \N__29585\,
            I => \current_shift_inst.un4_control_input_cry_1\
        );

    \I__5333\ : InMux
    port map (
            O => \N__29582\,
            I => \N__29578\
        );

    \I__5332\ : InMux
    port map (
            O => \N__29581\,
            I => \N__29575\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__29578\,
            I => \N__29570\
        );

    \I__5330\ : LocalMux
    port map (
            O => \N__29575\,
            I => \N__29570\
        );

    \I__5329\ : Span4Mux_h
    port map (
            O => \N__29570\,
            I => \N__29566\
        );

    \I__5328\ : InMux
    port map (
            O => \N__29569\,
            I => \N__29563\
        );

    \I__5327\ : Odrv4
    port map (
            O => \N__29566\,
            I => \current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__29563\,
            I => \current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0\
        );

    \I__5325\ : InMux
    port map (
            O => \N__29558\,
            I => \current_shift_inst.un4_control_input_cry_2\
        );

    \I__5324\ : InMux
    port map (
            O => \N__29555\,
            I => \N__29552\
        );

    \I__5323\ : LocalMux
    port map (
            O => \N__29552\,
            I => \N__29549\
        );

    \I__5322\ : Span4Mux_h
    port map (
            O => \N__29549\,
            I => \N__29545\
        );

    \I__5321\ : InMux
    port map (
            O => \N__29548\,
            I => \N__29542\
        );

    \I__5320\ : Odrv4
    port map (
            O => \N__29545\,
            I => \current_shift_inst.un4_control_input_cry_3_c_RNINL4GZ0\
        );

    \I__5319\ : LocalMux
    port map (
            O => \N__29542\,
            I => \current_shift_inst.un4_control_input_cry_3_c_RNINL4GZ0\
        );

    \I__5318\ : InMux
    port map (
            O => \N__29537\,
            I => \current_shift_inst.un4_control_input_cry_3\
        );

    \I__5317\ : CascadeMux
    port map (
            O => \N__29534\,
            I => \N__29531\
        );

    \I__5316\ : InMux
    port map (
            O => \N__29531\,
            I => \N__29526\
        );

    \I__5315\ : InMux
    port map (
            O => \N__29530\,
            I => \N__29523\
        );

    \I__5314\ : InMux
    port map (
            O => \N__29529\,
            I => \N__29520\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__29526\,
            I => \N__29514\
        );

    \I__5312\ : LocalMux
    port map (
            O => \N__29523\,
            I => \N__29514\
        );

    \I__5311\ : LocalMux
    port map (
            O => \N__29520\,
            I => \N__29511\
        );

    \I__5310\ : CascadeMux
    port map (
            O => \N__29519\,
            I => \N__29508\
        );

    \I__5309\ : Span4Mux_h
    port map (
            O => \N__29514\,
            I => \N__29505\
        );

    \I__5308\ : Span4Mux_h
    port map (
            O => \N__29511\,
            I => \N__29502\
        );

    \I__5307\ : InMux
    port map (
            O => \N__29508\,
            I => \N__29499\
        );

    \I__5306\ : Odrv4
    port map (
            O => \N__29505\,
            I => \current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0\
        );

    \I__5305\ : Odrv4
    port map (
            O => \N__29502\,
            I => \current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0\
        );

    \I__5304\ : LocalMux
    port map (
            O => \N__29499\,
            I => \current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0\
        );

    \I__5303\ : InMux
    port map (
            O => \N__29492\,
            I => \current_shift_inst.un4_control_input_cry_4\
        );

    \I__5302\ : InMux
    port map (
            O => \N__29489\,
            I => \N__29484\
        );

    \I__5301\ : InMux
    port map (
            O => \N__29488\,
            I => \N__29479\
        );

    \I__5300\ : InMux
    port map (
            O => \N__29487\,
            I => \N__29479\
        );

    \I__5299\ : LocalMux
    port map (
            O => \N__29484\,
            I => \N__29476\
        );

    \I__5298\ : LocalMux
    port map (
            O => \N__29479\,
            I => \N__29473\
        );

    \I__5297\ : Span4Mux_v
    port map (
            O => \N__29476\,
            I => \N__29469\
        );

    \I__5296\ : Span4Mux_h
    port map (
            O => \N__29473\,
            I => \N__29466\
        );

    \I__5295\ : InMux
    port map (
            O => \N__29472\,
            I => \N__29463\
        );

    \I__5294\ : Odrv4
    port map (
            O => \N__29469\,
            I => \current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0\
        );

    \I__5293\ : Odrv4
    port map (
            O => \N__29466\,
            I => \current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0\
        );

    \I__5292\ : LocalMux
    port map (
            O => \N__29463\,
            I => \current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0\
        );

    \I__5291\ : InMux
    port map (
            O => \N__29456\,
            I => \current_shift_inst.un4_control_input_cry_5\
        );

    \I__5290\ : InMux
    port map (
            O => \N__29453\,
            I => \N__29448\
        );

    \I__5289\ : InMux
    port map (
            O => \N__29452\,
            I => \N__29443\
        );

    \I__5288\ : InMux
    port map (
            O => \N__29451\,
            I => \N__29443\
        );

    \I__5287\ : LocalMux
    port map (
            O => \N__29448\,
            I => \N__29439\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__29443\,
            I => \N__29436\
        );

    \I__5285\ : CascadeMux
    port map (
            O => \N__29442\,
            I => \N__29433\
        );

    \I__5284\ : Span4Mux_h
    port map (
            O => \N__29439\,
            I => \N__29430\
        );

    \I__5283\ : Span4Mux_v
    port map (
            O => \N__29436\,
            I => \N__29427\
        );

    \I__5282\ : InMux
    port map (
            O => \N__29433\,
            I => \N__29424\
        );

    \I__5281\ : Odrv4
    port map (
            O => \N__29430\,
            I => \current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0\
        );

    \I__5280\ : Odrv4
    port map (
            O => \N__29427\,
            I => \current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0\
        );

    \I__5279\ : LocalMux
    port map (
            O => \N__29424\,
            I => \current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0\
        );

    \I__5278\ : InMux
    port map (
            O => \N__29417\,
            I => \current_shift_inst.un4_control_input_cry_6\
        );

    \I__5277\ : CascadeMux
    port map (
            O => \N__29414\,
            I => \N__29411\
        );

    \I__5276\ : InMux
    port map (
            O => \N__29411\,
            I => \N__29408\
        );

    \I__5275\ : LocalMux
    port map (
            O => \N__29408\,
            I => \N__29404\
        );

    \I__5274\ : CascadeMux
    port map (
            O => \N__29407\,
            I => \N__29400\
        );

    \I__5273\ : Span4Mux_h
    port map (
            O => \N__29404\,
            I => \N__29397\
        );

    \I__5272\ : InMux
    port map (
            O => \N__29403\,
            I => \N__29392\
        );

    \I__5271\ : InMux
    port map (
            O => \N__29400\,
            I => \N__29392\
        );

    \I__5270\ : Sp12to4
    port map (
            O => \N__29397\,
            I => \N__29388\
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__29392\,
            I => \N__29385\
        );

    \I__5268\ : CascadeMux
    port map (
            O => \N__29391\,
            I => \N__29382\
        );

    \I__5267\ : Span12Mux_v
    port map (
            O => \N__29388\,
            I => \N__29379\
        );

    \I__5266\ : Span4Mux_v
    port map (
            O => \N__29385\,
            I => \N__29376\
        );

    \I__5265\ : InMux
    port map (
            O => \N__29382\,
            I => \N__29373\
        );

    \I__5264\ : Odrv12
    port map (
            O => \N__29379\,
            I => \current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0\
        );

    \I__5263\ : Odrv4
    port map (
            O => \N__29376\,
            I => \current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0\
        );

    \I__5262\ : LocalMux
    port map (
            O => \N__29373\,
            I => \current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0\
        );

    \I__5261\ : InMux
    port map (
            O => \N__29366\,
            I => \current_shift_inst.un4_control_input_cry_7\
        );

    \I__5260\ : InMux
    port map (
            O => \N__29363\,
            I => \bfn_11_15_0_\
        );

    \I__5259\ : InMux
    port map (
            O => \N__29360\,
            I => \current_shift_inst.un4_control_input_cry_9\
        );

    \I__5258\ : CascadeMux
    port map (
            O => \N__29357\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6_cascade_\
        );

    \I__5257\ : CascadeMux
    port map (
            O => \N__29354\,
            I => \N__29351\
        );

    \I__5256\ : InMux
    port map (
            O => \N__29351\,
            I => \N__29348\
        );

    \I__5255\ : LocalMux
    port map (
            O => \N__29348\,
            I => \N__29345\
        );

    \I__5254\ : Odrv4
    port map (
            O => \N__29345\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\
        );

    \I__5253\ : CascadeMux
    port map (
            O => \N__29342\,
            I => \N__29339\
        );

    \I__5252\ : InMux
    port map (
            O => \N__29339\,
            I => \N__29336\
        );

    \I__5251\ : LocalMux
    port map (
            O => \N__29336\,
            I => \N__29333\
        );

    \I__5250\ : Span4Mux_h
    port map (
            O => \N__29333\,
            I => \N__29330\
        );

    \I__5249\ : Odrv4
    port map (
            O => \N__29330\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\
        );

    \I__5248\ : CascadeMux
    port map (
            O => \N__29327\,
            I => \N__29322\
        );

    \I__5247\ : InMux
    port map (
            O => \N__29326\,
            I => \N__29319\
        );

    \I__5246\ : InMux
    port map (
            O => \N__29325\,
            I => \N__29316\
        );

    \I__5245\ : InMux
    port map (
            O => \N__29322\,
            I => \N__29313\
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__29319\,
            I => \current_shift_inst.elapsed_time_ns_1_fast_31\
        );

    \I__5243\ : LocalMux
    port map (
            O => \N__29316\,
            I => \current_shift_inst.elapsed_time_ns_1_fast_31\
        );

    \I__5242\ : LocalMux
    port map (
            O => \N__29313\,
            I => \current_shift_inst.elapsed_time_ns_1_fast_31\
        );

    \I__5241\ : CascadeMux
    port map (
            O => \N__29306\,
            I => \N__29303\
        );

    \I__5240\ : InMux
    port map (
            O => \N__29303\,
            I => \N__29300\
        );

    \I__5239\ : LocalMux
    port map (
            O => \N__29300\,
            I => \N__29297\
        );

    \I__5238\ : Span4Mux_v
    port map (
            O => \N__29297\,
            I => \N__29294\
        );

    \I__5237\ : Span4Mux_h
    port map (
            O => \N__29294\,
            I => \N__29290\
        );

    \I__5236\ : InMux
    port map (
            O => \N__29293\,
            I => \N__29287\
        );

    \I__5235\ : Odrv4
    port map (
            O => \N__29290\,
            I => \current_shift_inst.un38_control_input_0\
        );

    \I__5234\ : LocalMux
    port map (
            O => \N__29287\,
            I => \current_shift_inst.un38_control_input_0\
        );

    \I__5233\ : InMux
    port map (
            O => \N__29282\,
            I => \N__29279\
        );

    \I__5232\ : LocalMux
    port map (
            O => \N__29279\,
            I => \N__29275\
        );

    \I__5231\ : InMux
    port map (
            O => \N__29278\,
            I => \N__29272\
        );

    \I__5230\ : Span4Mux_h
    port map (
            O => \N__29275\,
            I => \N__29269\
        );

    \I__5229\ : LocalMux
    port map (
            O => \N__29272\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__5228\ : Odrv4
    port map (
            O => \N__29269\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__5227\ : InMux
    port map (
            O => \N__29264\,
            I => \N__29261\
        );

    \I__5226\ : LocalMux
    port map (
            O => \N__29261\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13\
        );

    \I__5225\ : InMux
    port map (
            O => \N__29258\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\
        );

    \I__5224\ : InMux
    port map (
            O => \N__29255\,
            I => \N__29251\
        );

    \I__5223\ : InMux
    port map (
            O => \N__29254\,
            I => \N__29248\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__29251\,
            I => \N__29245\
        );

    \I__5221\ : LocalMux
    port map (
            O => \N__29248\,
            I => \N__29242\
        );

    \I__5220\ : Odrv12
    port map (
            O => \N__29245\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__5219\ : Odrv4
    port map (
            O => \N__29242\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__5218\ : InMux
    port map (
            O => \N__29237\,
            I => \N__29234\
        );

    \I__5217\ : LocalMux
    port map (
            O => \N__29234\,
            I => \N__29231\
        );

    \I__5216\ : Odrv4
    port map (
            O => \N__29231\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14\
        );

    \I__5215\ : InMux
    port map (
            O => \N__29228\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\
        );

    \I__5214\ : InMux
    port map (
            O => \N__29225\,
            I => \N__29222\
        );

    \I__5213\ : LocalMux
    port map (
            O => \N__29222\,
            I => \N__29218\
        );

    \I__5212\ : InMux
    port map (
            O => \N__29221\,
            I => \N__29215\
        );

    \I__5211\ : Span4Mux_v
    port map (
            O => \N__29218\,
            I => \N__29212\
        );

    \I__5210\ : LocalMux
    port map (
            O => \N__29215\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__5209\ : Odrv4
    port map (
            O => \N__29212\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__5208\ : InMux
    port map (
            O => \N__29207\,
            I => \N__29204\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__29204\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15\
        );

    \I__5206\ : InMux
    port map (
            O => \N__29201\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\
        );

    \I__5205\ : InMux
    port map (
            O => \N__29198\,
            I => \N__29195\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__29195\,
            I => \N__29191\
        );

    \I__5203\ : InMux
    port map (
            O => \N__29194\,
            I => \N__29188\
        );

    \I__5202\ : Span4Mux_h
    port map (
            O => \N__29191\,
            I => \N__29185\
        );

    \I__5201\ : LocalMux
    port map (
            O => \N__29188\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__5200\ : Odrv4
    port map (
            O => \N__29185\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__5199\ : InMux
    port map (
            O => \N__29180\,
            I => \N__29177\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__29177\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16\
        );

    \I__5197\ : InMux
    port map (
            O => \N__29174\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\
        );

    \I__5196\ : InMux
    port map (
            O => \N__29171\,
            I => \N__29168\
        );

    \I__5195\ : LocalMux
    port map (
            O => \N__29168\,
            I => \N__29164\
        );

    \I__5194\ : InMux
    port map (
            O => \N__29167\,
            I => \N__29161\
        );

    \I__5193\ : Span4Mux_h
    port map (
            O => \N__29164\,
            I => \N__29158\
        );

    \I__5192\ : LocalMux
    port map (
            O => \N__29161\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__5191\ : Odrv4
    port map (
            O => \N__29158\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__5190\ : InMux
    port map (
            O => \N__29153\,
            I => \N__29150\
        );

    \I__5189\ : LocalMux
    port map (
            O => \N__29150\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17\
        );

    \I__5188\ : InMux
    port map (
            O => \N__29147\,
            I => \bfn_11_10_0_\
        );

    \I__5187\ : InMux
    port map (
            O => \N__29144\,
            I => \N__29141\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__29141\,
            I => \N__29137\
        );

    \I__5185\ : InMux
    port map (
            O => \N__29140\,
            I => \N__29134\
        );

    \I__5184\ : Span4Mux_v
    port map (
            O => \N__29137\,
            I => \N__29131\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__29134\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__5182\ : Odrv4
    port map (
            O => \N__29131\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__5181\ : InMux
    port map (
            O => \N__29126\,
            I => \N__29123\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__29123\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18\
        );

    \I__5179\ : InMux
    port map (
            O => \N__29120\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\
        );

    \I__5178\ : InMux
    port map (
            O => \N__29117\,
            I => \N__29114\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__29114\,
            I => \N__29110\
        );

    \I__5176\ : InMux
    port map (
            O => \N__29113\,
            I => \N__29107\
        );

    \I__5175\ : Span4Mux_h
    port map (
            O => \N__29110\,
            I => \N__29104\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__29107\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__5173\ : Odrv4
    port map (
            O => \N__29104\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__5172\ : InMux
    port map (
            O => \N__29099\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17\
        );

    \I__5171\ : InMux
    port map (
            O => \N__29096\,
            I => \N__29093\
        );

    \I__5170\ : LocalMux
    port map (
            O => \N__29093\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19\
        );

    \I__5169\ : InMux
    port map (
            O => \N__29090\,
            I => \N__29087\
        );

    \I__5168\ : LocalMux
    port map (
            O => \N__29087\,
            I => \N__29084\
        );

    \I__5167\ : Odrv12
    port map (
            O => \N__29084\,
            I => \il_min_comp1_D1\
        );

    \I__5166\ : InMux
    port map (
            O => \N__29081\,
            I => \N__29078\
        );

    \I__5165\ : LocalMux
    port map (
            O => \N__29078\,
            I => \N__29075\
        );

    \I__5164\ : Span4Mux_v
    port map (
            O => \N__29075\,
            I => \N__29071\
        );

    \I__5163\ : InMux
    port map (
            O => \N__29074\,
            I => \N__29068\
        );

    \I__5162\ : Odrv4
    port map (
            O => \N__29071\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__5161\ : LocalMux
    port map (
            O => \N__29068\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__5160\ : InMux
    port map (
            O => \N__29063\,
            I => \N__29060\
        );

    \I__5159\ : LocalMux
    port map (
            O => \N__29060\,
            I => \N__29057\
        );

    \I__5158\ : Span4Mux_h
    port map (
            O => \N__29057\,
            I => \N__29054\
        );

    \I__5157\ : Odrv4
    port map (
            O => \N__29054\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5\
        );

    \I__5156\ : InMux
    port map (
            O => \N__29051\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\
        );

    \I__5155\ : InMux
    port map (
            O => \N__29048\,
            I => \N__29045\
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__29045\,
            I => \N__29042\
        );

    \I__5153\ : Span4Mux_h
    port map (
            O => \N__29042\,
            I => \N__29038\
        );

    \I__5152\ : InMux
    port map (
            O => \N__29041\,
            I => \N__29035\
        );

    \I__5151\ : Odrv4
    port map (
            O => \N__29038\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__29035\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__5149\ : InMux
    port map (
            O => \N__29030\,
            I => \N__29027\
        );

    \I__5148\ : LocalMux
    port map (
            O => \N__29027\,
            I => \N__29024\
        );

    \I__5147\ : Span4Mux_h
    port map (
            O => \N__29024\,
            I => \N__29021\
        );

    \I__5146\ : Odrv4
    port map (
            O => \N__29021\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6\
        );

    \I__5145\ : InMux
    port map (
            O => \N__29018\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\
        );

    \I__5144\ : InMux
    port map (
            O => \N__29015\,
            I => \N__29012\
        );

    \I__5143\ : LocalMux
    port map (
            O => \N__29012\,
            I => \N__29009\
        );

    \I__5142\ : Span4Mux_h
    port map (
            O => \N__29009\,
            I => \N__29005\
        );

    \I__5141\ : InMux
    port map (
            O => \N__29008\,
            I => \N__29002\
        );

    \I__5140\ : Odrv4
    port map (
            O => \N__29005\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__5139\ : LocalMux
    port map (
            O => \N__29002\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__5138\ : InMux
    port map (
            O => \N__28997\,
            I => \N__28994\
        );

    \I__5137\ : LocalMux
    port map (
            O => \N__28994\,
            I => \N__28991\
        );

    \I__5136\ : Span4Mux_h
    port map (
            O => \N__28991\,
            I => \N__28988\
        );

    \I__5135\ : Odrv4
    port map (
            O => \N__28988\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7\
        );

    \I__5134\ : InMux
    port map (
            O => \N__28985\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\
        );

    \I__5133\ : InMux
    port map (
            O => \N__28982\,
            I => \N__28979\
        );

    \I__5132\ : LocalMux
    port map (
            O => \N__28979\,
            I => \N__28975\
        );

    \I__5131\ : InMux
    port map (
            O => \N__28978\,
            I => \N__28972\
        );

    \I__5130\ : Span4Mux_h
    port map (
            O => \N__28975\,
            I => \N__28967\
        );

    \I__5129\ : LocalMux
    port map (
            O => \N__28972\,
            I => \N__28967\
        );

    \I__5128\ : Odrv4
    port map (
            O => \N__28967\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__5127\ : InMux
    port map (
            O => \N__28964\,
            I => \N__28961\
        );

    \I__5126\ : LocalMux
    port map (
            O => \N__28961\,
            I => \N__28958\
        );

    \I__5125\ : Span4Mux_h
    port map (
            O => \N__28958\,
            I => \N__28955\
        );

    \I__5124\ : Odrv4
    port map (
            O => \N__28955\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8\
        );

    \I__5123\ : InMux
    port map (
            O => \N__28952\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\
        );

    \I__5122\ : InMux
    port map (
            O => \N__28949\,
            I => \bfn_11_9_0_\
        );

    \I__5121\ : InMux
    port map (
            O => \N__28946\,
            I => \N__28942\
        );

    \I__5120\ : InMux
    port map (
            O => \N__28945\,
            I => \N__28939\
        );

    \I__5119\ : LocalMux
    port map (
            O => \N__28942\,
            I => \N__28936\
        );

    \I__5118\ : LocalMux
    port map (
            O => \N__28939\,
            I => \N__28933\
        );

    \I__5117\ : Odrv4
    port map (
            O => \N__28936\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__5116\ : Odrv4
    port map (
            O => \N__28933\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__5115\ : InMux
    port map (
            O => \N__28928\,
            I => \N__28925\
        );

    \I__5114\ : LocalMux
    port map (
            O => \N__28925\,
            I => \N__28922\
        );

    \I__5113\ : Odrv12
    port map (
            O => \N__28922\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10\
        );

    \I__5112\ : InMux
    port map (
            O => \N__28919\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\
        );

    \I__5111\ : InMux
    port map (
            O => \N__28916\,
            I => \N__28912\
        );

    \I__5110\ : CascadeMux
    port map (
            O => \N__28915\,
            I => \N__28909\
        );

    \I__5109\ : LocalMux
    port map (
            O => \N__28912\,
            I => \N__28906\
        );

    \I__5108\ : InMux
    port map (
            O => \N__28909\,
            I => \N__28903\
        );

    \I__5107\ : Span4Mux_v
    port map (
            O => \N__28906\,
            I => \N__28900\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__28903\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__5105\ : Odrv4
    port map (
            O => \N__28900\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__5104\ : InMux
    port map (
            O => \N__28895\,
            I => \N__28892\
        );

    \I__5103\ : LocalMux
    port map (
            O => \N__28892\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11\
        );

    \I__5102\ : InMux
    port map (
            O => \N__28889\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\
        );

    \I__5101\ : InMux
    port map (
            O => \N__28886\,
            I => \N__28882\
        );

    \I__5100\ : CascadeMux
    port map (
            O => \N__28885\,
            I => \N__28879\
        );

    \I__5099\ : LocalMux
    port map (
            O => \N__28882\,
            I => \N__28876\
        );

    \I__5098\ : InMux
    port map (
            O => \N__28879\,
            I => \N__28873\
        );

    \I__5097\ : Span4Mux_h
    port map (
            O => \N__28876\,
            I => \N__28870\
        );

    \I__5096\ : LocalMux
    port map (
            O => \N__28873\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__5095\ : Odrv4
    port map (
            O => \N__28870\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__5094\ : InMux
    port map (
            O => \N__28865\,
            I => \N__28862\
        );

    \I__5093\ : LocalMux
    port map (
            O => \N__28862\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12\
        );

    \I__5092\ : InMux
    port map (
            O => \N__28859\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\
        );

    \I__5091\ : InMux
    port map (
            O => \N__28856\,
            I => \N__28824\
        );

    \I__5090\ : InMux
    port map (
            O => \N__28855\,
            I => \N__28810\
        );

    \I__5089\ : InMux
    port map (
            O => \N__28854\,
            I => \N__28810\
        );

    \I__5088\ : InMux
    port map (
            O => \N__28853\,
            I => \N__28810\
        );

    \I__5087\ : InMux
    port map (
            O => \N__28852\,
            I => \N__28801\
        );

    \I__5086\ : InMux
    port map (
            O => \N__28851\,
            I => \N__28801\
        );

    \I__5085\ : InMux
    port map (
            O => \N__28850\,
            I => \N__28801\
        );

    \I__5084\ : InMux
    port map (
            O => \N__28849\,
            I => \N__28801\
        );

    \I__5083\ : CascadeMux
    port map (
            O => \N__28848\,
            I => \N__28797\
        );

    \I__5082\ : CascadeMux
    port map (
            O => \N__28847\,
            I => \N__28793\
        );

    \I__5081\ : CascadeMux
    port map (
            O => \N__28846\,
            I => \N__28789\
        );

    \I__5080\ : CascadeMux
    port map (
            O => \N__28845\,
            I => \N__28786\
        );

    \I__5079\ : CascadeMux
    port map (
            O => \N__28844\,
            I => \N__28783\
        );

    \I__5078\ : CascadeMux
    port map (
            O => \N__28843\,
            I => \N__28780\
        );

    \I__5077\ : CascadeMux
    port map (
            O => \N__28842\,
            I => \N__28777\
        );

    \I__5076\ : CascadeMux
    port map (
            O => \N__28841\,
            I => \N__28774\
        );

    \I__5075\ : CascadeMux
    port map (
            O => \N__28840\,
            I => \N__28771\
        );

    \I__5074\ : CascadeMux
    port map (
            O => \N__28839\,
            I => \N__28768\
        );

    \I__5073\ : CascadeMux
    port map (
            O => \N__28838\,
            I => \N__28765\
        );

    \I__5072\ : CascadeMux
    port map (
            O => \N__28837\,
            I => \N__28762\
        );

    \I__5071\ : CascadeMux
    port map (
            O => \N__28836\,
            I => \N__28759\
        );

    \I__5070\ : CascadeMux
    port map (
            O => \N__28835\,
            I => \N__28756\
        );

    \I__5069\ : CascadeMux
    port map (
            O => \N__28834\,
            I => \N__28753\
        );

    \I__5068\ : CascadeMux
    port map (
            O => \N__28833\,
            I => \N__28750\
        );

    \I__5067\ : CascadeMux
    port map (
            O => \N__28832\,
            I => \N__28747\
        );

    \I__5066\ : CascadeMux
    port map (
            O => \N__28831\,
            I => \N__28744\
        );

    \I__5065\ : CascadeMux
    port map (
            O => \N__28830\,
            I => \N__28741\
        );

    \I__5064\ : CascadeMux
    port map (
            O => \N__28829\,
            I => \N__28738\
        );

    \I__5063\ : CascadeMux
    port map (
            O => \N__28828\,
            I => \N__28735\
        );

    \I__5062\ : CascadeMux
    port map (
            O => \N__28827\,
            I => \N__28732\
        );

    \I__5061\ : LocalMux
    port map (
            O => \N__28824\,
            I => \N__28728\
        );

    \I__5060\ : InMux
    port map (
            O => \N__28823\,
            I => \N__28721\
        );

    \I__5059\ : InMux
    port map (
            O => \N__28822\,
            I => \N__28721\
        );

    \I__5058\ : InMux
    port map (
            O => \N__28821\,
            I => \N__28721\
        );

    \I__5057\ : InMux
    port map (
            O => \N__28820\,
            I => \N__28712\
        );

    \I__5056\ : InMux
    port map (
            O => \N__28819\,
            I => \N__28712\
        );

    \I__5055\ : InMux
    port map (
            O => \N__28818\,
            I => \N__28712\
        );

    \I__5054\ : InMux
    port map (
            O => \N__28817\,
            I => \N__28712\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__28810\,
            I => \N__28707\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__28801\,
            I => \N__28707\
        );

    \I__5051\ : InMux
    port map (
            O => \N__28800\,
            I => \N__28700\
        );

    \I__5050\ : InMux
    port map (
            O => \N__28797\,
            I => \N__28700\
        );

    \I__5049\ : InMux
    port map (
            O => \N__28796\,
            I => \N__28700\
        );

    \I__5048\ : InMux
    port map (
            O => \N__28793\,
            I => \N__28682\
        );

    \I__5047\ : InMux
    port map (
            O => \N__28792\,
            I => \N__28682\
        );

    \I__5046\ : InMux
    port map (
            O => \N__28789\,
            I => \N__28682\
        );

    \I__5045\ : InMux
    port map (
            O => \N__28786\,
            I => \N__28682\
        );

    \I__5044\ : InMux
    port map (
            O => \N__28783\,
            I => \N__28682\
        );

    \I__5043\ : InMux
    port map (
            O => \N__28780\,
            I => \N__28675\
        );

    \I__5042\ : InMux
    port map (
            O => \N__28777\,
            I => \N__28675\
        );

    \I__5041\ : InMux
    port map (
            O => \N__28774\,
            I => \N__28675\
        );

    \I__5040\ : InMux
    port map (
            O => \N__28771\,
            I => \N__28666\
        );

    \I__5039\ : InMux
    port map (
            O => \N__28768\,
            I => \N__28666\
        );

    \I__5038\ : InMux
    port map (
            O => \N__28765\,
            I => \N__28666\
        );

    \I__5037\ : InMux
    port map (
            O => \N__28762\,
            I => \N__28666\
        );

    \I__5036\ : InMux
    port map (
            O => \N__28759\,
            I => \N__28657\
        );

    \I__5035\ : InMux
    port map (
            O => \N__28756\,
            I => \N__28657\
        );

    \I__5034\ : InMux
    port map (
            O => \N__28753\,
            I => \N__28657\
        );

    \I__5033\ : InMux
    port map (
            O => \N__28750\,
            I => \N__28657\
        );

    \I__5032\ : InMux
    port map (
            O => \N__28747\,
            I => \N__28649\
        );

    \I__5031\ : InMux
    port map (
            O => \N__28744\,
            I => \N__28649\
        );

    \I__5030\ : InMux
    port map (
            O => \N__28741\,
            I => \N__28649\
        );

    \I__5029\ : InMux
    port map (
            O => \N__28738\,
            I => \N__28642\
        );

    \I__5028\ : InMux
    port map (
            O => \N__28735\,
            I => \N__28642\
        );

    \I__5027\ : InMux
    port map (
            O => \N__28732\,
            I => \N__28642\
        );

    \I__5026\ : InMux
    port map (
            O => \N__28731\,
            I => \N__28639\
        );

    \I__5025\ : Span4Mux_v
    port map (
            O => \N__28728\,
            I => \N__28632\
        );

    \I__5024\ : LocalMux
    port map (
            O => \N__28721\,
            I => \N__28632\
        );

    \I__5023\ : LocalMux
    port map (
            O => \N__28712\,
            I => \N__28632\
        );

    \I__5022\ : Span4Mux_s2_h
    port map (
            O => \N__28707\,
            I => \N__28627\
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__28700\,
            I => \N__28627\
        );

    \I__5020\ : CascadeMux
    port map (
            O => \N__28699\,
            I => \N__28624\
        );

    \I__5019\ : CascadeMux
    port map (
            O => \N__28698\,
            I => \N__28621\
        );

    \I__5018\ : CascadeMux
    port map (
            O => \N__28697\,
            I => \N__28618\
        );

    \I__5017\ : CascadeMux
    port map (
            O => \N__28696\,
            I => \N__28615\
        );

    \I__5016\ : CascadeMux
    port map (
            O => \N__28695\,
            I => \N__28612\
        );

    \I__5015\ : CascadeMux
    port map (
            O => \N__28694\,
            I => \N__28609\
        );

    \I__5014\ : CascadeMux
    port map (
            O => \N__28693\,
            I => \N__28606\
        );

    \I__5013\ : LocalMux
    port map (
            O => \N__28682\,
            I => \N__28603\
        );

    \I__5012\ : LocalMux
    port map (
            O => \N__28675\,
            I => \N__28600\
        );

    \I__5011\ : LocalMux
    port map (
            O => \N__28666\,
            I => \N__28595\
        );

    \I__5010\ : LocalMux
    port map (
            O => \N__28657\,
            I => \N__28595\
        );

    \I__5009\ : InMux
    port map (
            O => \N__28656\,
            I => \N__28592\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__28649\,
            I => \N__28587\
        );

    \I__5007\ : LocalMux
    port map (
            O => \N__28642\,
            I => \N__28587\
        );

    \I__5006\ : LocalMux
    port map (
            O => \N__28639\,
            I => \N__28582\
        );

    \I__5005\ : Span4Mux_v
    port map (
            O => \N__28632\,
            I => \N__28582\
        );

    \I__5004\ : Sp12to4
    port map (
            O => \N__28627\,
            I => \N__28579\
        );

    \I__5003\ : InMux
    port map (
            O => \N__28624\,
            I => \N__28572\
        );

    \I__5002\ : InMux
    port map (
            O => \N__28621\,
            I => \N__28572\
        );

    \I__5001\ : InMux
    port map (
            O => \N__28618\,
            I => \N__28572\
        );

    \I__5000\ : InMux
    port map (
            O => \N__28615\,
            I => \N__28563\
        );

    \I__4999\ : InMux
    port map (
            O => \N__28612\,
            I => \N__28563\
        );

    \I__4998\ : InMux
    port map (
            O => \N__28609\,
            I => \N__28563\
        );

    \I__4997\ : InMux
    port map (
            O => \N__28606\,
            I => \N__28563\
        );

    \I__4996\ : Span4Mux_v
    port map (
            O => \N__28603\,
            I => \N__28558\
        );

    \I__4995\ : Span4Mux_v
    port map (
            O => \N__28600\,
            I => \N__28558\
        );

    \I__4994\ : Span4Mux_v
    port map (
            O => \N__28595\,
            I => \N__28555\
        );

    \I__4993\ : LocalMux
    port map (
            O => \N__28592\,
            I => \N__28552\
        );

    \I__4992\ : Span4Mux_h
    port map (
            O => \N__28587\,
            I => \N__28549\
        );

    \I__4991\ : Span4Mux_h
    port map (
            O => \N__28582\,
            I => \N__28544\
        );

    \I__4990\ : Span12Mux_v
    port map (
            O => \N__28579\,
            I => \N__28537\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__28572\,
            I => \N__28537\
        );

    \I__4988\ : LocalMux
    port map (
            O => \N__28563\,
            I => \N__28537\
        );

    \I__4987\ : Span4Mux_v
    port map (
            O => \N__28558\,
            I => \N__28532\
        );

    \I__4986\ : Span4Mux_v
    port map (
            O => \N__28555\,
            I => \N__28532\
        );

    \I__4985\ : Span4Mux_v
    port map (
            O => \N__28552\,
            I => \N__28529\
        );

    \I__4984\ : Span4Mux_v
    port map (
            O => \N__28549\,
            I => \N__28525\
        );

    \I__4983\ : InMux
    port map (
            O => \N__28548\,
            I => \N__28522\
        );

    \I__4982\ : InMux
    port map (
            O => \N__28547\,
            I => \N__28519\
        );

    \I__4981\ : Sp12to4
    port map (
            O => \N__28544\,
            I => \N__28516\
        );

    \I__4980\ : Span12Mux_h
    port map (
            O => \N__28537\,
            I => \N__28513\
        );

    \I__4979\ : Span4Mux_v
    port map (
            O => \N__28532\,
            I => \N__28510\
        );

    \I__4978\ : Sp12to4
    port map (
            O => \N__28529\,
            I => \N__28507\
        );

    \I__4977\ : InMux
    port map (
            O => \N__28528\,
            I => \N__28504\
        );

    \I__4976\ : Span4Mux_v
    port map (
            O => \N__28525\,
            I => \N__28501\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__28522\,
            I => \N__28496\
        );

    \I__4974\ : LocalMux
    port map (
            O => \N__28519\,
            I => \N__28496\
        );

    \I__4973\ : Span12Mux_v
    port map (
            O => \N__28516\,
            I => \N__28493\
        );

    \I__4972\ : Span12Mux_v
    port map (
            O => \N__28513\,
            I => \N__28486\
        );

    \I__4971\ : Sp12to4
    port map (
            O => \N__28510\,
            I => \N__28486\
        );

    \I__4970\ : Span12Mux_s11_h
    port map (
            O => \N__28507\,
            I => \N__28486\
        );

    \I__4969\ : LocalMux
    port map (
            O => \N__28504\,
            I => \N__28483\
        );

    \I__4968\ : Span4Mux_h
    port map (
            O => \N__28501\,
            I => \N__28478\
        );

    \I__4967\ : Span4Mux_h
    port map (
            O => \N__28496\,
            I => \N__28478\
        );

    \I__4966\ : Odrv12
    port map (
            O => \N__28493\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4965\ : Odrv12
    port map (
            O => \N__28486\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4964\ : Odrv12
    port map (
            O => \N__28483\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4963\ : Odrv4
    port map (
            O => \N__28478\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4962\ : CascadeMux
    port map (
            O => \N__28469\,
            I => \N__28466\
        );

    \I__4961\ : InMux
    port map (
            O => \N__28466\,
            I => \N__28463\
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__28463\,
            I => \N__28460\
        );

    \I__4959\ : Span4Mux_h
    port map (
            O => \N__28460\,
            I => \N__28457\
        );

    \I__4958\ : Odrv4
    port map (
            O => \N__28457\,
            I => \current_shift_inst.z_5_30\
        );

    \I__4957\ : InMux
    port map (
            O => \N__28454\,
            I => \current_shift_inst.z_5_cry_29\
        );

    \I__4956\ : InMux
    port map (
            O => \N__28451\,
            I => \current_shift_inst.z_5_cry_30\
        );

    \I__4955\ : InMux
    port map (
            O => \N__28448\,
            I => \N__28445\
        );

    \I__4954\ : LocalMux
    port map (
            O => \N__28445\,
            I => \N__28442\
        );

    \I__4953\ : Span4Mux_v
    port map (
            O => \N__28442\,
            I => \N__28439\
        );

    \I__4952\ : Odrv4
    port map (
            O => \N__28439\,
            I => \current_shift_inst.z_5_cry_30_THRU_CO\
        );

    \I__4951\ : IoInMux
    port map (
            O => \N__28436\,
            I => \N__28433\
        );

    \I__4950\ : LocalMux
    port map (
            O => \N__28433\,
            I => \N__28430\
        );

    \I__4949\ : IoSpan4Mux
    port map (
            O => \N__28430\,
            I => \N__28427\
        );

    \I__4948\ : Span4Mux_s2_v
    port map (
            O => \N__28427\,
            I => \N__28424\
        );

    \I__4947\ : Odrv4
    port map (
            O => \N__28424\,
            I => s4_phy_c
        );

    \I__4946\ : InMux
    port map (
            O => \N__28421\,
            I => \N__28418\
        );

    \I__4945\ : LocalMux
    port map (
            O => \N__28418\,
            I => \N__28415\
        );

    \I__4944\ : Span4Mux_h
    port map (
            O => \N__28415\,
            I => \N__28412\
        );

    \I__4943\ : Span4Mux_v
    port map (
            O => \N__28412\,
            I => \N__28409\
        );

    \I__4942\ : Odrv4
    port map (
            O => \N__28409\,
            I => il_min_comp1_c
        );

    \I__4941\ : InMux
    port map (
            O => \N__28406\,
            I => \N__28403\
        );

    \I__4940\ : LocalMux
    port map (
            O => \N__28403\,
            I => \N__28400\
        );

    \I__4939\ : Span4Mux_h
    port map (
            O => \N__28400\,
            I => \N__28397\
        );

    \I__4938\ : Span4Mux_v
    port map (
            O => \N__28397\,
            I => \N__28394\
        );

    \I__4937\ : Odrv4
    port map (
            O => \N__28394\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0\
        );

    \I__4936\ : CascadeMux
    port map (
            O => \N__28391\,
            I => \N__28388\
        );

    \I__4935\ : InMux
    port map (
            O => \N__28388\,
            I => \N__28384\
        );

    \I__4934\ : InMux
    port map (
            O => \N__28387\,
            I => \N__28381\
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__28384\,
            I => \N__28378\
        );

    \I__4932\ : LocalMux
    port map (
            O => \N__28381\,
            I => \N__28374\
        );

    \I__4931\ : Span4Mux_h
    port map (
            O => \N__28378\,
            I => \N__28371\
        );

    \I__4930\ : InMux
    port map (
            O => \N__28377\,
            I => \N__28368\
        );

    \I__4929\ : Odrv4
    port map (
            O => \N__28374\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__4928\ : Odrv4
    port map (
            O => \N__28371\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__4927\ : LocalMux
    port map (
            O => \N__28368\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__4926\ : InMux
    port map (
            O => \N__28361\,
            I => \N__28358\
        );

    \I__4925\ : LocalMux
    port map (
            O => \N__28358\,
            I => \N__28355\
        );

    \I__4924\ : Span4Mux_h
    port map (
            O => \N__28355\,
            I => \N__28351\
        );

    \I__4923\ : InMux
    port map (
            O => \N__28354\,
            I => \N__28348\
        );

    \I__4922\ : Odrv4
    port map (
            O => \N__28351\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__4921\ : LocalMux
    port map (
            O => \N__28348\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__4920\ : InMux
    port map (
            O => \N__28343\,
            I => \N__28340\
        );

    \I__4919\ : LocalMux
    port map (
            O => \N__28340\,
            I => \N__28337\
        );

    \I__4918\ : Span4Mux_h
    port map (
            O => \N__28337\,
            I => \N__28334\
        );

    \I__4917\ : Odrv4
    port map (
            O => \N__28334\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2\
        );

    \I__4916\ : InMux
    port map (
            O => \N__28331\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\
        );

    \I__4915\ : InMux
    port map (
            O => \N__28328\,
            I => \N__28325\
        );

    \I__4914\ : LocalMux
    port map (
            O => \N__28325\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0\
        );

    \I__4913\ : CascadeMux
    port map (
            O => \N__28322\,
            I => \N__28319\
        );

    \I__4912\ : InMux
    port map (
            O => \N__28319\,
            I => \N__28316\
        );

    \I__4911\ : LocalMux
    port map (
            O => \N__28316\,
            I => \N__28313\
        );

    \I__4910\ : Span4Mux_h
    port map (
            O => \N__28313\,
            I => \N__28309\
        );

    \I__4909\ : InMux
    port map (
            O => \N__28312\,
            I => \N__28306\
        );

    \I__4908\ : Odrv4
    port map (
            O => \N__28309\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__4907\ : LocalMux
    port map (
            O => \N__28306\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__4906\ : InMux
    port map (
            O => \N__28301\,
            I => \N__28298\
        );

    \I__4905\ : LocalMux
    port map (
            O => \N__28298\,
            I => \N__28295\
        );

    \I__4904\ : Span4Mux_v
    port map (
            O => \N__28295\,
            I => \N__28292\
        );

    \I__4903\ : Odrv4
    port map (
            O => \N__28292\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3\
        );

    \I__4902\ : InMux
    port map (
            O => \N__28289\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\
        );

    \I__4901\ : InMux
    port map (
            O => \N__28286\,
            I => \N__28283\
        );

    \I__4900\ : LocalMux
    port map (
            O => \N__28283\,
            I => \N__28280\
        );

    \I__4899\ : Span4Mux_v
    port map (
            O => \N__28280\,
            I => \N__28276\
        );

    \I__4898\ : InMux
    port map (
            O => \N__28279\,
            I => \N__28273\
        );

    \I__4897\ : Odrv4
    port map (
            O => \N__28276\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__4896\ : LocalMux
    port map (
            O => \N__28273\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__4895\ : InMux
    port map (
            O => \N__28268\,
            I => \N__28265\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__28265\,
            I => \N__28262\
        );

    \I__4893\ : Span4Mux_v
    port map (
            O => \N__28262\,
            I => \N__28259\
        );

    \I__4892\ : Odrv4
    port map (
            O => \N__28259\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4\
        );

    \I__4891\ : InMux
    port map (
            O => \N__28256\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\
        );

    \I__4890\ : InMux
    port map (
            O => \N__28253\,
            I => \current_shift_inst.z_5_cry_20\
        );

    \I__4889\ : InMux
    port map (
            O => \N__28250\,
            I => \N__28240\
        );

    \I__4888\ : InMux
    port map (
            O => \N__28249\,
            I => \N__28240\
        );

    \I__4887\ : InMux
    port map (
            O => \N__28248\,
            I => \N__28240\
        );

    \I__4886\ : InMux
    port map (
            O => \N__28247\,
            I => \N__28237\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__28240\,
            I => \N__28234\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__28237\,
            I => \N__28231\
        );

    \I__4883\ : Odrv4
    port map (
            O => \N__28234\,
            I => \current_shift_inst.elapsed_time_ns_phase_22\
        );

    \I__4882\ : Odrv4
    port map (
            O => \N__28231\,
            I => \current_shift_inst.elapsed_time_ns_phase_22\
        );

    \I__4881\ : InMux
    port map (
            O => \N__28226\,
            I => \N__28223\
        );

    \I__4880\ : LocalMux
    port map (
            O => \N__28223\,
            I => \N__28220\
        );

    \I__4879\ : Span4Mux_h
    port map (
            O => \N__28220\,
            I => \N__28217\
        );

    \I__4878\ : Odrv4
    port map (
            O => \N__28217\,
            I => \current_shift_inst.z_5_22\
        );

    \I__4877\ : InMux
    port map (
            O => \N__28214\,
            I => \current_shift_inst.z_5_cry_21\
        );

    \I__4876\ : CascadeMux
    port map (
            O => \N__28211\,
            I => \N__28208\
        );

    \I__4875\ : InMux
    port map (
            O => \N__28208\,
            I => \N__28205\
        );

    \I__4874\ : LocalMux
    port map (
            O => \N__28205\,
            I => \N__28202\
        );

    \I__4873\ : Span4Mux_v
    port map (
            O => \N__28202\,
            I => \N__28199\
        );

    \I__4872\ : Odrv4
    port map (
            O => \N__28199\,
            I => \current_shift_inst.z_5_23\
        );

    \I__4871\ : InMux
    port map (
            O => \N__28196\,
            I => \current_shift_inst.z_5_cry_22\
        );

    \I__4870\ : InMux
    port map (
            O => \N__28193\,
            I => \N__28190\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__28190\,
            I => \N__28187\
        );

    \I__4868\ : Span4Mux_h
    port map (
            O => \N__28187\,
            I => \N__28184\
        );

    \I__4867\ : Odrv4
    port map (
            O => \N__28184\,
            I => \current_shift_inst.z_5_24\
        );

    \I__4866\ : InMux
    port map (
            O => \N__28181\,
            I => \current_shift_inst.z_5_cry_23\
        );

    \I__4865\ : CascadeMux
    port map (
            O => \N__28178\,
            I => \N__28175\
        );

    \I__4864\ : InMux
    port map (
            O => \N__28175\,
            I => \N__28172\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__28172\,
            I => \N__28169\
        );

    \I__4862\ : Span4Mux_h
    port map (
            O => \N__28169\,
            I => \N__28166\
        );

    \I__4861\ : Odrv4
    port map (
            O => \N__28166\,
            I => \current_shift_inst.z_5_25\
        );

    \I__4860\ : InMux
    port map (
            O => \N__28163\,
            I => \bfn_10_21_0_\
        );

    \I__4859\ : InMux
    port map (
            O => \N__28160\,
            I => \N__28157\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__28157\,
            I => \N__28154\
        );

    \I__4857\ : Span4Mux_h
    port map (
            O => \N__28154\,
            I => \N__28151\
        );

    \I__4856\ : Odrv4
    port map (
            O => \N__28151\,
            I => \current_shift_inst.z_5_26\
        );

    \I__4855\ : InMux
    port map (
            O => \N__28148\,
            I => \current_shift_inst.z_5_cry_25\
        );

    \I__4854\ : CascadeMux
    port map (
            O => \N__28145\,
            I => \N__28141\
        );

    \I__4853\ : InMux
    port map (
            O => \N__28144\,
            I => \N__28136\
        );

    \I__4852\ : InMux
    port map (
            O => \N__28141\,
            I => \N__28131\
        );

    \I__4851\ : InMux
    port map (
            O => \N__28140\,
            I => \N__28131\
        );

    \I__4850\ : InMux
    port map (
            O => \N__28139\,
            I => \N__28128\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__28136\,
            I => \N__28123\
        );

    \I__4848\ : LocalMux
    port map (
            O => \N__28131\,
            I => \N__28123\
        );

    \I__4847\ : LocalMux
    port map (
            O => \N__28128\,
            I => \N__28120\
        );

    \I__4846\ : Span4Mux_v
    port map (
            O => \N__28123\,
            I => \N__28115\
        );

    \I__4845\ : Span4Mux_h
    port map (
            O => \N__28120\,
            I => \N__28115\
        );

    \I__4844\ : Odrv4
    port map (
            O => \N__28115\,
            I => \current_shift_inst.elapsed_time_ns_phase_27\
        );

    \I__4843\ : InMux
    port map (
            O => \N__28112\,
            I => \N__28109\
        );

    \I__4842\ : LocalMux
    port map (
            O => \N__28109\,
            I => \N__28106\
        );

    \I__4841\ : Span4Mux_h
    port map (
            O => \N__28106\,
            I => \N__28103\
        );

    \I__4840\ : Odrv4
    port map (
            O => \N__28103\,
            I => \current_shift_inst.z_5_27\
        );

    \I__4839\ : InMux
    port map (
            O => \N__28100\,
            I => \current_shift_inst.z_5_cry_26\
        );

    \I__4838\ : InMux
    port map (
            O => \N__28097\,
            I => \N__28094\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__28094\,
            I => \N__28091\
        );

    \I__4836\ : Span4Mux_h
    port map (
            O => \N__28091\,
            I => \N__28088\
        );

    \I__4835\ : Odrv4
    port map (
            O => \N__28088\,
            I => \current_shift_inst.z_5_28\
        );

    \I__4834\ : InMux
    port map (
            O => \N__28085\,
            I => \current_shift_inst.z_5_cry_27\
        );

    \I__4833\ : CascadeMux
    port map (
            O => \N__28082\,
            I => \N__28079\
        );

    \I__4832\ : InMux
    port map (
            O => \N__28079\,
            I => \N__28076\
        );

    \I__4831\ : LocalMux
    port map (
            O => \N__28076\,
            I => \N__28073\
        );

    \I__4830\ : Span4Mux_h
    port map (
            O => \N__28073\,
            I => \N__28070\
        );

    \I__4829\ : Odrv4
    port map (
            O => \N__28070\,
            I => \current_shift_inst.z_5_29\
        );

    \I__4828\ : InMux
    port map (
            O => \N__28067\,
            I => \current_shift_inst.z_5_cry_28\
        );

    \I__4827\ : InMux
    port map (
            O => \N__28064\,
            I => \N__28061\
        );

    \I__4826\ : LocalMux
    port map (
            O => \N__28061\,
            I => \N__28058\
        );

    \I__4825\ : Span4Mux_h
    port map (
            O => \N__28058\,
            I => \N__28055\
        );

    \I__4824\ : Odrv4
    port map (
            O => \N__28055\,
            I => \current_shift_inst.z_5_13\
        );

    \I__4823\ : InMux
    port map (
            O => \N__28052\,
            I => \current_shift_inst.z_5_cry_12\
        );

    \I__4822\ : InMux
    port map (
            O => \N__28049\,
            I => \N__28046\
        );

    \I__4821\ : LocalMux
    port map (
            O => \N__28046\,
            I => \N__28043\
        );

    \I__4820\ : Span4Mux_h
    port map (
            O => \N__28043\,
            I => \N__28040\
        );

    \I__4819\ : Odrv4
    port map (
            O => \N__28040\,
            I => \current_shift_inst.z_5_14\
        );

    \I__4818\ : InMux
    port map (
            O => \N__28037\,
            I => \current_shift_inst.z_5_cry_13\
        );

    \I__4817\ : InMux
    port map (
            O => \N__28034\,
            I => \N__28031\
        );

    \I__4816\ : LocalMux
    port map (
            O => \N__28031\,
            I => \N__28028\
        );

    \I__4815\ : Span4Mux_v
    port map (
            O => \N__28028\,
            I => \N__28025\
        );

    \I__4814\ : Odrv4
    port map (
            O => \N__28025\,
            I => \current_shift_inst.z_5_15\
        );

    \I__4813\ : InMux
    port map (
            O => \N__28022\,
            I => \current_shift_inst.z_5_cry_14\
        );

    \I__4812\ : CascadeMux
    port map (
            O => \N__28019\,
            I => \N__28016\
        );

    \I__4811\ : InMux
    port map (
            O => \N__28016\,
            I => \N__28013\
        );

    \I__4810\ : LocalMux
    port map (
            O => \N__28013\,
            I => \N__28010\
        );

    \I__4809\ : Span4Mux_v
    port map (
            O => \N__28010\,
            I => \N__28007\
        );

    \I__4808\ : Odrv4
    port map (
            O => \N__28007\,
            I => \current_shift_inst.z_5_16\
        );

    \I__4807\ : InMux
    port map (
            O => \N__28004\,
            I => \current_shift_inst.z_5_cry_15\
        );

    \I__4806\ : InMux
    port map (
            O => \N__28001\,
            I => \N__27997\
        );

    \I__4805\ : CascadeMux
    port map (
            O => \N__28000\,
            I => \N__27994\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__27997\,
            I => \N__27989\
        );

    \I__4803\ : InMux
    port map (
            O => \N__27994\,
            I => \N__27984\
        );

    \I__4802\ : InMux
    port map (
            O => \N__27993\,
            I => \N__27984\
        );

    \I__4801\ : InMux
    port map (
            O => \N__27992\,
            I => \N__27981\
        );

    \I__4800\ : Span12Mux_s9_h
    port map (
            O => \N__27989\,
            I => \N__27976\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__27984\,
            I => \N__27976\
        );

    \I__4798\ : LocalMux
    port map (
            O => \N__27981\,
            I => \N__27973\
        );

    \I__4797\ : Odrv12
    port map (
            O => \N__27976\,
            I => \current_shift_inst.elapsed_time_ns_phase_17\
        );

    \I__4796\ : Odrv4
    port map (
            O => \N__27973\,
            I => \current_shift_inst.elapsed_time_ns_phase_17\
        );

    \I__4795\ : InMux
    port map (
            O => \N__27968\,
            I => \N__27965\
        );

    \I__4794\ : LocalMux
    port map (
            O => \N__27965\,
            I => \N__27962\
        );

    \I__4793\ : Span4Mux_v
    port map (
            O => \N__27962\,
            I => \N__27959\
        );

    \I__4792\ : Odrv4
    port map (
            O => \N__27959\,
            I => \current_shift_inst.z_5_17\
        );

    \I__4791\ : InMux
    port map (
            O => \N__27956\,
            I => \bfn_10_20_0_\
        );

    \I__4790\ : CascadeMux
    port map (
            O => \N__27953\,
            I => \N__27950\
        );

    \I__4789\ : InMux
    port map (
            O => \N__27950\,
            I => \N__27945\
        );

    \I__4788\ : InMux
    port map (
            O => \N__27949\,
            I => \N__27940\
        );

    \I__4787\ : InMux
    port map (
            O => \N__27948\,
            I => \N__27940\
        );

    \I__4786\ : LocalMux
    port map (
            O => \N__27945\,
            I => \N__27934\
        );

    \I__4785\ : LocalMux
    port map (
            O => \N__27940\,
            I => \N__27934\
        );

    \I__4784\ : InMux
    port map (
            O => \N__27939\,
            I => \N__27931\
        );

    \I__4783\ : Span4Mux_v
    port map (
            O => \N__27934\,
            I => \N__27928\
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__27931\,
            I => \N__27925\
        );

    \I__4781\ : Odrv4
    port map (
            O => \N__27928\,
            I => \current_shift_inst.elapsed_time_ns_phase_18\
        );

    \I__4780\ : Odrv4
    port map (
            O => \N__27925\,
            I => \current_shift_inst.elapsed_time_ns_phase_18\
        );

    \I__4779\ : CascadeMux
    port map (
            O => \N__27920\,
            I => \N__27917\
        );

    \I__4778\ : InMux
    port map (
            O => \N__27917\,
            I => \N__27914\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__27914\,
            I => \N__27911\
        );

    \I__4776\ : Span4Mux_h
    port map (
            O => \N__27911\,
            I => \N__27908\
        );

    \I__4775\ : Odrv4
    port map (
            O => \N__27908\,
            I => \current_shift_inst.z_5_18\
        );

    \I__4774\ : InMux
    port map (
            O => \N__27905\,
            I => \current_shift_inst.z_5_cry_17\
        );

    \I__4773\ : InMux
    port map (
            O => \N__27902\,
            I => \N__27899\
        );

    \I__4772\ : LocalMux
    port map (
            O => \N__27899\,
            I => \N__27896\
        );

    \I__4771\ : Span4Mux_h
    port map (
            O => \N__27896\,
            I => \N__27893\
        );

    \I__4770\ : Odrv4
    port map (
            O => \N__27893\,
            I => \current_shift_inst.z_5_19\
        );

    \I__4769\ : InMux
    port map (
            O => \N__27890\,
            I => \current_shift_inst.z_5_cry_18\
        );

    \I__4768\ : InMux
    port map (
            O => \N__27887\,
            I => \N__27884\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__27884\,
            I => \N__27881\
        );

    \I__4766\ : Span4Mux_v
    port map (
            O => \N__27881\,
            I => \N__27878\
        );

    \I__4765\ : Odrv4
    port map (
            O => \N__27878\,
            I => \current_shift_inst.z_5_20\
        );

    \I__4764\ : InMux
    port map (
            O => \N__27875\,
            I => \current_shift_inst.z_5_cry_19\
        );

    \I__4763\ : CascadeMux
    port map (
            O => \N__27872\,
            I => \N__27869\
        );

    \I__4762\ : InMux
    port map (
            O => \N__27869\,
            I => \N__27866\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__27866\,
            I => \N__27863\
        );

    \I__4760\ : Span4Mux_h
    port map (
            O => \N__27863\,
            I => \N__27860\
        );

    \I__4759\ : Odrv4
    port map (
            O => \N__27860\,
            I => \current_shift_inst.z_5_21\
        );

    \I__4758\ : CascadeMux
    port map (
            O => \N__27857\,
            I => \N__27854\
        );

    \I__4757\ : InMux
    port map (
            O => \N__27854\,
            I => \N__27849\
        );

    \I__4756\ : InMux
    port map (
            O => \N__27853\,
            I => \N__27846\
        );

    \I__4755\ : InMux
    port map (
            O => \N__27852\,
            I => \N__27843\
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__27849\,
            I => \N__27835\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__27846\,
            I => \N__27835\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__27843\,
            I => \N__27835\
        );

    \I__4751\ : InMux
    port map (
            O => \N__27842\,
            I => \N__27832\
        );

    \I__4750\ : Span4Mux_v
    port map (
            O => \N__27835\,
            I => \N__27829\
        );

    \I__4749\ : LocalMux
    port map (
            O => \N__27832\,
            I => \N__27826\
        );

    \I__4748\ : Odrv4
    port map (
            O => \N__27829\,
            I => \current_shift_inst.elapsed_time_ns_phase_5\
        );

    \I__4747\ : Odrv4
    port map (
            O => \N__27826\,
            I => \current_shift_inst.elapsed_time_ns_phase_5\
        );

    \I__4746\ : CascadeMux
    port map (
            O => \N__27821\,
            I => \N__27818\
        );

    \I__4745\ : InMux
    port map (
            O => \N__27818\,
            I => \N__27815\
        );

    \I__4744\ : LocalMux
    port map (
            O => \N__27815\,
            I => \N__27812\
        );

    \I__4743\ : Span4Mux_h
    port map (
            O => \N__27812\,
            I => \N__27809\
        );

    \I__4742\ : Odrv4
    port map (
            O => \N__27809\,
            I => \current_shift_inst.z_5_5\
        );

    \I__4741\ : InMux
    port map (
            O => \N__27806\,
            I => \current_shift_inst.z_5_cry_4\
        );

    \I__4740\ : InMux
    port map (
            O => \N__27803\,
            I => \N__27800\
        );

    \I__4739\ : LocalMux
    port map (
            O => \N__27800\,
            I => \N__27794\
        );

    \I__4738\ : InMux
    port map (
            O => \N__27799\,
            I => \N__27789\
        );

    \I__4737\ : InMux
    port map (
            O => \N__27798\,
            I => \N__27789\
        );

    \I__4736\ : InMux
    port map (
            O => \N__27797\,
            I => \N__27786\
        );

    \I__4735\ : Span4Mux_v
    port map (
            O => \N__27794\,
            I => \N__27783\
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__27789\,
            I => \N__27778\
        );

    \I__4733\ : LocalMux
    port map (
            O => \N__27786\,
            I => \N__27778\
        );

    \I__4732\ : Odrv4
    port map (
            O => \N__27783\,
            I => \current_shift_inst.elapsed_time_ns_phase_6\
        );

    \I__4731\ : Odrv4
    port map (
            O => \N__27778\,
            I => \current_shift_inst.elapsed_time_ns_phase_6\
        );

    \I__4730\ : InMux
    port map (
            O => \N__27773\,
            I => \N__27770\
        );

    \I__4729\ : LocalMux
    port map (
            O => \N__27770\,
            I => \N__27767\
        );

    \I__4728\ : Span4Mux_h
    port map (
            O => \N__27767\,
            I => \N__27764\
        );

    \I__4727\ : Odrv4
    port map (
            O => \N__27764\,
            I => \current_shift_inst.z_5_6\
        );

    \I__4726\ : InMux
    port map (
            O => \N__27761\,
            I => \current_shift_inst.z_5_cry_5\
        );

    \I__4725\ : CascadeMux
    port map (
            O => \N__27758\,
            I => \N__27753\
        );

    \I__4724\ : InMux
    port map (
            O => \N__27757\,
            I => \N__27749\
        );

    \I__4723\ : InMux
    port map (
            O => \N__27756\,
            I => \N__27746\
        );

    \I__4722\ : InMux
    port map (
            O => \N__27753\,
            I => \N__27741\
        );

    \I__4721\ : InMux
    port map (
            O => \N__27752\,
            I => \N__27741\
        );

    \I__4720\ : LocalMux
    port map (
            O => \N__27749\,
            I => \N__27738\
        );

    \I__4719\ : LocalMux
    port map (
            O => \N__27746\,
            I => \N__27735\
        );

    \I__4718\ : LocalMux
    port map (
            O => \N__27741\,
            I => \N__27732\
        );

    \I__4717\ : Span4Mux_v
    port map (
            O => \N__27738\,
            I => \N__27729\
        );

    \I__4716\ : Odrv12
    port map (
            O => \N__27735\,
            I => \current_shift_inst.elapsed_time_ns_phase_7\
        );

    \I__4715\ : Odrv4
    port map (
            O => \N__27732\,
            I => \current_shift_inst.elapsed_time_ns_phase_7\
        );

    \I__4714\ : Odrv4
    port map (
            O => \N__27729\,
            I => \current_shift_inst.elapsed_time_ns_phase_7\
        );

    \I__4713\ : InMux
    port map (
            O => \N__27722\,
            I => \N__27719\
        );

    \I__4712\ : LocalMux
    port map (
            O => \N__27719\,
            I => \N__27716\
        );

    \I__4711\ : Span4Mux_v
    port map (
            O => \N__27716\,
            I => \N__27713\
        );

    \I__4710\ : Odrv4
    port map (
            O => \N__27713\,
            I => \current_shift_inst.z_5_7\
        );

    \I__4709\ : InMux
    port map (
            O => \N__27710\,
            I => \current_shift_inst.z_5_cry_6\
        );

    \I__4708\ : InMux
    port map (
            O => \N__27707\,
            I => \N__27704\
        );

    \I__4707\ : LocalMux
    port map (
            O => \N__27704\,
            I => \N__27701\
        );

    \I__4706\ : Span4Mux_v
    port map (
            O => \N__27701\,
            I => \N__27698\
        );

    \I__4705\ : Odrv4
    port map (
            O => \N__27698\,
            I => \current_shift_inst.z_5_8\
        );

    \I__4704\ : InMux
    port map (
            O => \N__27695\,
            I => \current_shift_inst.z_5_cry_7\
        );

    \I__4703\ : InMux
    port map (
            O => \N__27692\,
            I => \N__27689\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__27689\,
            I => \N__27686\
        );

    \I__4701\ : Span4Mux_v
    port map (
            O => \N__27686\,
            I => \N__27683\
        );

    \I__4700\ : Odrv4
    port map (
            O => \N__27683\,
            I => \current_shift_inst.z_5_9\
        );

    \I__4699\ : InMux
    port map (
            O => \N__27680\,
            I => \bfn_10_19_0_\
        );

    \I__4698\ : InMux
    port map (
            O => \N__27677\,
            I => \N__27669\
        );

    \I__4697\ : InMux
    port map (
            O => \N__27676\,
            I => \N__27669\
        );

    \I__4696\ : InMux
    port map (
            O => \N__27675\,
            I => \N__27666\
        );

    \I__4695\ : InMux
    port map (
            O => \N__27674\,
            I => \N__27663\
        );

    \I__4694\ : LocalMux
    port map (
            O => \N__27669\,
            I => \N__27660\
        );

    \I__4693\ : LocalMux
    port map (
            O => \N__27666\,
            I => \N__27655\
        );

    \I__4692\ : LocalMux
    port map (
            O => \N__27663\,
            I => \N__27655\
        );

    \I__4691\ : Odrv12
    port map (
            O => \N__27660\,
            I => \current_shift_inst.elapsed_time_ns_phase_10\
        );

    \I__4690\ : Odrv4
    port map (
            O => \N__27655\,
            I => \current_shift_inst.elapsed_time_ns_phase_10\
        );

    \I__4689\ : CascadeMux
    port map (
            O => \N__27650\,
            I => \N__27647\
        );

    \I__4688\ : InMux
    port map (
            O => \N__27647\,
            I => \N__27644\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__27644\,
            I => \N__27641\
        );

    \I__4686\ : Span4Mux_h
    port map (
            O => \N__27641\,
            I => \N__27638\
        );

    \I__4685\ : Odrv4
    port map (
            O => \N__27638\,
            I => \current_shift_inst.z_5_10\
        );

    \I__4684\ : InMux
    port map (
            O => \N__27635\,
            I => \current_shift_inst.z_5_cry_9\
        );

    \I__4683\ : InMux
    port map (
            O => \N__27632\,
            I => \N__27629\
        );

    \I__4682\ : LocalMux
    port map (
            O => \N__27629\,
            I => \N__27626\
        );

    \I__4681\ : Span4Mux_h
    port map (
            O => \N__27626\,
            I => \N__27623\
        );

    \I__4680\ : Odrv4
    port map (
            O => \N__27623\,
            I => \current_shift_inst.z_5_11\
        );

    \I__4679\ : InMux
    port map (
            O => \N__27620\,
            I => \current_shift_inst.z_5_cry_10\
        );

    \I__4678\ : InMux
    port map (
            O => \N__27617\,
            I => \N__27614\
        );

    \I__4677\ : LocalMux
    port map (
            O => \N__27614\,
            I => \N__27611\
        );

    \I__4676\ : Span4Mux_h
    port map (
            O => \N__27611\,
            I => \N__27608\
        );

    \I__4675\ : Odrv4
    port map (
            O => \N__27608\,
            I => \current_shift_inst.z_5_12\
        );

    \I__4674\ : InMux
    port map (
            O => \N__27605\,
            I => \current_shift_inst.z_5_cry_11\
        );

    \I__4673\ : InMux
    port map (
            O => \N__27602\,
            I => \current_shift_inst.z_cry_30\
        );

    \I__4672\ : InMux
    port map (
            O => \N__27599\,
            I => \N__27592\
        );

    \I__4671\ : InMux
    port map (
            O => \N__27598\,
            I => \N__27582\
        );

    \I__4670\ : InMux
    port map (
            O => \N__27597\,
            I => \N__27582\
        );

    \I__4669\ : InMux
    port map (
            O => \N__27596\,
            I => \N__27582\
        );

    \I__4668\ : InMux
    port map (
            O => \N__27595\,
            I => \N__27582\
        );

    \I__4667\ : LocalMux
    port map (
            O => \N__27592\,
            I => \N__27579\
        );

    \I__4666\ : InMux
    port map (
            O => \N__27591\,
            I => \N__27576\
        );

    \I__4665\ : LocalMux
    port map (
            O => \N__27582\,
            I => \current_shift_inst.elapsed_time_ns_phase_1\
        );

    \I__4664\ : Odrv4
    port map (
            O => \N__27579\,
            I => \current_shift_inst.elapsed_time_ns_phase_1\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__27576\,
            I => \current_shift_inst.elapsed_time_ns_phase_1\
        );

    \I__4662\ : CascadeMux
    port map (
            O => \N__27569\,
            I => \N__27565\
        );

    \I__4661\ : InMux
    port map (
            O => \N__27568\,
            I => \N__27560\
        );

    \I__4660\ : InMux
    port map (
            O => \N__27565\,
            I => \N__27555\
        );

    \I__4659\ : InMux
    port map (
            O => \N__27564\,
            I => \N__27555\
        );

    \I__4658\ : InMux
    port map (
            O => \N__27563\,
            I => \N__27552\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__27560\,
            I => \current_shift_inst.elapsed_time_ns_phase_2\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__27555\,
            I => \current_shift_inst.elapsed_time_ns_phase_2\
        );

    \I__4655\ : LocalMux
    port map (
            O => \N__27552\,
            I => \current_shift_inst.elapsed_time_ns_phase_2\
        );

    \I__4654\ : CascadeMux
    port map (
            O => \N__27545\,
            I => \N__27542\
        );

    \I__4653\ : InMux
    port map (
            O => \N__27542\,
            I => \N__27539\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__27539\,
            I => \N__27536\
        );

    \I__4651\ : Span4Mux_h
    port map (
            O => \N__27536\,
            I => \N__27533\
        );

    \I__4650\ : Odrv4
    port map (
            O => \N__27533\,
            I => \current_shift_inst.z_5_2\
        );

    \I__4649\ : InMux
    port map (
            O => \N__27530\,
            I => \current_shift_inst.z_5_cry_1\
        );

    \I__4648\ : InMux
    port map (
            O => \N__27527\,
            I => \N__27521\
        );

    \I__4647\ : InMux
    port map (
            O => \N__27526\,
            I => \N__27521\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__27521\,
            I => \N__27517\
        );

    \I__4645\ : InMux
    port map (
            O => \N__27520\,
            I => \N__27514\
        );

    \I__4644\ : Span4Mux_h
    port map (
            O => \N__27517\,
            I => \N__27509\
        );

    \I__4643\ : LocalMux
    port map (
            O => \N__27514\,
            I => \N__27509\
        );

    \I__4642\ : Odrv4
    port map (
            O => \N__27509\,
            I => \current_shift_inst.elapsed_time_ns_phase_3\
        );

    \I__4641\ : CascadeMux
    port map (
            O => \N__27506\,
            I => \N__27503\
        );

    \I__4640\ : InMux
    port map (
            O => \N__27503\,
            I => \N__27500\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__27500\,
            I => \N__27497\
        );

    \I__4638\ : Span4Mux_h
    port map (
            O => \N__27497\,
            I => \N__27494\
        );

    \I__4637\ : Odrv4
    port map (
            O => \N__27494\,
            I => \current_shift_inst.z_5_3\
        );

    \I__4636\ : InMux
    port map (
            O => \N__27491\,
            I => \current_shift_inst.z_5_cry_2\
        );

    \I__4635\ : InMux
    port map (
            O => \N__27488\,
            I => \N__27480\
        );

    \I__4634\ : InMux
    port map (
            O => \N__27487\,
            I => \N__27480\
        );

    \I__4633\ : InMux
    port map (
            O => \N__27486\,
            I => \N__27477\
        );

    \I__4632\ : InMux
    port map (
            O => \N__27485\,
            I => \N__27474\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__27480\,
            I => \N__27469\
        );

    \I__4630\ : LocalMux
    port map (
            O => \N__27477\,
            I => \N__27469\
        );

    \I__4629\ : LocalMux
    port map (
            O => \N__27474\,
            I => \N__27466\
        );

    \I__4628\ : Span4Mux_v
    port map (
            O => \N__27469\,
            I => \N__27461\
        );

    \I__4627\ : Span4Mux_h
    port map (
            O => \N__27466\,
            I => \N__27461\
        );

    \I__4626\ : Odrv4
    port map (
            O => \N__27461\,
            I => \current_shift_inst.elapsed_time_ns_phase_4\
        );

    \I__4625\ : InMux
    port map (
            O => \N__27458\,
            I => \N__27455\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__27455\,
            I => \N__27452\
        );

    \I__4623\ : Span4Mux_h
    port map (
            O => \N__27452\,
            I => \N__27449\
        );

    \I__4622\ : Odrv4
    port map (
            O => \N__27449\,
            I => \current_shift_inst.z_5_4\
        );

    \I__4621\ : InMux
    port map (
            O => \N__27446\,
            I => \current_shift_inst.z_5_cry_3\
        );

    \I__4620\ : InMux
    port map (
            O => \N__27443\,
            I => \N__27440\
        );

    \I__4619\ : LocalMux
    port map (
            O => \N__27440\,
            I => \G_406\
        );

    \I__4618\ : CascadeMux
    port map (
            O => \N__27437\,
            I => \N__27434\
        );

    \I__4617\ : InMux
    port map (
            O => \N__27434\,
            I => \N__27431\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__27431\,
            I => \N__27428\
        );

    \I__4615\ : Span4Mux_h
    port map (
            O => \N__27428\,
            I => \N__27425\
        );

    \I__4614\ : Odrv4
    port map (
            O => \N__27425\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\
        );

    \I__4613\ : CascadeMux
    port map (
            O => \N__27422\,
            I => \N__27419\
        );

    \I__4612\ : InMux
    port map (
            O => \N__27419\,
            I => \N__27416\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__27416\,
            I => \N__27413\
        );

    \I__4610\ : Odrv4
    port map (
            O => \N__27413\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\
        );

    \I__4609\ : CascadeMux
    port map (
            O => \N__27410\,
            I => \N__27407\
        );

    \I__4608\ : InMux
    port map (
            O => \N__27407\,
            I => \N__27404\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__27404\,
            I => \N__27401\
        );

    \I__4606\ : Odrv4
    port map (
            O => \N__27401\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\
        );

    \I__4605\ : InMux
    port map (
            O => \N__27398\,
            I => \N__27394\
        );

    \I__4604\ : InMux
    port map (
            O => \N__27397\,
            I => \N__27390\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__27394\,
            I => \N__27386\
        );

    \I__4602\ : InMux
    port map (
            O => \N__27393\,
            I => \N__27383\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__27390\,
            I => \N__27380\
        );

    \I__4600\ : InMux
    port map (
            O => \N__27389\,
            I => \N__27377\
        );

    \I__4599\ : Odrv4
    port map (
            O => \N__27386\,
            I => \phase_controller_inst1.stoper_hc.time_passed11\
        );

    \I__4598\ : LocalMux
    port map (
            O => \N__27383\,
            I => \phase_controller_inst1.stoper_hc.time_passed11\
        );

    \I__4597\ : Odrv12
    port map (
            O => \N__27380\,
            I => \phase_controller_inst1.stoper_hc.time_passed11\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__27377\,
            I => \phase_controller_inst1.stoper_hc.time_passed11\
        );

    \I__4595\ : CascadeMux
    port map (
            O => \N__27368\,
            I => \N__27365\
        );

    \I__4594\ : InMux
    port map (
            O => \N__27365\,
            I => \N__27362\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__27362\,
            I => \N__27359\
        );

    \I__4592\ : Odrv4
    port map (
            O => \N__27359\,
            I => \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa\
        );

    \I__4591\ : CascadeMux
    port map (
            O => \N__27356\,
            I => \N__27353\
        );

    \I__4590\ : InMux
    port map (
            O => \N__27353\,
            I => \N__27350\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__27350\,
            I => \G_407\
        );

    \I__4588\ : InMux
    port map (
            O => \N__27347\,
            I => \N__27342\
        );

    \I__4587\ : InMux
    port map (
            O => \N__27346\,
            I => \N__27339\
        );

    \I__4586\ : InMux
    port map (
            O => \N__27345\,
            I => \N__27336\
        );

    \I__4585\ : LocalMux
    port map (
            O => \N__27342\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__4584\ : LocalMux
    port map (
            O => \N__27339\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__27336\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__4582\ : InMux
    port map (
            O => \N__27329\,
            I => \pwm_generator_inst.counter_cry_5\
        );

    \I__4581\ : InMux
    port map (
            O => \N__27326\,
            I => \N__27321\
        );

    \I__4580\ : InMux
    port map (
            O => \N__27325\,
            I => \N__27318\
        );

    \I__4579\ : InMux
    port map (
            O => \N__27324\,
            I => \N__27315\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__27321\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__27318\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__4576\ : LocalMux
    port map (
            O => \N__27315\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__4575\ : InMux
    port map (
            O => \N__27308\,
            I => \pwm_generator_inst.counter_cry_6\
        );

    \I__4574\ : InMux
    port map (
            O => \N__27305\,
            I => \N__27300\
        );

    \I__4573\ : InMux
    port map (
            O => \N__27304\,
            I => \N__27297\
        );

    \I__4572\ : InMux
    port map (
            O => \N__27303\,
            I => \N__27294\
        );

    \I__4571\ : LocalMux
    port map (
            O => \N__27300\,
            I => \N__27291\
        );

    \I__4570\ : LocalMux
    port map (
            O => \N__27297\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__4569\ : LocalMux
    port map (
            O => \N__27294\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__4568\ : Odrv4
    port map (
            O => \N__27291\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__4567\ : InMux
    port map (
            O => \N__27284\,
            I => \bfn_10_10_0_\
        );

    \I__4566\ : InMux
    port map (
            O => \N__27281\,
            I => \N__27269\
        );

    \I__4565\ : InMux
    port map (
            O => \N__27280\,
            I => \N__27266\
        );

    \I__4564\ : InMux
    port map (
            O => \N__27279\,
            I => \N__27257\
        );

    \I__4563\ : InMux
    port map (
            O => \N__27278\,
            I => \N__27257\
        );

    \I__4562\ : InMux
    port map (
            O => \N__27277\,
            I => \N__27257\
        );

    \I__4561\ : InMux
    port map (
            O => \N__27276\,
            I => \N__27257\
        );

    \I__4560\ : InMux
    port map (
            O => \N__27275\,
            I => \N__27248\
        );

    \I__4559\ : InMux
    port map (
            O => \N__27274\,
            I => \N__27248\
        );

    \I__4558\ : InMux
    port map (
            O => \N__27273\,
            I => \N__27248\
        );

    \I__4557\ : InMux
    port map (
            O => \N__27272\,
            I => \N__27248\
        );

    \I__4556\ : LocalMux
    port map (
            O => \N__27269\,
            I => \N__27245\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__27266\,
            I => \N__27242\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__27257\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__4553\ : LocalMux
    port map (
            O => \N__27248\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__4552\ : Odrv12
    port map (
            O => \N__27245\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__4551\ : Odrv4
    port map (
            O => \N__27242\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__4550\ : InMux
    port map (
            O => \N__27233\,
            I => \pwm_generator_inst.counter_cry_8\
        );

    \I__4549\ : InMux
    port map (
            O => \N__27230\,
            I => \N__27225\
        );

    \I__4548\ : InMux
    port map (
            O => \N__27229\,
            I => \N__27222\
        );

    \I__4547\ : InMux
    port map (
            O => \N__27228\,
            I => \N__27219\
        );

    \I__4546\ : LocalMux
    port map (
            O => \N__27225\,
            I => \N__27216\
        );

    \I__4545\ : LocalMux
    port map (
            O => \N__27222\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__27219\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__4543\ : Odrv4
    port map (
            O => \N__27216\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__4542\ : CascadeMux
    port map (
            O => \N__27209\,
            I => \pwm_generator_inst.un1_counterlto2_0_cascade_\
        );

    \I__4541\ : CascadeMux
    port map (
            O => \N__27206\,
            I => \pwm_generator_inst.un1_counterlt9_cascade_\
        );

    \I__4540\ : InMux
    port map (
            O => \N__27203\,
            I => \N__27200\
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__27200\,
            I => \pwm_generator_inst.un1_counterlto9_2\
        );

    \I__4538\ : InMux
    port map (
            O => \N__27197\,
            I => \N__27192\
        );

    \I__4537\ : InMux
    port map (
            O => \N__27196\,
            I => \N__27189\
        );

    \I__4536\ : InMux
    port map (
            O => \N__27195\,
            I => \N__27186\
        );

    \I__4535\ : LocalMux
    port map (
            O => \N__27192\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__4534\ : LocalMux
    port map (
            O => \N__27189\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__4533\ : LocalMux
    port map (
            O => \N__27186\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__4532\ : InMux
    port map (
            O => \N__27179\,
            I => \bfn_10_9_0_\
        );

    \I__4531\ : InMux
    port map (
            O => \N__27176\,
            I => \N__27171\
        );

    \I__4530\ : InMux
    port map (
            O => \N__27175\,
            I => \N__27168\
        );

    \I__4529\ : InMux
    port map (
            O => \N__27174\,
            I => \N__27165\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__27171\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__27168\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__4526\ : LocalMux
    port map (
            O => \N__27165\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__4525\ : InMux
    port map (
            O => \N__27158\,
            I => \pwm_generator_inst.counter_cry_0\
        );

    \I__4524\ : InMux
    port map (
            O => \N__27155\,
            I => \N__27150\
        );

    \I__4523\ : InMux
    port map (
            O => \N__27154\,
            I => \N__27147\
        );

    \I__4522\ : InMux
    port map (
            O => \N__27153\,
            I => \N__27144\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__27150\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__27147\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__4519\ : LocalMux
    port map (
            O => \N__27144\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__4518\ : InMux
    port map (
            O => \N__27137\,
            I => \pwm_generator_inst.counter_cry_1\
        );

    \I__4517\ : InMux
    port map (
            O => \N__27134\,
            I => \N__27129\
        );

    \I__4516\ : InMux
    port map (
            O => \N__27133\,
            I => \N__27126\
        );

    \I__4515\ : InMux
    port map (
            O => \N__27132\,
            I => \N__27123\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__27129\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__27126\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__27123\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__4511\ : InMux
    port map (
            O => \N__27116\,
            I => \pwm_generator_inst.counter_cry_2\
        );

    \I__4510\ : InMux
    port map (
            O => \N__27113\,
            I => \N__27108\
        );

    \I__4509\ : InMux
    port map (
            O => \N__27112\,
            I => \N__27105\
        );

    \I__4508\ : InMux
    port map (
            O => \N__27111\,
            I => \N__27102\
        );

    \I__4507\ : LocalMux
    port map (
            O => \N__27108\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__4506\ : LocalMux
    port map (
            O => \N__27105\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__27102\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__4504\ : InMux
    port map (
            O => \N__27095\,
            I => \pwm_generator_inst.counter_cry_3\
        );

    \I__4503\ : InMux
    port map (
            O => \N__27092\,
            I => \N__27087\
        );

    \I__4502\ : InMux
    port map (
            O => \N__27091\,
            I => \N__27084\
        );

    \I__4501\ : InMux
    port map (
            O => \N__27090\,
            I => \N__27081\
        );

    \I__4500\ : LocalMux
    port map (
            O => \N__27087\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__4499\ : LocalMux
    port map (
            O => \N__27084\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__4498\ : LocalMux
    port map (
            O => \N__27081\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__4497\ : InMux
    port map (
            O => \N__27074\,
            I => \pwm_generator_inst.counter_cry_4\
        );

    \I__4496\ : InMux
    port map (
            O => \N__27071\,
            I => \N__27067\
        );

    \I__4495\ : InMux
    port map (
            O => \N__27070\,
            I => \N__27064\
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__27067\,
            I => \N__27058\
        );

    \I__4493\ : LocalMux
    port map (
            O => \N__27064\,
            I => \N__27058\
        );

    \I__4492\ : InMux
    port map (
            O => \N__27063\,
            I => \N__27055\
        );

    \I__4491\ : Span4Mux_v
    port map (
            O => \N__27058\,
            I => \N__27052\
        );

    \I__4490\ : LocalMux
    port map (
            O => \N__27055\,
            I => \current_shift_inst.timer_phase.counterZ0Z_24\
        );

    \I__4489\ : Odrv4
    port map (
            O => \N__27052\,
            I => \current_shift_inst.timer_phase.counterZ0Z_24\
        );

    \I__4488\ : InMux
    port map (
            O => \N__27047\,
            I => \bfn_9_28_0_\
        );

    \I__4487\ : InMux
    port map (
            O => \N__27044\,
            I => \N__27040\
        );

    \I__4486\ : InMux
    port map (
            O => \N__27043\,
            I => \N__27037\
        );

    \I__4485\ : LocalMux
    port map (
            O => \N__27040\,
            I => \N__27031\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__27037\,
            I => \N__27031\
        );

    \I__4483\ : InMux
    port map (
            O => \N__27036\,
            I => \N__27028\
        );

    \I__4482\ : Span4Mux_v
    port map (
            O => \N__27031\,
            I => \N__27025\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__27028\,
            I => \current_shift_inst.timer_phase.counterZ0Z_25\
        );

    \I__4480\ : Odrv4
    port map (
            O => \N__27025\,
            I => \current_shift_inst.timer_phase.counterZ0Z_25\
        );

    \I__4479\ : InMux
    port map (
            O => \N__27020\,
            I => \current_shift_inst.timer_phase.counter_cry_24\
        );

    \I__4478\ : CascadeMux
    port map (
            O => \N__27017\,
            I => \N__27013\
        );

    \I__4477\ : CascadeMux
    port map (
            O => \N__27016\,
            I => \N__27010\
        );

    \I__4476\ : InMux
    port map (
            O => \N__27013\,
            I => \N__27005\
        );

    \I__4475\ : InMux
    port map (
            O => \N__27010\,
            I => \N__27005\
        );

    \I__4474\ : LocalMux
    port map (
            O => \N__27005\,
            I => \N__27001\
        );

    \I__4473\ : InMux
    port map (
            O => \N__27004\,
            I => \N__26998\
        );

    \I__4472\ : Span4Mux_h
    port map (
            O => \N__27001\,
            I => \N__26995\
        );

    \I__4471\ : LocalMux
    port map (
            O => \N__26998\,
            I => \current_shift_inst.timer_phase.counterZ0Z_26\
        );

    \I__4470\ : Odrv4
    port map (
            O => \N__26995\,
            I => \current_shift_inst.timer_phase.counterZ0Z_26\
        );

    \I__4469\ : InMux
    port map (
            O => \N__26990\,
            I => \current_shift_inst.timer_phase.counter_cry_25\
        );

    \I__4468\ : CascadeMux
    port map (
            O => \N__26987\,
            I => \N__26983\
        );

    \I__4467\ : CascadeMux
    port map (
            O => \N__26986\,
            I => \N__26980\
        );

    \I__4466\ : InMux
    port map (
            O => \N__26983\,
            I => \N__26974\
        );

    \I__4465\ : InMux
    port map (
            O => \N__26980\,
            I => \N__26974\
        );

    \I__4464\ : InMux
    port map (
            O => \N__26979\,
            I => \N__26971\
        );

    \I__4463\ : LocalMux
    port map (
            O => \N__26974\,
            I => \N__26968\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__26971\,
            I => \current_shift_inst.timer_phase.counterZ0Z_27\
        );

    \I__4461\ : Odrv12
    port map (
            O => \N__26968\,
            I => \current_shift_inst.timer_phase.counterZ0Z_27\
        );

    \I__4460\ : InMux
    port map (
            O => \N__26963\,
            I => \current_shift_inst.timer_phase.counter_cry_26\
        );

    \I__4459\ : InMux
    port map (
            O => \N__26960\,
            I => \N__26957\
        );

    \I__4458\ : LocalMux
    port map (
            O => \N__26957\,
            I => \N__26953\
        );

    \I__4457\ : InMux
    port map (
            O => \N__26956\,
            I => \N__26950\
        );

    \I__4456\ : Span4Mux_h
    port map (
            O => \N__26953\,
            I => \N__26947\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__26950\,
            I => \current_shift_inst.timer_phase.counterZ0Z_28\
        );

    \I__4454\ : Odrv4
    port map (
            O => \N__26947\,
            I => \current_shift_inst.timer_phase.counterZ0Z_28\
        );

    \I__4453\ : InMux
    port map (
            O => \N__26942\,
            I => \current_shift_inst.timer_phase.counter_cry_27\
        );

    \I__4452\ : InMux
    port map (
            O => \N__26939\,
            I => \current_shift_inst.timer_phase.counter_cry_28\
        );

    \I__4451\ : InMux
    port map (
            O => \N__26936\,
            I => \N__26932\
        );

    \I__4450\ : InMux
    port map (
            O => \N__26935\,
            I => \N__26929\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__26932\,
            I => \N__26926\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__26929\,
            I => \current_shift_inst.timer_phase.counterZ0Z_29\
        );

    \I__4447\ : Odrv12
    port map (
            O => \N__26926\,
            I => \current_shift_inst.timer_phase.counterZ0Z_29\
        );

    \I__4446\ : InMux
    port map (
            O => \N__26921\,
            I => \N__26918\
        );

    \I__4445\ : LocalMux
    port map (
            O => \N__26918\,
            I => \il_max_comp1_D1\
        );

    \I__4444\ : InMux
    port map (
            O => \N__26915\,
            I => \N__26911\
        );

    \I__4443\ : InMux
    port map (
            O => \N__26914\,
            I => \N__26908\
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__26911\,
            I => \N__26902\
        );

    \I__4441\ : LocalMux
    port map (
            O => \N__26908\,
            I => \N__26902\
        );

    \I__4440\ : InMux
    port map (
            O => \N__26907\,
            I => \N__26899\
        );

    \I__4439\ : Span4Mux_v
    port map (
            O => \N__26902\,
            I => \N__26896\
        );

    \I__4438\ : LocalMux
    port map (
            O => \N__26899\,
            I => \current_shift_inst.timer_phase.counterZ0Z_16\
        );

    \I__4437\ : Odrv4
    port map (
            O => \N__26896\,
            I => \current_shift_inst.timer_phase.counterZ0Z_16\
        );

    \I__4436\ : InMux
    port map (
            O => \N__26891\,
            I => \bfn_9_27_0_\
        );

    \I__4435\ : InMux
    port map (
            O => \N__26888\,
            I => \N__26884\
        );

    \I__4434\ : InMux
    port map (
            O => \N__26887\,
            I => \N__26881\
        );

    \I__4433\ : LocalMux
    port map (
            O => \N__26884\,
            I => \N__26875\
        );

    \I__4432\ : LocalMux
    port map (
            O => \N__26881\,
            I => \N__26875\
        );

    \I__4431\ : InMux
    port map (
            O => \N__26880\,
            I => \N__26872\
        );

    \I__4430\ : Span4Mux_v
    port map (
            O => \N__26875\,
            I => \N__26869\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__26872\,
            I => \current_shift_inst.timer_phase.counterZ0Z_17\
        );

    \I__4428\ : Odrv4
    port map (
            O => \N__26869\,
            I => \current_shift_inst.timer_phase.counterZ0Z_17\
        );

    \I__4427\ : InMux
    port map (
            O => \N__26864\,
            I => \current_shift_inst.timer_phase.counter_cry_16\
        );

    \I__4426\ : CascadeMux
    port map (
            O => \N__26861\,
            I => \N__26857\
        );

    \I__4425\ : CascadeMux
    port map (
            O => \N__26860\,
            I => \N__26854\
        );

    \I__4424\ : InMux
    port map (
            O => \N__26857\,
            I => \N__26849\
        );

    \I__4423\ : InMux
    port map (
            O => \N__26854\,
            I => \N__26849\
        );

    \I__4422\ : LocalMux
    port map (
            O => \N__26849\,
            I => \N__26845\
        );

    \I__4421\ : InMux
    port map (
            O => \N__26848\,
            I => \N__26842\
        );

    \I__4420\ : Span4Mux_h
    port map (
            O => \N__26845\,
            I => \N__26839\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__26842\,
            I => \current_shift_inst.timer_phase.counterZ0Z_18\
        );

    \I__4418\ : Odrv4
    port map (
            O => \N__26839\,
            I => \current_shift_inst.timer_phase.counterZ0Z_18\
        );

    \I__4417\ : InMux
    port map (
            O => \N__26834\,
            I => \current_shift_inst.timer_phase.counter_cry_17\
        );

    \I__4416\ : CascadeMux
    port map (
            O => \N__26831\,
            I => \N__26827\
        );

    \I__4415\ : CascadeMux
    port map (
            O => \N__26830\,
            I => \N__26824\
        );

    \I__4414\ : InMux
    port map (
            O => \N__26827\,
            I => \N__26819\
        );

    \I__4413\ : InMux
    port map (
            O => \N__26824\,
            I => \N__26819\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__26819\,
            I => \N__26815\
        );

    \I__4411\ : InMux
    port map (
            O => \N__26818\,
            I => \N__26812\
        );

    \I__4410\ : Span4Mux_h
    port map (
            O => \N__26815\,
            I => \N__26809\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__26812\,
            I => \current_shift_inst.timer_phase.counterZ0Z_19\
        );

    \I__4408\ : Odrv4
    port map (
            O => \N__26809\,
            I => \current_shift_inst.timer_phase.counterZ0Z_19\
        );

    \I__4407\ : InMux
    port map (
            O => \N__26804\,
            I => \current_shift_inst.timer_phase.counter_cry_18\
        );

    \I__4406\ : InMux
    port map (
            O => \N__26801\,
            I => \N__26795\
        );

    \I__4405\ : InMux
    port map (
            O => \N__26800\,
            I => \N__26795\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__26795\,
            I => \N__26791\
        );

    \I__4403\ : InMux
    port map (
            O => \N__26794\,
            I => \N__26788\
        );

    \I__4402\ : Span4Mux_h
    port map (
            O => \N__26791\,
            I => \N__26785\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__26788\,
            I => \current_shift_inst.timer_phase.counterZ0Z_20\
        );

    \I__4400\ : Odrv4
    port map (
            O => \N__26785\,
            I => \current_shift_inst.timer_phase.counterZ0Z_20\
        );

    \I__4399\ : InMux
    port map (
            O => \N__26780\,
            I => \current_shift_inst.timer_phase.counter_cry_19\
        );

    \I__4398\ : InMux
    port map (
            O => \N__26777\,
            I => \N__26771\
        );

    \I__4397\ : InMux
    port map (
            O => \N__26776\,
            I => \N__26771\
        );

    \I__4396\ : LocalMux
    port map (
            O => \N__26771\,
            I => \N__26767\
        );

    \I__4395\ : InMux
    port map (
            O => \N__26770\,
            I => \N__26764\
        );

    \I__4394\ : Span4Mux_h
    port map (
            O => \N__26767\,
            I => \N__26761\
        );

    \I__4393\ : LocalMux
    port map (
            O => \N__26764\,
            I => \current_shift_inst.timer_phase.counterZ0Z_21\
        );

    \I__4392\ : Odrv4
    port map (
            O => \N__26761\,
            I => \current_shift_inst.timer_phase.counterZ0Z_21\
        );

    \I__4391\ : InMux
    port map (
            O => \N__26756\,
            I => \current_shift_inst.timer_phase.counter_cry_20\
        );

    \I__4390\ : CascadeMux
    port map (
            O => \N__26753\,
            I => \N__26749\
        );

    \I__4389\ : CascadeMux
    port map (
            O => \N__26752\,
            I => \N__26746\
        );

    \I__4388\ : InMux
    port map (
            O => \N__26749\,
            I => \N__26741\
        );

    \I__4387\ : InMux
    port map (
            O => \N__26746\,
            I => \N__26741\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__26741\,
            I => \N__26737\
        );

    \I__4385\ : InMux
    port map (
            O => \N__26740\,
            I => \N__26734\
        );

    \I__4384\ : Span4Mux_v
    port map (
            O => \N__26737\,
            I => \N__26731\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__26734\,
            I => \current_shift_inst.timer_phase.counterZ0Z_22\
        );

    \I__4382\ : Odrv4
    port map (
            O => \N__26731\,
            I => \current_shift_inst.timer_phase.counterZ0Z_22\
        );

    \I__4381\ : InMux
    port map (
            O => \N__26726\,
            I => \current_shift_inst.timer_phase.counter_cry_21\
        );

    \I__4380\ : CascadeMux
    port map (
            O => \N__26723\,
            I => \N__26719\
        );

    \I__4379\ : CascadeMux
    port map (
            O => \N__26722\,
            I => \N__26716\
        );

    \I__4378\ : InMux
    port map (
            O => \N__26719\,
            I => \N__26710\
        );

    \I__4377\ : InMux
    port map (
            O => \N__26716\,
            I => \N__26710\
        );

    \I__4376\ : InMux
    port map (
            O => \N__26715\,
            I => \N__26707\
        );

    \I__4375\ : LocalMux
    port map (
            O => \N__26710\,
            I => \N__26704\
        );

    \I__4374\ : LocalMux
    port map (
            O => \N__26707\,
            I => \current_shift_inst.timer_phase.counterZ0Z_23\
        );

    \I__4373\ : Odrv12
    port map (
            O => \N__26704\,
            I => \current_shift_inst.timer_phase.counterZ0Z_23\
        );

    \I__4372\ : InMux
    port map (
            O => \N__26699\,
            I => \current_shift_inst.timer_phase.counter_cry_22\
        );

    \I__4371\ : CascadeMux
    port map (
            O => \N__26696\,
            I => \N__26692\
        );

    \I__4370\ : InMux
    port map (
            O => \N__26695\,
            I => \N__26689\
        );

    \I__4369\ : InMux
    port map (
            O => \N__26692\,
            I => \N__26686\
        );

    \I__4368\ : LocalMux
    port map (
            O => \N__26689\,
            I => \N__26680\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__26686\,
            I => \N__26680\
        );

    \I__4366\ : InMux
    port map (
            O => \N__26685\,
            I => \N__26677\
        );

    \I__4365\ : Span4Mux_v
    port map (
            O => \N__26680\,
            I => \N__26674\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__26677\,
            I => \current_shift_inst.timer_phase.counterZ0Z_8\
        );

    \I__4363\ : Odrv4
    port map (
            O => \N__26674\,
            I => \current_shift_inst.timer_phase.counterZ0Z_8\
        );

    \I__4362\ : InMux
    port map (
            O => \N__26669\,
            I => \bfn_9_26_0_\
        );

    \I__4361\ : InMux
    port map (
            O => \N__26666\,
            I => \N__26662\
        );

    \I__4360\ : InMux
    port map (
            O => \N__26665\,
            I => \N__26659\
        );

    \I__4359\ : LocalMux
    port map (
            O => \N__26662\,
            I => \N__26653\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__26659\,
            I => \N__26653\
        );

    \I__4357\ : InMux
    port map (
            O => \N__26658\,
            I => \N__26650\
        );

    \I__4356\ : Span4Mux_v
    port map (
            O => \N__26653\,
            I => \N__26647\
        );

    \I__4355\ : LocalMux
    port map (
            O => \N__26650\,
            I => \current_shift_inst.timer_phase.counterZ0Z_9\
        );

    \I__4354\ : Odrv4
    port map (
            O => \N__26647\,
            I => \current_shift_inst.timer_phase.counterZ0Z_9\
        );

    \I__4353\ : InMux
    port map (
            O => \N__26642\,
            I => \current_shift_inst.timer_phase.counter_cry_8\
        );

    \I__4352\ : CascadeMux
    port map (
            O => \N__26639\,
            I => \N__26635\
        );

    \I__4351\ : CascadeMux
    port map (
            O => \N__26638\,
            I => \N__26632\
        );

    \I__4350\ : InMux
    port map (
            O => \N__26635\,
            I => \N__26627\
        );

    \I__4349\ : InMux
    port map (
            O => \N__26632\,
            I => \N__26627\
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__26627\,
            I => \N__26623\
        );

    \I__4347\ : InMux
    port map (
            O => \N__26626\,
            I => \N__26620\
        );

    \I__4346\ : Span4Mux_h
    port map (
            O => \N__26623\,
            I => \N__26617\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__26620\,
            I => \current_shift_inst.timer_phase.counterZ0Z_10\
        );

    \I__4344\ : Odrv4
    port map (
            O => \N__26617\,
            I => \current_shift_inst.timer_phase.counterZ0Z_10\
        );

    \I__4343\ : InMux
    port map (
            O => \N__26612\,
            I => \current_shift_inst.timer_phase.counter_cry_9\
        );

    \I__4342\ : CascadeMux
    port map (
            O => \N__26609\,
            I => \N__26605\
        );

    \I__4341\ : CascadeMux
    port map (
            O => \N__26608\,
            I => \N__26602\
        );

    \I__4340\ : InMux
    port map (
            O => \N__26605\,
            I => \N__26596\
        );

    \I__4339\ : InMux
    port map (
            O => \N__26602\,
            I => \N__26596\
        );

    \I__4338\ : InMux
    port map (
            O => \N__26601\,
            I => \N__26593\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__26596\,
            I => \N__26590\
        );

    \I__4336\ : LocalMux
    port map (
            O => \N__26593\,
            I => \current_shift_inst.timer_phase.counterZ0Z_11\
        );

    \I__4335\ : Odrv12
    port map (
            O => \N__26590\,
            I => \current_shift_inst.timer_phase.counterZ0Z_11\
        );

    \I__4334\ : InMux
    port map (
            O => \N__26585\,
            I => \current_shift_inst.timer_phase.counter_cry_10\
        );

    \I__4333\ : InMux
    port map (
            O => \N__26582\,
            I => \N__26575\
        );

    \I__4332\ : InMux
    port map (
            O => \N__26581\,
            I => \N__26575\
        );

    \I__4331\ : InMux
    port map (
            O => \N__26580\,
            I => \N__26572\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__26575\,
            I => \N__26569\
        );

    \I__4329\ : LocalMux
    port map (
            O => \N__26572\,
            I => \current_shift_inst.timer_phase.counterZ0Z_12\
        );

    \I__4328\ : Odrv12
    port map (
            O => \N__26569\,
            I => \current_shift_inst.timer_phase.counterZ0Z_12\
        );

    \I__4327\ : InMux
    port map (
            O => \N__26564\,
            I => \current_shift_inst.timer_phase.counter_cry_11\
        );

    \I__4326\ : InMux
    port map (
            O => \N__26561\,
            I => \N__26555\
        );

    \I__4325\ : InMux
    port map (
            O => \N__26560\,
            I => \N__26555\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__26555\,
            I => \N__26551\
        );

    \I__4323\ : InMux
    port map (
            O => \N__26554\,
            I => \N__26548\
        );

    \I__4322\ : Span4Mux_h
    port map (
            O => \N__26551\,
            I => \N__26545\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__26548\,
            I => \current_shift_inst.timer_phase.counterZ0Z_13\
        );

    \I__4320\ : Odrv4
    port map (
            O => \N__26545\,
            I => \current_shift_inst.timer_phase.counterZ0Z_13\
        );

    \I__4319\ : InMux
    port map (
            O => \N__26540\,
            I => \current_shift_inst.timer_phase.counter_cry_12\
        );

    \I__4318\ : CascadeMux
    port map (
            O => \N__26537\,
            I => \N__26533\
        );

    \I__4317\ : CascadeMux
    port map (
            O => \N__26536\,
            I => \N__26530\
        );

    \I__4316\ : InMux
    port map (
            O => \N__26533\,
            I => \N__26524\
        );

    \I__4315\ : InMux
    port map (
            O => \N__26530\,
            I => \N__26524\
        );

    \I__4314\ : InMux
    port map (
            O => \N__26529\,
            I => \N__26521\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__26524\,
            I => \N__26518\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__26521\,
            I => \current_shift_inst.timer_phase.counterZ0Z_14\
        );

    \I__4311\ : Odrv12
    port map (
            O => \N__26518\,
            I => \current_shift_inst.timer_phase.counterZ0Z_14\
        );

    \I__4310\ : InMux
    port map (
            O => \N__26513\,
            I => \current_shift_inst.timer_phase.counter_cry_13\
        );

    \I__4309\ : CascadeMux
    port map (
            O => \N__26510\,
            I => \N__26506\
        );

    \I__4308\ : CascadeMux
    port map (
            O => \N__26509\,
            I => \N__26503\
        );

    \I__4307\ : InMux
    port map (
            O => \N__26506\,
            I => \N__26498\
        );

    \I__4306\ : InMux
    port map (
            O => \N__26503\,
            I => \N__26498\
        );

    \I__4305\ : LocalMux
    port map (
            O => \N__26498\,
            I => \N__26494\
        );

    \I__4304\ : InMux
    port map (
            O => \N__26497\,
            I => \N__26491\
        );

    \I__4303\ : Span4Mux_v
    port map (
            O => \N__26494\,
            I => \N__26488\
        );

    \I__4302\ : LocalMux
    port map (
            O => \N__26491\,
            I => \current_shift_inst.timer_phase.counterZ0Z_15\
        );

    \I__4301\ : Odrv4
    port map (
            O => \N__26488\,
            I => \current_shift_inst.timer_phase.counterZ0Z_15\
        );

    \I__4300\ : InMux
    port map (
            O => \N__26483\,
            I => \current_shift_inst.timer_phase.counter_cry_14\
        );

    \I__4299\ : InMux
    port map (
            O => \N__26480\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_29\
        );

    \I__4298\ : CEMux
    port map (
            O => \N__26477\,
            I => \N__26462\
        );

    \I__4297\ : CEMux
    port map (
            O => \N__26476\,
            I => \N__26462\
        );

    \I__4296\ : CEMux
    port map (
            O => \N__26475\,
            I => \N__26462\
        );

    \I__4295\ : CEMux
    port map (
            O => \N__26474\,
            I => \N__26462\
        );

    \I__4294\ : CEMux
    port map (
            O => \N__26473\,
            I => \N__26462\
        );

    \I__4293\ : GlobalMux
    port map (
            O => \N__26462\,
            I => \N__26459\
        );

    \I__4292\ : gio2CtrlBuf
    port map (
            O => \N__26459\,
            I => \current_shift_inst.timer_phase.N_188_i_g\
        );

    \I__4291\ : InMux
    port map (
            O => \N__26456\,
            I => \N__26452\
        );

    \I__4290\ : InMux
    port map (
            O => \N__26455\,
            I => \N__26449\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__26452\,
            I => \N__26446\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__26449\,
            I => \N__26443\
        );

    \I__4287\ : Span12Mux_v
    port map (
            O => \N__26446\,
            I => \N__26439\
        );

    \I__4286\ : Span4Mux_h
    port map (
            O => \N__26443\,
            I => \N__26436\
        );

    \I__4285\ : InMux
    port map (
            O => \N__26442\,
            I => \N__26433\
        );

    \I__4284\ : Odrv12
    port map (
            O => \N__26439\,
            I => \current_shift_inst.timer_phase.counterZ0Z_0\
        );

    \I__4283\ : Odrv4
    port map (
            O => \N__26436\,
            I => \current_shift_inst.timer_phase.counterZ0Z_0\
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__26433\,
            I => \current_shift_inst.timer_phase.counterZ0Z_0\
        );

    \I__4281\ : InMux
    port map (
            O => \N__26426\,
            I => \bfn_9_25_0_\
        );

    \I__4280\ : InMux
    port map (
            O => \N__26423\,
            I => \N__26419\
        );

    \I__4279\ : InMux
    port map (
            O => \N__26422\,
            I => \N__26416\
        );

    \I__4278\ : LocalMux
    port map (
            O => \N__26419\,
            I => \N__26410\
        );

    \I__4277\ : LocalMux
    port map (
            O => \N__26416\,
            I => \N__26410\
        );

    \I__4276\ : InMux
    port map (
            O => \N__26415\,
            I => \N__26407\
        );

    \I__4275\ : Odrv12
    port map (
            O => \N__26410\,
            I => \current_shift_inst.timer_phase.counterZ0Z_1\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__26407\,
            I => \current_shift_inst.timer_phase.counterZ0Z_1\
        );

    \I__4273\ : InMux
    port map (
            O => \N__26402\,
            I => \current_shift_inst.timer_phase.counter_cry_0\
        );

    \I__4272\ : CascadeMux
    port map (
            O => \N__26399\,
            I => \N__26395\
        );

    \I__4271\ : CascadeMux
    port map (
            O => \N__26398\,
            I => \N__26392\
        );

    \I__4270\ : InMux
    port map (
            O => \N__26395\,
            I => \N__26386\
        );

    \I__4269\ : InMux
    port map (
            O => \N__26392\,
            I => \N__26386\
        );

    \I__4268\ : InMux
    port map (
            O => \N__26391\,
            I => \N__26383\
        );

    \I__4267\ : LocalMux
    port map (
            O => \N__26386\,
            I => \N__26380\
        );

    \I__4266\ : LocalMux
    port map (
            O => \N__26383\,
            I => \current_shift_inst.timer_phase.counterZ0Z_2\
        );

    \I__4265\ : Odrv12
    port map (
            O => \N__26380\,
            I => \current_shift_inst.timer_phase.counterZ0Z_2\
        );

    \I__4264\ : InMux
    port map (
            O => \N__26375\,
            I => \current_shift_inst.timer_phase.counter_cry_1\
        );

    \I__4263\ : CascadeMux
    port map (
            O => \N__26372\,
            I => \N__26368\
        );

    \I__4262\ : CascadeMux
    port map (
            O => \N__26371\,
            I => \N__26365\
        );

    \I__4261\ : InMux
    port map (
            O => \N__26368\,
            I => \N__26360\
        );

    \I__4260\ : InMux
    port map (
            O => \N__26365\,
            I => \N__26360\
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__26360\,
            I => \N__26356\
        );

    \I__4258\ : InMux
    port map (
            O => \N__26359\,
            I => \N__26353\
        );

    \I__4257\ : Span4Mux_h
    port map (
            O => \N__26356\,
            I => \N__26350\
        );

    \I__4256\ : LocalMux
    port map (
            O => \N__26353\,
            I => \current_shift_inst.timer_phase.counterZ0Z_3\
        );

    \I__4255\ : Odrv4
    port map (
            O => \N__26350\,
            I => \current_shift_inst.timer_phase.counterZ0Z_3\
        );

    \I__4254\ : InMux
    port map (
            O => \N__26345\,
            I => \current_shift_inst.timer_phase.counter_cry_2\
        );

    \I__4253\ : InMux
    port map (
            O => \N__26342\,
            I => \N__26335\
        );

    \I__4252\ : InMux
    port map (
            O => \N__26341\,
            I => \N__26335\
        );

    \I__4251\ : InMux
    port map (
            O => \N__26340\,
            I => \N__26332\
        );

    \I__4250\ : LocalMux
    port map (
            O => \N__26335\,
            I => \N__26329\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__26332\,
            I => \current_shift_inst.timer_phase.counterZ0Z_4\
        );

    \I__4248\ : Odrv12
    port map (
            O => \N__26329\,
            I => \current_shift_inst.timer_phase.counterZ0Z_4\
        );

    \I__4247\ : InMux
    port map (
            O => \N__26324\,
            I => \current_shift_inst.timer_phase.counter_cry_3\
        );

    \I__4246\ : InMux
    port map (
            O => \N__26321\,
            I => \N__26315\
        );

    \I__4245\ : InMux
    port map (
            O => \N__26320\,
            I => \N__26315\
        );

    \I__4244\ : LocalMux
    port map (
            O => \N__26315\,
            I => \N__26311\
        );

    \I__4243\ : InMux
    port map (
            O => \N__26314\,
            I => \N__26308\
        );

    \I__4242\ : Span4Mux_h
    port map (
            O => \N__26311\,
            I => \N__26305\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__26308\,
            I => \current_shift_inst.timer_phase.counterZ0Z_5\
        );

    \I__4240\ : Odrv4
    port map (
            O => \N__26305\,
            I => \current_shift_inst.timer_phase.counterZ0Z_5\
        );

    \I__4239\ : InMux
    port map (
            O => \N__26300\,
            I => \current_shift_inst.timer_phase.counter_cry_4\
        );

    \I__4238\ : CascadeMux
    port map (
            O => \N__26297\,
            I => \N__26293\
        );

    \I__4237\ : InMux
    port map (
            O => \N__26296\,
            I => \N__26290\
        );

    \I__4236\ : InMux
    port map (
            O => \N__26293\,
            I => \N__26287\
        );

    \I__4235\ : LocalMux
    port map (
            O => \N__26290\,
            I => \N__26283\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__26287\,
            I => \N__26280\
        );

    \I__4233\ : InMux
    port map (
            O => \N__26286\,
            I => \N__26277\
        );

    \I__4232\ : Span4Mux_v
    port map (
            O => \N__26283\,
            I => \N__26272\
        );

    \I__4231\ : Span4Mux_v
    port map (
            O => \N__26280\,
            I => \N__26272\
        );

    \I__4230\ : LocalMux
    port map (
            O => \N__26277\,
            I => \current_shift_inst.timer_phase.counterZ0Z_6\
        );

    \I__4229\ : Odrv4
    port map (
            O => \N__26272\,
            I => \current_shift_inst.timer_phase.counterZ0Z_6\
        );

    \I__4228\ : InMux
    port map (
            O => \N__26267\,
            I => \current_shift_inst.timer_phase.counter_cry_5\
        );

    \I__4227\ : CascadeMux
    port map (
            O => \N__26264\,
            I => \N__26260\
        );

    \I__4226\ : CascadeMux
    port map (
            O => \N__26263\,
            I => \N__26257\
        );

    \I__4225\ : InMux
    port map (
            O => \N__26260\,
            I => \N__26251\
        );

    \I__4224\ : InMux
    port map (
            O => \N__26257\,
            I => \N__26251\
        );

    \I__4223\ : InMux
    port map (
            O => \N__26256\,
            I => \N__26248\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__26251\,
            I => \N__26245\
        );

    \I__4221\ : LocalMux
    port map (
            O => \N__26248\,
            I => \current_shift_inst.timer_phase.counterZ0Z_7\
        );

    \I__4220\ : Odrv12
    port map (
            O => \N__26245\,
            I => \current_shift_inst.timer_phase.counterZ0Z_7\
        );

    \I__4219\ : InMux
    port map (
            O => \N__26240\,
            I => \current_shift_inst.timer_phase.counter_cry_6\
        );

    \I__4218\ : InMux
    port map (
            O => \N__26237\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_20\
        );

    \I__4217\ : InMux
    port map (
            O => \N__26234\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_21\
        );

    \I__4216\ : InMux
    port map (
            O => \N__26231\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_22\
        );

    \I__4215\ : InMux
    port map (
            O => \N__26228\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_23\
        );

    \I__4214\ : InMux
    port map (
            O => \N__26225\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_24\
        );

    \I__4213\ : InMux
    port map (
            O => \N__26222\,
            I => \bfn_9_24_0_\
        );

    \I__4212\ : InMux
    port map (
            O => \N__26219\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_26\
        );

    \I__4211\ : InMux
    port map (
            O => \N__26216\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_27\
        );

    \I__4210\ : InMux
    port map (
            O => \N__26213\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_28\
        );

    \I__4209\ : InMux
    port map (
            O => \N__26210\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_11\
        );

    \I__4208\ : InMux
    port map (
            O => \N__26207\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_12\
        );

    \I__4207\ : InMux
    port map (
            O => \N__26204\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_13\
        );

    \I__4206\ : InMux
    port map (
            O => \N__26201\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_14\
        );

    \I__4205\ : InMux
    port map (
            O => \N__26198\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_15\
        );

    \I__4204\ : InMux
    port map (
            O => \N__26195\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_16\
        );

    \I__4203\ : InMux
    port map (
            O => \N__26192\,
            I => \bfn_9_23_0_\
        );

    \I__4202\ : InMux
    port map (
            O => \N__26189\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_18\
        );

    \I__4201\ : InMux
    port map (
            O => \N__26186\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_19\
        );

    \I__4200\ : InMux
    port map (
            O => \N__26183\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_2\
        );

    \I__4199\ : InMux
    port map (
            O => \N__26180\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_3\
        );

    \I__4198\ : InMux
    port map (
            O => \N__26177\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_4\
        );

    \I__4197\ : InMux
    port map (
            O => \N__26174\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_5\
        );

    \I__4196\ : InMux
    port map (
            O => \N__26171\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_6\
        );

    \I__4195\ : InMux
    port map (
            O => \N__26168\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_7\
        );

    \I__4194\ : InMux
    port map (
            O => \N__26165\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_8\
        );

    \I__4193\ : InMux
    port map (
            O => \N__26162\,
            I => \bfn_9_22_0_\
        );

    \I__4192\ : InMux
    port map (
            O => \N__26159\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_10\
        );

    \I__4191\ : CascadeMux
    port map (
            O => \N__26156\,
            I => \N__26153\
        );

    \I__4190\ : InMux
    port map (
            O => \N__26153\,
            I => \N__26150\
        );

    \I__4189\ : LocalMux
    port map (
            O => \N__26150\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIR32K_22\
        );

    \I__4188\ : InMux
    port map (
            O => \N__26147\,
            I => \N__26144\
        );

    \I__4187\ : LocalMux
    port map (
            O => \N__26144\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPB581_22\
        );

    \I__4186\ : InMux
    port map (
            O => \N__26141\,
            I => \N__26138\
        );

    \I__4185\ : LocalMux
    port map (
            O => \N__26138\,
            I => \N__26135\
        );

    \I__4184\ : Odrv4
    port map (
            O => \N__26135\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJ3381_21\
        );

    \I__4183\ : InMux
    port map (
            O => \N__26132\,
            I => \N__26129\
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__26129\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIVQF91_30\
        );

    \I__4181\ : CascadeMux
    port map (
            O => \N__26126\,
            I => \N__26123\
        );

    \I__4180\ : InMux
    port map (
            O => \N__26123\,
            I => \N__26120\
        );

    \I__4179\ : LocalMux
    port map (
            O => \N__26120\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIAO7K_27\
        );

    \I__4178\ : CascadeMux
    port map (
            O => \N__26117\,
            I => \N__26114\
        );

    \I__4177\ : InMux
    port map (
            O => \N__26114\,
            I => \N__26111\
        );

    \I__4176\ : LocalMux
    port map (
            O => \N__26111\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI4D1J_16\
        );

    \I__4175\ : InMux
    port map (
            O => \N__26108\,
            I => \N__26105\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__26105\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIKKJ81_29\
        );

    \I__4173\ : InMux
    port map (
            O => \N__26102\,
            I => \N__26099\
        );

    \I__4172\ : LocalMux
    port map (
            O => \N__26099\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIHCE81_26\
        );

    \I__4171\ : InMux
    port map (
            O => \N__26096\,
            I => \N__26093\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__26093\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI7DM51_10\
        );

    \I__4169\ : InMux
    port map (
            O => \N__26090\,
            I => \N__26087\
        );

    \I__4168\ : LocalMux
    port map (
            O => \N__26087\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI53NU1_6\
        );

    \I__4167\ : InMux
    port map (
            O => \N__26084\,
            I => \N__26081\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__26081\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI7H2J_17\
        );

    \I__4165\ : CascadeMux
    port map (
            O => \N__26078\,
            I => \N__26075\
        );

    \I__4164\ : InMux
    port map (
            O => \N__26075\,
            I => \N__26072\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__26072\,
            I => \N__26069\
        );

    \I__4162\ : Odrv4
    port map (
            O => \N__26069\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIIKQI_10\
        );

    \I__4161\ : CascadeMux
    port map (
            O => \N__26066\,
            I => \N__26063\
        );

    \I__4160\ : InMux
    port map (
            O => \N__26063\,
            I => \N__26060\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__26060\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIU4VI_14\
        );

    \I__4158\ : InMux
    port map (
            O => \N__26057\,
            I => \N__26054\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__26054\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIBU361_16\
        );

    \I__4156\ : InMux
    port map (
            O => \N__26051\,
            I => \N__26048\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__26048\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIBBPU1_7\
        );

    \I__4154\ : InMux
    port map (
            O => \N__26045\,
            I => \N__26042\
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__26042\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI1PG21_9\
        );

    \I__4152\ : InMux
    port map (
            O => \N__26039\,
            I => \N__26036\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__26036\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINKG81_27\
        );

    \I__4150\ : CascadeMux
    port map (
            O => \N__26033\,
            I => \N__26030\
        );

    \I__4149\ : InMux
    port map (
            O => \N__26030\,
            I => \N__26027\
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__26027\,
            I => \current_shift_inst.un38_control_input_0_cry_2_c_RNOZ0\
        );

    \I__4147\ : CascadeMux
    port map (
            O => \N__26024\,
            I => \N__26021\
        );

    \I__4146\ : InMux
    port map (
            O => \N__26021\,
            I => \N__26018\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__26018\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3\
        );

    \I__4144\ : CascadeMux
    port map (
            O => \N__26015\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3_cascade_\
        );

    \I__4143\ : InMux
    port map (
            O => \N__26012\,
            I => \N__26009\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__26009\,
            I => \current_shift_inst.un38_control_input_0_cry_4_c_RNOZ0\
        );

    \I__4141\ : CascadeMux
    port map (
            O => \N__26006\,
            I => \N__26003\
        );

    \I__4140\ : InMux
    port map (
            O => \N__26003\,
            I => \N__26000\
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__26000\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIK3CV_7\
        );

    \I__4138\ : InMux
    port map (
            O => \N__25997\,
            I => \N__25994\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__25994\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP5T51_13\
        );

    \I__4136\ : CascadeMux
    port map (
            O => \N__25991\,
            I => \N__25988\
        );

    \I__4135\ : InMux
    port map (
            O => \N__25988\,
            I => \N__25985\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__25985\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIER9V_5\
        );

    \I__4133\ : CascadeMux
    port map (
            O => \N__25982\,
            I => \N__25979\
        );

    \I__4132\ : InMux
    port map (
            O => \N__25979\,
            I => \N__25976\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__25976\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJDBL1_10\
        );

    \I__4130\ : InMux
    port map (
            O => \N__25973\,
            I => \N__25970\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__25970\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIE6961_18\
        );

    \I__4128\ : CascadeMux
    port map (
            O => \N__25967\,
            I => \N__25964\
        );

    \I__4127\ : InMux
    port map (
            O => \N__25964\,
            I => \N__25961\
        );

    \I__4126\ : LocalMux
    port map (
            O => \N__25961\,
            I => \N__25958\
        );

    \I__4125\ : Odrv4
    port map (
            O => \N__25958\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIHVAV_6\
        );

    \I__4124\ : InMux
    port map (
            O => \N__25955\,
            I => \N__25951\
        );

    \I__4123\ : InMux
    port map (
            O => \N__25954\,
            I => \N__25947\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__25951\,
            I => \N__25943\
        );

    \I__4121\ : InMux
    port map (
            O => \N__25950\,
            I => \N__25940\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__25947\,
            I => \N__25937\
        );

    \I__4119\ : InMux
    port map (
            O => \N__25946\,
            I => \N__25934\
        );

    \I__4118\ : Span4Mux_h
    port map (
            O => \N__25943\,
            I => \N__25927\
        );

    \I__4117\ : LocalMux
    port map (
            O => \N__25940\,
            I => \N__25927\
        );

    \I__4116\ : Span4Mux_v
    port map (
            O => \N__25937\,
            I => \N__25927\
        );

    \I__4115\ : LocalMux
    port map (
            O => \N__25934\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__4114\ : Odrv4
    port map (
            O => \N__25927\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__4113\ : InMux
    port map (
            O => \N__25922\,
            I => \N__25919\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__25919\,
            I => \N__25916\
        );

    \I__4111\ : Span4Mux_h
    port map (
            O => \N__25916\,
            I => \N__25913\
        );

    \I__4110\ : Odrv4
    port map (
            O => \N__25913\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\
        );

    \I__4109\ : InMux
    port map (
            O => \N__25910\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\
        );

    \I__4108\ : InMux
    port map (
            O => \N__25907\,
            I => \N__25902\
        );

    \I__4107\ : CascadeMux
    port map (
            O => \N__25906\,
            I => \N__25899\
        );

    \I__4106\ : CascadeMux
    port map (
            O => \N__25905\,
            I => \N__25896\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__25902\,
            I => \N__25893\
        );

    \I__4104\ : InMux
    port map (
            O => \N__25899\,
            I => \N__25890\
        );

    \I__4103\ : InMux
    port map (
            O => \N__25896\,
            I => \N__25887\
        );

    \I__4102\ : Span4Mux_v
    port map (
            O => \N__25893\,
            I => \N__25883\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__25890\,
            I => \N__25878\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__25887\,
            I => \N__25878\
        );

    \I__4099\ : InMux
    port map (
            O => \N__25886\,
            I => \N__25875\
        );

    \I__4098\ : Span4Mux_h
    port map (
            O => \N__25883\,
            I => \N__25872\
        );

    \I__4097\ : Odrv12
    port map (
            O => \N__25878\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__4096\ : LocalMux
    port map (
            O => \N__25875\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__4095\ : Odrv4
    port map (
            O => \N__25872\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__4094\ : InMux
    port map (
            O => \N__25865\,
            I => \N__25862\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__25862\,
            I => \N__25859\
        );

    \I__4092\ : Odrv4
    port map (
            O => \N__25859\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\
        );

    \I__4091\ : InMux
    port map (
            O => \N__25856\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\
        );

    \I__4090\ : CascadeMux
    port map (
            O => \N__25853\,
            I => \N__25849\
        );

    \I__4089\ : CascadeMux
    port map (
            O => \N__25852\,
            I => \N__25844\
        );

    \I__4088\ : InMux
    port map (
            O => \N__25849\,
            I => \N__25841\
        );

    \I__4087\ : InMux
    port map (
            O => \N__25848\,
            I => \N__25838\
        );

    \I__4086\ : InMux
    port map (
            O => \N__25847\,
            I => \N__25835\
        );

    \I__4085\ : InMux
    port map (
            O => \N__25844\,
            I => \N__25832\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__25841\,
            I => \N__25829\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__25838\,
            I => \N__25826\
        );

    \I__4082\ : LocalMux
    port map (
            O => \N__25835\,
            I => \N__25823\
        );

    \I__4081\ : LocalMux
    port map (
            O => \N__25832\,
            I => \N__25820\
        );

    \I__4080\ : Span4Mux_h
    port map (
            O => \N__25829\,
            I => \N__25817\
        );

    \I__4079\ : Odrv4
    port map (
            O => \N__25826\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__4078\ : Odrv4
    port map (
            O => \N__25823\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__4077\ : Odrv4
    port map (
            O => \N__25820\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__4076\ : Odrv4
    port map (
            O => \N__25817\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__4075\ : InMux
    port map (
            O => \N__25808\,
            I => \N__25805\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__25805\,
            I => \N__25802\
        );

    \I__4073\ : Odrv4
    port map (
            O => \N__25802\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\
        );

    \I__4072\ : InMux
    port map (
            O => \N__25799\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\
        );

    \I__4071\ : CascadeMux
    port map (
            O => \N__25796\,
            I => \N__25792\
        );

    \I__4070\ : CascadeMux
    port map (
            O => \N__25795\,
            I => \N__25788\
        );

    \I__4069\ : InMux
    port map (
            O => \N__25792\,
            I => \N__25784\
        );

    \I__4068\ : CascadeMux
    port map (
            O => \N__25791\,
            I => \N__25781\
        );

    \I__4067\ : InMux
    port map (
            O => \N__25788\,
            I => \N__25778\
        );

    \I__4066\ : CascadeMux
    port map (
            O => \N__25787\,
            I => \N__25775\
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__25784\,
            I => \N__25772\
        );

    \I__4064\ : InMux
    port map (
            O => \N__25781\,
            I => \N__25769\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__25778\,
            I => \N__25766\
        );

    \I__4062\ : InMux
    port map (
            O => \N__25775\,
            I => \N__25763\
        );

    \I__4061\ : Span4Mux_h
    port map (
            O => \N__25772\,
            I => \N__25760\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__25769\,
            I => \N__25755\
        );

    \I__4059\ : Span4Mux_h
    port map (
            O => \N__25766\,
            I => \N__25755\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__25763\,
            I => \N__25752\
        );

    \I__4057\ : Odrv4
    port map (
            O => \N__25760\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__4056\ : Odrv4
    port map (
            O => \N__25755\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__4055\ : Odrv4
    port map (
            O => \N__25752\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__4054\ : InMux
    port map (
            O => \N__25745\,
            I => \N__25742\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__25742\,
            I => \N__25739\
        );

    \I__4052\ : Odrv12
    port map (
            O => \N__25739\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\
        );

    \I__4051\ : InMux
    port map (
            O => \N__25736\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\
        );

    \I__4050\ : CascadeMux
    port map (
            O => \N__25733\,
            I => \N__25725\
        );

    \I__4049\ : CascadeMux
    port map (
            O => \N__25732\,
            I => \N__25721\
        );

    \I__4048\ : CascadeMux
    port map (
            O => \N__25731\,
            I => \N__25717\
        );

    \I__4047\ : InMux
    port map (
            O => \N__25730\,
            I => \N__25714\
        );

    \I__4046\ : InMux
    port map (
            O => \N__25729\,
            I => \N__25699\
        );

    \I__4045\ : InMux
    port map (
            O => \N__25728\,
            I => \N__25699\
        );

    \I__4044\ : InMux
    port map (
            O => \N__25725\,
            I => \N__25699\
        );

    \I__4043\ : InMux
    port map (
            O => \N__25724\,
            I => \N__25699\
        );

    \I__4042\ : InMux
    port map (
            O => \N__25721\,
            I => \N__25699\
        );

    \I__4041\ : InMux
    port map (
            O => \N__25720\,
            I => \N__25699\
        );

    \I__4040\ : InMux
    port map (
            O => \N__25717\,
            I => \N__25699\
        );

    \I__4039\ : LocalMux
    port map (
            O => \N__25714\,
            I => \N__25696\
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__25699\,
            I => \N__25693\
        );

    \I__4037\ : Span4Mux_h
    port map (
            O => \N__25696\,
            I => \N__25690\
        );

    \I__4036\ : Span4Mux_v
    port map (
            O => \N__25693\,
            I => \N__25687\
        );

    \I__4035\ : Odrv4
    port map (
            O => \N__25690\,
            I => \current_shift_inst.control_inputZ0Z_25\
        );

    \I__4034\ : Odrv4
    port map (
            O => \N__25687\,
            I => \current_shift_inst.control_inputZ0Z_25\
        );

    \I__4033\ : CascadeMux
    port map (
            O => \N__25682\,
            I => \N__25679\
        );

    \I__4032\ : InMux
    port map (
            O => \N__25679\,
            I => \N__25659\
        );

    \I__4031\ : InMux
    port map (
            O => \N__25678\,
            I => \N__25659\
        );

    \I__4030\ : CascadeMux
    port map (
            O => \N__25677\,
            I => \N__25655\
        );

    \I__4029\ : CascadeMux
    port map (
            O => \N__25676\,
            I => \N__25650\
        );

    \I__4028\ : CascadeMux
    port map (
            O => \N__25675\,
            I => \N__25646\
        );

    \I__4027\ : CascadeMux
    port map (
            O => \N__25674\,
            I => \N__25642\
        );

    \I__4026\ : CascadeMux
    port map (
            O => \N__25673\,
            I => \N__25639\
        );

    \I__4025\ : CascadeMux
    port map (
            O => \N__25672\,
            I => \N__25636\
        );

    \I__4024\ : CascadeMux
    port map (
            O => \N__25671\,
            I => \N__25629\
        );

    \I__4023\ : CascadeMux
    port map (
            O => \N__25670\,
            I => \N__25626\
        );

    \I__4022\ : CascadeMux
    port map (
            O => \N__25669\,
            I => \N__25623\
        );

    \I__4021\ : CascadeMux
    port map (
            O => \N__25668\,
            I => \N__25620\
        );

    \I__4020\ : CascadeMux
    port map (
            O => \N__25667\,
            I => \N__25615\
        );

    \I__4019\ : CascadeMux
    port map (
            O => \N__25666\,
            I => \N__25610\
        );

    \I__4018\ : CascadeMux
    port map (
            O => \N__25665\,
            I => \N__25607\
        );

    \I__4017\ : CascadeMux
    port map (
            O => \N__25664\,
            I => \N__25604\
        );

    \I__4016\ : LocalMux
    port map (
            O => \N__25659\,
            I => \N__25598\
        );

    \I__4015\ : InMux
    port map (
            O => \N__25658\,
            I => \N__25595\
        );

    \I__4014\ : InMux
    port map (
            O => \N__25655\,
            I => \N__25590\
        );

    \I__4013\ : InMux
    port map (
            O => \N__25654\,
            I => \N__25590\
        );

    \I__4012\ : InMux
    port map (
            O => \N__25653\,
            I => \N__25587\
        );

    \I__4011\ : InMux
    port map (
            O => \N__25650\,
            I => \N__25582\
        );

    \I__4010\ : InMux
    port map (
            O => \N__25649\,
            I => \N__25582\
        );

    \I__4009\ : InMux
    port map (
            O => \N__25646\,
            I => \N__25579\
        );

    \I__4008\ : InMux
    port map (
            O => \N__25645\,
            I => \N__25564\
        );

    \I__4007\ : InMux
    port map (
            O => \N__25642\,
            I => \N__25564\
        );

    \I__4006\ : InMux
    port map (
            O => \N__25639\,
            I => \N__25564\
        );

    \I__4005\ : InMux
    port map (
            O => \N__25636\,
            I => \N__25564\
        );

    \I__4004\ : InMux
    port map (
            O => \N__25635\,
            I => \N__25564\
        );

    \I__4003\ : InMux
    port map (
            O => \N__25634\,
            I => \N__25564\
        );

    \I__4002\ : InMux
    port map (
            O => \N__25633\,
            I => \N__25564\
        );

    \I__4001\ : InMux
    port map (
            O => \N__25632\,
            I => \N__25561\
        );

    \I__4000\ : InMux
    port map (
            O => \N__25629\,
            I => \N__25548\
        );

    \I__3999\ : InMux
    port map (
            O => \N__25626\,
            I => \N__25548\
        );

    \I__3998\ : InMux
    port map (
            O => \N__25623\,
            I => \N__25548\
        );

    \I__3997\ : InMux
    port map (
            O => \N__25620\,
            I => \N__25548\
        );

    \I__3996\ : InMux
    port map (
            O => \N__25619\,
            I => \N__25548\
        );

    \I__3995\ : InMux
    port map (
            O => \N__25618\,
            I => \N__25548\
        );

    \I__3994\ : InMux
    port map (
            O => \N__25615\,
            I => \N__25543\
        );

    \I__3993\ : InMux
    port map (
            O => \N__25614\,
            I => \N__25543\
        );

    \I__3992\ : InMux
    port map (
            O => \N__25613\,
            I => \N__25528\
        );

    \I__3991\ : InMux
    port map (
            O => \N__25610\,
            I => \N__25528\
        );

    \I__3990\ : InMux
    port map (
            O => \N__25607\,
            I => \N__25528\
        );

    \I__3989\ : InMux
    port map (
            O => \N__25604\,
            I => \N__25528\
        );

    \I__3988\ : InMux
    port map (
            O => \N__25603\,
            I => \N__25528\
        );

    \I__3987\ : InMux
    port map (
            O => \N__25602\,
            I => \N__25528\
        );

    \I__3986\ : InMux
    port map (
            O => \N__25601\,
            I => \N__25528\
        );

    \I__3985\ : Span4Mux_v
    port map (
            O => \N__25598\,
            I => \N__25525\
        );

    \I__3984\ : LocalMux
    port map (
            O => \N__25595\,
            I => \N__25518\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__25590\,
            I => \N__25518\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__25587\,
            I => \N__25518\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__25582\,
            I => \N__25513\
        );

    \I__3980\ : LocalMux
    port map (
            O => \N__25579\,
            I => \N__25513\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__25564\,
            I => \N__25508\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__25561\,
            I => \N__25508\
        );

    \I__3977\ : LocalMux
    port map (
            O => \N__25548\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3976\ : LocalMux
    port map (
            O => \N__25543\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__25528\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3974\ : Odrv4
    port map (
            O => \N__25525\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3973\ : Odrv12
    port map (
            O => \N__25518\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3972\ : Odrv12
    port map (
            O => \N__25513\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3971\ : Odrv4
    port map (
            O => \N__25508\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3970\ : InMux
    port map (
            O => \N__25493\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_30\
        );

    \I__3969\ : InMux
    port map (
            O => \N__25490\,
            I => \N__25487\
        );

    \I__3968\ : LocalMux
    port map (
            O => \N__25487\,
            I => \N__25484\
        );

    \I__3967\ : Odrv4
    port map (
            O => \N__25484\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\
        );

    \I__3966\ : InMux
    port map (
            O => \N__25481\,
            I => \N__25478\
        );

    \I__3965\ : LocalMux
    port map (
            O => \N__25478\,
            I => \current_shift_inst.un38_control_input_0_cry_1_c_RNOZ0\
        );

    \I__3964\ : InMux
    port map (
            O => \N__25475\,
            I => \N__25472\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__25472\,
            I => \current_shift_inst.N_1717_i\
        );

    \I__3962\ : CascadeMux
    port map (
            O => \N__25469\,
            I => \N__25466\
        );

    \I__3961\ : InMux
    port map (
            O => \N__25466\,
            I => \N__25463\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__25463\,
            I => \N__25457\
        );

    \I__3959\ : InMux
    port map (
            O => \N__25462\,
            I => \N__25454\
        );

    \I__3958\ : InMux
    port map (
            O => \N__25461\,
            I => \N__25449\
        );

    \I__3957\ : InMux
    port map (
            O => \N__25460\,
            I => \N__25449\
        );

    \I__3956\ : Odrv12
    port map (
            O => \N__25457\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__25454\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__3954\ : LocalMux
    port map (
            O => \N__25449\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__3953\ : InMux
    port map (
            O => \N__25442\,
            I => \N__25438\
        );

    \I__3952\ : CascadeMux
    port map (
            O => \N__25441\,
            I => \N__25435\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__25438\,
            I => \N__25432\
        );

    \I__3950\ : InMux
    port map (
            O => \N__25435\,
            I => \N__25429\
        );

    \I__3949\ : Span4Mux_h
    port map (
            O => \N__25432\,
            I => \N__25426\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__25429\,
            I => \N__25423\
        );

    \I__3947\ : Span4Mux_v
    port map (
            O => \N__25426\,
            I => \N__25420\
        );

    \I__3946\ : Span4Mux_h
    port map (
            O => \N__25423\,
            I => \N__25417\
        );

    \I__3945\ : Odrv4
    port map (
            O => \N__25420\,
            I => \current_shift_inst.control_inputZ0Z_20\
        );

    \I__3944\ : Odrv4
    port map (
            O => \N__25417\,
            I => \current_shift_inst.control_inputZ0Z_20\
        );

    \I__3943\ : InMux
    port map (
            O => \N__25412\,
            I => \N__25409\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__25409\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\
        );

    \I__3941\ : InMux
    port map (
            O => \N__25406\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\
        );

    \I__3940\ : CascadeMux
    port map (
            O => \N__25403\,
            I => \N__25400\
        );

    \I__3939\ : InMux
    port map (
            O => \N__25400\,
            I => \N__25397\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__25397\,
            I => \N__25393\
        );

    \I__3937\ : InMux
    port map (
            O => \N__25396\,
            I => \N__25390\
        );

    \I__3936\ : Span4Mux_v
    port map (
            O => \N__25393\,
            I => \N__25387\
        );

    \I__3935\ : LocalMux
    port map (
            O => \N__25390\,
            I => \N__25382\
        );

    \I__3934\ : Span4Mux_h
    port map (
            O => \N__25387\,
            I => \N__25379\
        );

    \I__3933\ : InMux
    port map (
            O => \N__25386\,
            I => \N__25376\
        );

    \I__3932\ : InMux
    port map (
            O => \N__25385\,
            I => \N__25373\
        );

    \I__3931\ : Span4Mux_v
    port map (
            O => \N__25382\,
            I => \N__25370\
        );

    \I__3930\ : Odrv4
    port map (
            O => \N__25379\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__25376\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__25373\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__3927\ : Odrv4
    port map (
            O => \N__25370\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__3926\ : InMux
    port map (
            O => \N__25361\,
            I => \N__25357\
        );

    \I__3925\ : CascadeMux
    port map (
            O => \N__25360\,
            I => \N__25354\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__25357\,
            I => \N__25351\
        );

    \I__3923\ : InMux
    port map (
            O => \N__25354\,
            I => \N__25348\
        );

    \I__3922\ : Span4Mux_v
    port map (
            O => \N__25351\,
            I => \N__25345\
        );

    \I__3921\ : LocalMux
    port map (
            O => \N__25348\,
            I => \N__25342\
        );

    \I__3920\ : Sp12to4
    port map (
            O => \N__25345\,
            I => \N__25339\
        );

    \I__3919\ : Span4Mux_h
    port map (
            O => \N__25342\,
            I => \N__25336\
        );

    \I__3918\ : Odrv12
    port map (
            O => \N__25339\,
            I => \current_shift_inst.control_inputZ0Z_21\
        );

    \I__3917\ : Odrv4
    port map (
            O => \N__25336\,
            I => \current_shift_inst.control_inputZ0Z_21\
        );

    \I__3916\ : InMux
    port map (
            O => \N__25331\,
            I => \N__25328\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__25328\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\
        );

    \I__3914\ : InMux
    port map (
            O => \N__25325\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\
        );

    \I__3913\ : InMux
    port map (
            O => \N__25322\,
            I => \N__25317\
        );

    \I__3912\ : CascadeMux
    port map (
            O => \N__25321\,
            I => \N__25313\
        );

    \I__3911\ : CascadeMux
    port map (
            O => \N__25320\,
            I => \N__25310\
        );

    \I__3910\ : LocalMux
    port map (
            O => \N__25317\,
            I => \N__25307\
        );

    \I__3909\ : InMux
    port map (
            O => \N__25316\,
            I => \N__25304\
        );

    \I__3908\ : InMux
    port map (
            O => \N__25313\,
            I => \N__25299\
        );

    \I__3907\ : InMux
    port map (
            O => \N__25310\,
            I => \N__25299\
        );

    \I__3906\ : Odrv12
    port map (
            O => \N__25307\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__25304\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__3904\ : LocalMux
    port map (
            O => \N__25299\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__3903\ : CascadeMux
    port map (
            O => \N__25292\,
            I => \N__25289\
        );

    \I__3902\ : InMux
    port map (
            O => \N__25289\,
            I => \N__25285\
        );

    \I__3901\ : InMux
    port map (
            O => \N__25288\,
            I => \N__25282\
        );

    \I__3900\ : LocalMux
    port map (
            O => \N__25285\,
            I => \N__25279\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__25282\,
            I => \N__25274\
        );

    \I__3898\ : Span4Mux_h
    port map (
            O => \N__25279\,
            I => \N__25274\
        );

    \I__3897\ : Span4Mux_v
    port map (
            O => \N__25274\,
            I => \N__25271\
        );

    \I__3896\ : Odrv4
    port map (
            O => \N__25271\,
            I => \current_shift_inst.control_inputZ0Z_22\
        );

    \I__3895\ : InMux
    port map (
            O => \N__25268\,
            I => \N__25265\
        );

    \I__3894\ : LocalMux
    port map (
            O => \N__25265\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\
        );

    \I__3893\ : InMux
    port map (
            O => \N__25262\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\
        );

    \I__3892\ : InMux
    port map (
            O => \N__25259\,
            I => \N__25254\
        );

    \I__3891\ : InMux
    port map (
            O => \N__25258\,
            I => \N__25251\
        );

    \I__3890\ : InMux
    port map (
            O => \N__25257\,
            I => \N__25247\
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__25254\,
            I => \N__25244\
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__25251\,
            I => \N__25241\
        );

    \I__3887\ : InMux
    port map (
            O => \N__25250\,
            I => \N__25238\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__25247\,
            I => \N__25235\
        );

    \I__3885\ : Odrv12
    port map (
            O => \N__25244\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__3884\ : Odrv4
    port map (
            O => \N__25241\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__25238\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__3882\ : Odrv4
    port map (
            O => \N__25235\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__3881\ : CascadeMux
    port map (
            O => \N__25226\,
            I => \N__25223\
        );

    \I__3880\ : InMux
    port map (
            O => \N__25223\,
            I => \N__25219\
        );

    \I__3879\ : InMux
    port map (
            O => \N__25222\,
            I => \N__25216\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__25219\,
            I => \N__25213\
        );

    \I__3877\ : LocalMux
    port map (
            O => \N__25216\,
            I => \N__25208\
        );

    \I__3876\ : Span4Mux_h
    port map (
            O => \N__25213\,
            I => \N__25208\
        );

    \I__3875\ : Span4Mux_v
    port map (
            O => \N__25208\,
            I => \N__25205\
        );

    \I__3874\ : Odrv4
    port map (
            O => \N__25205\,
            I => \current_shift_inst.control_inputZ0Z_23\
        );

    \I__3873\ : CascadeMux
    port map (
            O => \N__25202\,
            I => \N__25199\
        );

    \I__3872\ : InMux
    port map (
            O => \N__25199\,
            I => \N__25196\
        );

    \I__3871\ : LocalMux
    port map (
            O => \N__25196\,
            I => \N__25193\
        );

    \I__3870\ : Span4Mux_h
    port map (
            O => \N__25193\,
            I => \N__25190\
        );

    \I__3869\ : Odrv4
    port map (
            O => \N__25190\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\
        );

    \I__3868\ : InMux
    port map (
            O => \N__25187\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\
        );

    \I__3867\ : CascadeMux
    port map (
            O => \N__25184\,
            I => \N__25181\
        );

    \I__3866\ : InMux
    port map (
            O => \N__25181\,
            I => \N__25177\
        );

    \I__3865\ : InMux
    port map (
            O => \N__25180\,
            I => \N__25173\
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__25177\,
            I => \N__25170\
        );

    \I__3863\ : InMux
    port map (
            O => \N__25176\,
            I => \N__25167\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__25173\,
            I => \N__25163\
        );

    \I__3861\ : Span4Mux_h
    port map (
            O => \N__25170\,
            I => \N__25158\
        );

    \I__3860\ : LocalMux
    port map (
            O => \N__25167\,
            I => \N__25158\
        );

    \I__3859\ : InMux
    port map (
            O => \N__25166\,
            I => \N__25155\
        );

    \I__3858\ : Span4Mux_h
    port map (
            O => \N__25163\,
            I => \N__25152\
        );

    \I__3857\ : Odrv4
    port map (
            O => \N__25158\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__25155\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__3855\ : Odrv4
    port map (
            O => \N__25152\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__3854\ : CascadeMux
    port map (
            O => \N__25145\,
            I => \N__25141\
        );

    \I__3853\ : InMux
    port map (
            O => \N__25144\,
            I => \N__25138\
        );

    \I__3852\ : InMux
    port map (
            O => \N__25141\,
            I => \N__25135\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__25138\,
            I => \N__25132\
        );

    \I__3850\ : LocalMux
    port map (
            O => \N__25135\,
            I => \N__25129\
        );

    \I__3849\ : Span4Mux_h
    port map (
            O => \N__25132\,
            I => \N__25126\
        );

    \I__3848\ : Span4Mux_h
    port map (
            O => \N__25129\,
            I => \N__25123\
        );

    \I__3847\ : Odrv4
    port map (
            O => \N__25126\,
            I => \current_shift_inst.control_inputZ0Z_24\
        );

    \I__3846\ : Odrv4
    port map (
            O => \N__25123\,
            I => \current_shift_inst.control_inputZ0Z_24\
        );

    \I__3845\ : InMux
    port map (
            O => \N__25118\,
            I => \N__25115\
        );

    \I__3844\ : LocalMux
    port map (
            O => \N__25115\,
            I => \N__25112\
        );

    \I__3843\ : Odrv12
    port map (
            O => \N__25112\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\
        );

    \I__3842\ : InMux
    port map (
            O => \N__25109\,
            I => \bfn_9_16_0_\
        );

    \I__3841\ : InMux
    port map (
            O => \N__25106\,
            I => \N__25102\
        );

    \I__3840\ : InMux
    port map (
            O => \N__25105\,
            I => \N__25098\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__25102\,
            I => \N__25095\
        );

    \I__3838\ : InMux
    port map (
            O => \N__25101\,
            I => \N__25092\
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__25098\,
            I => \N__25088\
        );

    \I__3836\ : Span4Mux_h
    port map (
            O => \N__25095\,
            I => \N__25083\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__25092\,
            I => \N__25083\
        );

    \I__3834\ : InMux
    port map (
            O => \N__25091\,
            I => \N__25080\
        );

    \I__3833\ : Span4Mux_h
    port map (
            O => \N__25088\,
            I => \N__25077\
        );

    \I__3832\ : Odrv4
    port map (
            O => \N__25083\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__3831\ : LocalMux
    port map (
            O => \N__25080\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__3830\ : Odrv4
    port map (
            O => \N__25077\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__3829\ : InMux
    port map (
            O => \N__25070\,
            I => \N__25067\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__25067\,
            I => \N__25064\
        );

    \I__3827\ : Span4Mux_h
    port map (
            O => \N__25064\,
            I => \N__25061\
        );

    \I__3826\ : Odrv4
    port map (
            O => \N__25061\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\
        );

    \I__3825\ : InMux
    port map (
            O => \N__25058\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\
        );

    \I__3824\ : CascadeMux
    port map (
            O => \N__25055\,
            I => \N__25051\
        );

    \I__3823\ : CascadeMux
    port map (
            O => \N__25054\,
            I => \N__25047\
        );

    \I__3822\ : InMux
    port map (
            O => \N__25051\,
            I => \N__25044\
        );

    \I__3821\ : CascadeMux
    port map (
            O => \N__25050\,
            I => \N__25041\
        );

    \I__3820\ : InMux
    port map (
            O => \N__25047\,
            I => \N__25037\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__25044\,
            I => \N__25034\
        );

    \I__3818\ : InMux
    port map (
            O => \N__25041\,
            I => \N__25031\
        );

    \I__3817\ : CascadeMux
    port map (
            O => \N__25040\,
            I => \N__25028\
        );

    \I__3816\ : LocalMux
    port map (
            O => \N__25037\,
            I => \N__25025\
        );

    \I__3815\ : Span4Mux_h
    port map (
            O => \N__25034\,
            I => \N__25020\
        );

    \I__3814\ : LocalMux
    port map (
            O => \N__25031\,
            I => \N__25020\
        );

    \I__3813\ : InMux
    port map (
            O => \N__25028\,
            I => \N__25017\
        );

    \I__3812\ : Span4Mux_h
    port map (
            O => \N__25025\,
            I => \N__25014\
        );

    \I__3811\ : Odrv4
    port map (
            O => \N__25020\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__25017\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__3809\ : Odrv4
    port map (
            O => \N__25014\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__3808\ : InMux
    port map (
            O => \N__25007\,
            I => \N__25004\
        );

    \I__3807\ : LocalMux
    port map (
            O => \N__25004\,
            I => \N__25001\
        );

    \I__3806\ : Span4Mux_h
    port map (
            O => \N__25001\,
            I => \N__24998\
        );

    \I__3805\ : Odrv4
    port map (
            O => \N__24998\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\
        );

    \I__3804\ : InMux
    port map (
            O => \N__24995\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\
        );

    \I__3803\ : InMux
    port map (
            O => \N__24992\,
            I => \N__24989\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__24989\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\
        );

    \I__3801\ : InMux
    port map (
            O => \N__24986\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\
        );

    \I__3800\ : CascadeMux
    port map (
            O => \N__24983\,
            I => \N__24979\
        );

    \I__3799\ : InMux
    port map (
            O => \N__24982\,
            I => \N__24976\
        );

    \I__3798\ : InMux
    port map (
            O => \N__24979\,
            I => \N__24973\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__24976\,
            I => \N__24968\
        );

    \I__3796\ : LocalMux
    port map (
            O => \N__24973\,
            I => \N__24965\
        );

    \I__3795\ : InMux
    port map (
            O => \N__24972\,
            I => \N__24962\
        );

    \I__3794\ : InMux
    port map (
            O => \N__24971\,
            I => \N__24959\
        );

    \I__3793\ : Span4Mux_h
    port map (
            O => \N__24968\,
            I => \N__24956\
        );

    \I__3792\ : Odrv12
    port map (
            O => \N__24965\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__24962\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__24959\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__3789\ : Odrv4
    port map (
            O => \N__24956\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__3788\ : CascadeMux
    port map (
            O => \N__24947\,
            I => \N__24943\
        );

    \I__3787\ : InMux
    port map (
            O => \N__24946\,
            I => \N__24940\
        );

    \I__3786\ : InMux
    port map (
            O => \N__24943\,
            I => \N__24937\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__24940\,
            I => \N__24934\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__24937\,
            I => \N__24931\
        );

    \I__3783\ : Span4Mux_h
    port map (
            O => \N__24934\,
            I => \N__24926\
        );

    \I__3782\ : Span4Mux_h
    port map (
            O => \N__24931\,
            I => \N__24926\
        );

    \I__3781\ : Odrv4
    port map (
            O => \N__24926\,
            I => \current_shift_inst.control_inputZ0Z_13\
        );

    \I__3780\ : InMux
    port map (
            O => \N__24923\,
            I => \N__24920\
        );

    \I__3779\ : LocalMux
    port map (
            O => \N__24920\,
            I => \N__24917\
        );

    \I__3778\ : Odrv4
    port map (
            O => \N__24917\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\
        );

    \I__3777\ : InMux
    port map (
            O => \N__24914\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\
        );

    \I__3776\ : InMux
    port map (
            O => \N__24911\,
            I => \N__24907\
        );

    \I__3775\ : InMux
    port map (
            O => \N__24910\,
            I => \N__24904\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__24907\,
            I => \N__24901\
        );

    \I__3773\ : LocalMux
    port map (
            O => \N__24904\,
            I => \N__24898\
        );

    \I__3772\ : Span12Mux_v
    port map (
            O => \N__24901\,
            I => \N__24895\
        );

    \I__3771\ : Span12Mux_v
    port map (
            O => \N__24898\,
            I => \N__24892\
        );

    \I__3770\ : Odrv12
    port map (
            O => \N__24895\,
            I => \current_shift_inst.control_inputZ0Z_14\
        );

    \I__3769\ : Odrv12
    port map (
            O => \N__24892\,
            I => \current_shift_inst.control_inputZ0Z_14\
        );

    \I__3768\ : CascadeMux
    port map (
            O => \N__24887\,
            I => \N__24884\
        );

    \I__3767\ : InMux
    port map (
            O => \N__24884\,
            I => \N__24881\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__24881\,
            I => \N__24876\
        );

    \I__3765\ : InMux
    port map (
            O => \N__24880\,
            I => \N__24872\
        );

    \I__3764\ : CascadeMux
    port map (
            O => \N__24879\,
            I => \N__24869\
        );

    \I__3763\ : Span4Mux_v
    port map (
            O => \N__24876\,
            I => \N__24866\
        );

    \I__3762\ : InMux
    port map (
            O => \N__24875\,
            I => \N__24863\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__24872\,
            I => \N__24860\
        );

    \I__3760\ : InMux
    port map (
            O => \N__24869\,
            I => \N__24857\
        );

    \I__3759\ : Span4Mux_h
    port map (
            O => \N__24866\,
            I => \N__24852\
        );

    \I__3758\ : LocalMux
    port map (
            O => \N__24863\,
            I => \N__24852\
        );

    \I__3757\ : Odrv4
    port map (
            O => \N__24860\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__24857\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__3755\ : Odrv4
    port map (
            O => \N__24852\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__3754\ : InMux
    port map (
            O => \N__24845\,
            I => \N__24842\
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__24842\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\
        );

    \I__3752\ : InMux
    port map (
            O => \N__24839\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\
        );

    \I__3751\ : CascadeMux
    port map (
            O => \N__24836\,
            I => \N__24833\
        );

    \I__3750\ : InMux
    port map (
            O => \N__24833\,
            I => \N__24829\
        );

    \I__3749\ : InMux
    port map (
            O => \N__24832\,
            I => \N__24826\
        );

    \I__3748\ : LocalMux
    port map (
            O => \N__24829\,
            I => \N__24822\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__24826\,
            I => \N__24818\
        );

    \I__3746\ : InMux
    port map (
            O => \N__24825\,
            I => \N__24815\
        );

    \I__3745\ : Span4Mux_h
    port map (
            O => \N__24822\,
            I => \N__24812\
        );

    \I__3744\ : InMux
    port map (
            O => \N__24821\,
            I => \N__24809\
        );

    \I__3743\ : Span4Mux_v
    port map (
            O => \N__24818\,
            I => \N__24804\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__24815\,
            I => \N__24804\
        );

    \I__3741\ : Odrv4
    port map (
            O => \N__24812\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__24809\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__3739\ : Odrv4
    port map (
            O => \N__24804\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__3738\ : InMux
    port map (
            O => \N__24797\,
            I => \N__24793\
        );

    \I__3737\ : CascadeMux
    port map (
            O => \N__24796\,
            I => \N__24790\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__24793\,
            I => \N__24787\
        );

    \I__3735\ : InMux
    port map (
            O => \N__24790\,
            I => \N__24784\
        );

    \I__3734\ : Span4Mux_h
    port map (
            O => \N__24787\,
            I => \N__24779\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__24784\,
            I => \N__24779\
        );

    \I__3732\ : Span4Mux_h
    port map (
            O => \N__24779\,
            I => \N__24776\
        );

    \I__3731\ : Span4Mux_v
    port map (
            O => \N__24776\,
            I => \N__24773\
        );

    \I__3730\ : Odrv4
    port map (
            O => \N__24773\,
            I => \current_shift_inst.control_inputZ0Z_15\
        );

    \I__3729\ : InMux
    port map (
            O => \N__24770\,
            I => \N__24767\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__24767\,
            I => \N__24764\
        );

    \I__3727\ : Span4Mux_h
    port map (
            O => \N__24764\,
            I => \N__24761\
        );

    \I__3726\ : Odrv4
    port map (
            O => \N__24761\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\
        );

    \I__3725\ : InMux
    port map (
            O => \N__24758\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\
        );

    \I__3724\ : CascadeMux
    port map (
            O => \N__24755\,
            I => \N__24750\
        );

    \I__3723\ : InMux
    port map (
            O => \N__24754\,
            I => \N__24747\
        );

    \I__3722\ : CascadeMux
    port map (
            O => \N__24753\,
            I => \N__24743\
        );

    \I__3721\ : InMux
    port map (
            O => \N__24750\,
            I => \N__24740\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__24747\,
            I => \N__24737\
        );

    \I__3719\ : InMux
    port map (
            O => \N__24746\,
            I => \N__24734\
        );

    \I__3718\ : InMux
    port map (
            O => \N__24743\,
            I => \N__24731\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__24740\,
            I => \N__24728\
        );

    \I__3716\ : Odrv12
    port map (
            O => \N__24737\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__24734\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__24731\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__3713\ : Odrv4
    port map (
            O => \N__24728\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__3712\ : CascadeMux
    port map (
            O => \N__24719\,
            I => \N__24715\
        );

    \I__3711\ : InMux
    port map (
            O => \N__24718\,
            I => \N__24712\
        );

    \I__3710\ : InMux
    port map (
            O => \N__24715\,
            I => \N__24709\
        );

    \I__3709\ : LocalMux
    port map (
            O => \N__24712\,
            I => \N__24706\
        );

    \I__3708\ : LocalMux
    port map (
            O => \N__24709\,
            I => \N__24703\
        );

    \I__3707\ : Span4Mux_h
    port map (
            O => \N__24706\,
            I => \N__24700\
        );

    \I__3706\ : Span4Mux_h
    port map (
            O => \N__24703\,
            I => \N__24697\
        );

    \I__3705\ : Odrv4
    port map (
            O => \N__24700\,
            I => \current_shift_inst.control_inputZ0Z_16\
        );

    \I__3704\ : Odrv4
    port map (
            O => \N__24697\,
            I => \current_shift_inst.control_inputZ0Z_16\
        );

    \I__3703\ : InMux
    port map (
            O => \N__24692\,
            I => \N__24689\
        );

    \I__3702\ : LocalMux
    port map (
            O => \N__24689\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\
        );

    \I__3701\ : InMux
    port map (
            O => \N__24686\,
            I => \bfn_9_15_0_\
        );

    \I__3700\ : InMux
    port map (
            O => \N__24683\,
            I => \N__24680\
        );

    \I__3699\ : LocalMux
    port map (
            O => \N__24680\,
            I => \N__24674\
        );

    \I__3698\ : InMux
    port map (
            O => \N__24679\,
            I => \N__24671\
        );

    \I__3697\ : InMux
    port map (
            O => \N__24678\,
            I => \N__24666\
        );

    \I__3696\ : InMux
    port map (
            O => \N__24677\,
            I => \N__24666\
        );

    \I__3695\ : Odrv12
    port map (
            O => \N__24674\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__3694\ : LocalMux
    port map (
            O => \N__24671\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__24666\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__3692\ : InMux
    port map (
            O => \N__24659\,
            I => \N__24655\
        );

    \I__3691\ : CascadeMux
    port map (
            O => \N__24658\,
            I => \N__24652\
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__24655\,
            I => \N__24649\
        );

    \I__3689\ : InMux
    port map (
            O => \N__24652\,
            I => \N__24646\
        );

    \I__3688\ : Span4Mux_h
    port map (
            O => \N__24649\,
            I => \N__24643\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__24646\,
            I => \N__24640\
        );

    \I__3686\ : Span4Mux_v
    port map (
            O => \N__24643\,
            I => \N__24637\
        );

    \I__3685\ : Span4Mux_h
    port map (
            O => \N__24640\,
            I => \N__24634\
        );

    \I__3684\ : Odrv4
    port map (
            O => \N__24637\,
            I => \current_shift_inst.control_inputZ0Z_17\
        );

    \I__3683\ : Odrv4
    port map (
            O => \N__24634\,
            I => \current_shift_inst.control_inputZ0Z_17\
        );

    \I__3682\ : InMux
    port map (
            O => \N__24629\,
            I => \N__24626\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__24626\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\
        );

    \I__3680\ : InMux
    port map (
            O => \N__24623\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\
        );

    \I__3679\ : CascadeMux
    port map (
            O => \N__24620\,
            I => \N__24617\
        );

    \I__3678\ : InMux
    port map (
            O => \N__24617\,
            I => \N__24614\
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__24614\,
            I => \N__24607\
        );

    \I__3676\ : InMux
    port map (
            O => \N__24613\,
            I => \N__24600\
        );

    \I__3675\ : InMux
    port map (
            O => \N__24612\,
            I => \N__24600\
        );

    \I__3674\ : InMux
    port map (
            O => \N__24611\,
            I => \N__24600\
        );

    \I__3673\ : InMux
    port map (
            O => \N__24610\,
            I => \N__24596\
        );

    \I__3672\ : Span4Mux_h
    port map (
            O => \N__24607\,
            I => \N__24593\
        );

    \I__3671\ : LocalMux
    port map (
            O => \N__24600\,
            I => \N__24590\
        );

    \I__3670\ : InMux
    port map (
            O => \N__24599\,
            I => \N__24587\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__24596\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__3668\ : Odrv4
    port map (
            O => \N__24593\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__3667\ : Odrv4
    port map (
            O => \N__24590\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__3666\ : LocalMux
    port map (
            O => \N__24587\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__3665\ : CascadeMux
    port map (
            O => \N__24578\,
            I => \N__24574\
        );

    \I__3664\ : InMux
    port map (
            O => \N__24577\,
            I => \N__24571\
        );

    \I__3663\ : InMux
    port map (
            O => \N__24574\,
            I => \N__24568\
        );

    \I__3662\ : LocalMux
    port map (
            O => \N__24571\,
            I => \N__24565\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__24568\,
            I => \N__24562\
        );

    \I__3660\ : Span4Mux_h
    port map (
            O => \N__24565\,
            I => \N__24559\
        );

    \I__3659\ : Span4Mux_h
    port map (
            O => \N__24562\,
            I => \N__24556\
        );

    \I__3658\ : Odrv4
    port map (
            O => \N__24559\,
            I => \current_shift_inst.control_inputZ0Z_18\
        );

    \I__3657\ : Odrv4
    port map (
            O => \N__24556\,
            I => \current_shift_inst.control_inputZ0Z_18\
        );

    \I__3656\ : InMux
    port map (
            O => \N__24551\,
            I => \N__24548\
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__24548\,
            I => \N__24545\
        );

    \I__3654\ : Odrv4
    port map (
            O => \N__24545\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\
        );

    \I__3653\ : InMux
    port map (
            O => \N__24542\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\
        );

    \I__3652\ : InMux
    port map (
            O => \N__24539\,
            I => \N__24536\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__24536\,
            I => \N__24530\
        );

    \I__3650\ : InMux
    port map (
            O => \N__24535\,
            I => \N__24527\
        );

    \I__3649\ : InMux
    port map (
            O => \N__24534\,
            I => \N__24522\
        );

    \I__3648\ : InMux
    port map (
            O => \N__24533\,
            I => \N__24522\
        );

    \I__3647\ : Odrv12
    port map (
            O => \N__24530\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__24527\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__24522\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__3644\ : InMux
    port map (
            O => \N__24515\,
            I => \N__24511\
        );

    \I__3643\ : CascadeMux
    port map (
            O => \N__24514\,
            I => \N__24508\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__24511\,
            I => \N__24505\
        );

    \I__3641\ : InMux
    port map (
            O => \N__24508\,
            I => \N__24502\
        );

    \I__3640\ : Span4Mux_h
    port map (
            O => \N__24505\,
            I => \N__24499\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__24502\,
            I => \N__24496\
        );

    \I__3638\ : Span4Mux_v
    port map (
            O => \N__24499\,
            I => \N__24493\
        );

    \I__3637\ : Span4Mux_h
    port map (
            O => \N__24496\,
            I => \N__24490\
        );

    \I__3636\ : Odrv4
    port map (
            O => \N__24493\,
            I => \current_shift_inst.control_inputZ0Z_19\
        );

    \I__3635\ : Odrv4
    port map (
            O => \N__24490\,
            I => \current_shift_inst.control_inputZ0Z_19\
        );

    \I__3634\ : InMux
    port map (
            O => \N__24485\,
            I => \N__24482\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__24482\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\
        );

    \I__3632\ : InMux
    port map (
            O => \N__24479\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\
        );

    \I__3631\ : InMux
    port map (
            O => \N__24476\,
            I => \N__24473\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__24473\,
            I => \N__24469\
        );

    \I__3629\ : InMux
    port map (
            O => \N__24472\,
            I => \N__24466\
        );

    \I__3628\ : Span4Mux_h
    port map (
            O => \N__24469\,
            I => \N__24460\
        );

    \I__3627\ : LocalMux
    port map (
            O => \N__24466\,
            I => \N__24460\
        );

    \I__3626\ : CascadeMux
    port map (
            O => \N__24465\,
            I => \N__24456\
        );

    \I__3625\ : Span4Mux_h
    port map (
            O => \N__24460\,
            I => \N__24453\
        );

    \I__3624\ : InMux
    port map (
            O => \N__24459\,
            I => \N__24448\
        );

    \I__3623\ : InMux
    port map (
            O => \N__24456\,
            I => \N__24448\
        );

    \I__3622\ : Odrv4
    port map (
            O => \N__24453\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__24448\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__3620\ : InMux
    port map (
            O => \N__24443\,
            I => \N__24439\
        );

    \I__3619\ : CascadeMux
    port map (
            O => \N__24442\,
            I => \N__24436\
        );

    \I__3618\ : LocalMux
    port map (
            O => \N__24439\,
            I => \N__24433\
        );

    \I__3617\ : InMux
    port map (
            O => \N__24436\,
            I => \N__24430\
        );

    \I__3616\ : Span4Mux_h
    port map (
            O => \N__24433\,
            I => \N__24427\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__24430\,
            I => \N__24424\
        );

    \I__3614\ : Span4Mux_v
    port map (
            O => \N__24427\,
            I => \N__24421\
        );

    \I__3613\ : Span4Mux_h
    port map (
            O => \N__24424\,
            I => \N__24418\
        );

    \I__3612\ : Odrv4
    port map (
            O => \N__24421\,
            I => \current_shift_inst.control_inputZ0Z_5\
        );

    \I__3611\ : Odrv4
    port map (
            O => \N__24418\,
            I => \current_shift_inst.control_inputZ0Z_5\
        );

    \I__3610\ : InMux
    port map (
            O => \N__24413\,
            I => \N__24410\
        );

    \I__3609\ : LocalMux
    port map (
            O => \N__24410\,
            I => \N__24407\
        );

    \I__3608\ : Span4Mux_h
    port map (
            O => \N__24407\,
            I => \N__24404\
        );

    \I__3607\ : Odrv4
    port map (
            O => \N__24404\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\
        );

    \I__3606\ : InMux
    port map (
            O => \N__24401\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\
        );

    \I__3605\ : InMux
    port map (
            O => \N__24398\,
            I => \N__24395\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__24395\,
            I => \N__24391\
        );

    \I__3603\ : InMux
    port map (
            O => \N__24394\,
            I => \N__24388\
        );

    \I__3602\ : Span4Mux_h
    port map (
            O => \N__24391\,
            I => \N__24381\
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__24388\,
            I => \N__24381\
        );

    \I__3600\ : InMux
    port map (
            O => \N__24387\,
            I => \N__24376\
        );

    \I__3599\ : InMux
    port map (
            O => \N__24386\,
            I => \N__24376\
        );

    \I__3598\ : Span4Mux_h
    port map (
            O => \N__24381\,
            I => \N__24373\
        );

    \I__3597\ : LocalMux
    port map (
            O => \N__24376\,
            I => \N__24370\
        );

    \I__3596\ : Odrv4
    port map (
            O => \N__24373\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__3595\ : Odrv4
    port map (
            O => \N__24370\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__3594\ : CascadeMux
    port map (
            O => \N__24365\,
            I => \N__24361\
        );

    \I__3593\ : InMux
    port map (
            O => \N__24364\,
            I => \N__24358\
        );

    \I__3592\ : InMux
    port map (
            O => \N__24361\,
            I => \N__24355\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__24358\,
            I => \N__24352\
        );

    \I__3590\ : LocalMux
    port map (
            O => \N__24355\,
            I => \N__24349\
        );

    \I__3589\ : Span4Mux_h
    port map (
            O => \N__24352\,
            I => \N__24344\
        );

    \I__3588\ : Span4Mux_h
    port map (
            O => \N__24349\,
            I => \N__24344\
        );

    \I__3587\ : Span4Mux_v
    port map (
            O => \N__24344\,
            I => \N__24341\
        );

    \I__3586\ : Odrv4
    port map (
            O => \N__24341\,
            I => \current_shift_inst.control_inputZ0Z_6\
        );

    \I__3585\ : InMux
    port map (
            O => \N__24338\,
            I => \N__24335\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__24335\,
            I => \N__24332\
        );

    \I__3583\ : Span4Mux_h
    port map (
            O => \N__24332\,
            I => \N__24329\
        );

    \I__3582\ : Odrv4
    port map (
            O => \N__24329\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\
        );

    \I__3581\ : InMux
    port map (
            O => \N__24326\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\
        );

    \I__3580\ : InMux
    port map (
            O => \N__24323\,
            I => \N__24320\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__24320\,
            I => \N__24317\
        );

    \I__3578\ : Span4Mux_h
    port map (
            O => \N__24317\,
            I => \N__24313\
        );

    \I__3577\ : InMux
    port map (
            O => \N__24316\,
            I => \N__24310\
        );

    \I__3576\ : Span4Mux_v
    port map (
            O => \N__24313\,
            I => \N__24307\
        );

    \I__3575\ : LocalMux
    port map (
            O => \N__24310\,
            I => \current_shift_inst.control_inputZ0Z_7\
        );

    \I__3574\ : Odrv4
    port map (
            O => \N__24307\,
            I => \current_shift_inst.control_inputZ0Z_7\
        );

    \I__3573\ : InMux
    port map (
            O => \N__24302\,
            I => \N__24299\
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__24299\,
            I => \N__24295\
        );

    \I__3571\ : CascadeMux
    port map (
            O => \N__24298\,
            I => \N__24292\
        );

    \I__3570\ : Span4Mux_h
    port map (
            O => \N__24295\,
            I => \N__24287\
        );

    \I__3569\ : InMux
    port map (
            O => \N__24292\,
            I => \N__24284\
        );

    \I__3568\ : InMux
    port map (
            O => \N__24291\,
            I => \N__24279\
        );

    \I__3567\ : InMux
    port map (
            O => \N__24290\,
            I => \N__24279\
        );

    \I__3566\ : Odrv4
    port map (
            O => \N__24287\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__3565\ : LocalMux
    port map (
            O => \N__24284\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__24279\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__3563\ : InMux
    port map (
            O => \N__24272\,
            I => \N__24269\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__24269\,
            I => \N__24266\
        );

    \I__3561\ : Odrv4
    port map (
            O => \N__24266\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\
        );

    \I__3560\ : InMux
    port map (
            O => \N__24263\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\
        );

    \I__3559\ : InMux
    port map (
            O => \N__24260\,
            I => \N__24257\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__24257\,
            I => \N__24251\
        );

    \I__3557\ : InMux
    port map (
            O => \N__24256\,
            I => \N__24248\
        );

    \I__3556\ : InMux
    port map (
            O => \N__24255\,
            I => \N__24243\
        );

    \I__3555\ : InMux
    port map (
            O => \N__24254\,
            I => \N__24243\
        );

    \I__3554\ : Odrv12
    port map (
            O => \N__24251\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__24248\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__3552\ : LocalMux
    port map (
            O => \N__24243\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__3551\ : InMux
    port map (
            O => \N__24236\,
            I => \N__24232\
        );

    \I__3550\ : CascadeMux
    port map (
            O => \N__24235\,
            I => \N__24229\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__24232\,
            I => \N__24226\
        );

    \I__3548\ : InMux
    port map (
            O => \N__24229\,
            I => \N__24223\
        );

    \I__3547\ : Span4Mux_v
    port map (
            O => \N__24226\,
            I => \N__24220\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__24223\,
            I => \N__24217\
        );

    \I__3545\ : Span4Mux_v
    port map (
            O => \N__24220\,
            I => \N__24214\
        );

    \I__3544\ : Span4Mux_h
    port map (
            O => \N__24217\,
            I => \N__24211\
        );

    \I__3543\ : Odrv4
    port map (
            O => \N__24214\,
            I => \current_shift_inst.control_inputZ0Z_8\
        );

    \I__3542\ : Odrv4
    port map (
            O => \N__24211\,
            I => \current_shift_inst.control_inputZ0Z_8\
        );

    \I__3541\ : InMux
    port map (
            O => \N__24206\,
            I => \N__24203\
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__24203\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\
        );

    \I__3539\ : InMux
    port map (
            O => \N__24200\,
            I => \bfn_9_14_0_\
        );

    \I__3538\ : InMux
    port map (
            O => \N__24197\,
            I => \N__24194\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__24194\,
            I => \N__24191\
        );

    \I__3536\ : Span4Mux_h
    port map (
            O => \N__24191\,
            I => \N__24185\
        );

    \I__3535\ : InMux
    port map (
            O => \N__24190\,
            I => \N__24180\
        );

    \I__3534\ : InMux
    port map (
            O => \N__24189\,
            I => \N__24180\
        );

    \I__3533\ : InMux
    port map (
            O => \N__24188\,
            I => \N__24177\
        );

    \I__3532\ : Odrv4
    port map (
            O => \N__24185\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__24180\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__24177\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__3529\ : InMux
    port map (
            O => \N__24170\,
            I => \N__24166\
        );

    \I__3528\ : CascadeMux
    port map (
            O => \N__24169\,
            I => \N__24163\
        );

    \I__3527\ : LocalMux
    port map (
            O => \N__24166\,
            I => \N__24160\
        );

    \I__3526\ : InMux
    port map (
            O => \N__24163\,
            I => \N__24157\
        );

    \I__3525\ : Span4Mux_h
    port map (
            O => \N__24160\,
            I => \N__24154\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__24157\,
            I => \N__24151\
        );

    \I__3523\ : Span4Mux_v
    port map (
            O => \N__24154\,
            I => \N__24148\
        );

    \I__3522\ : Span4Mux_h
    port map (
            O => \N__24151\,
            I => \N__24145\
        );

    \I__3521\ : Odrv4
    port map (
            O => \N__24148\,
            I => \current_shift_inst.control_inputZ0Z_9\
        );

    \I__3520\ : Odrv4
    port map (
            O => \N__24145\,
            I => \current_shift_inst.control_inputZ0Z_9\
        );

    \I__3519\ : InMux
    port map (
            O => \N__24140\,
            I => \N__24137\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__24137\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\
        );

    \I__3517\ : InMux
    port map (
            O => \N__24134\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\
        );

    \I__3516\ : InMux
    port map (
            O => \N__24131\,
            I => \N__24128\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__24128\,
            I => \N__24123\
        );

    \I__3514\ : InMux
    port map (
            O => \N__24127\,
            I => \N__24120\
        );

    \I__3513\ : InMux
    port map (
            O => \N__24126\,
            I => \N__24116\
        );

    \I__3512\ : Span4Mux_h
    port map (
            O => \N__24123\,
            I => \N__24111\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__24120\,
            I => \N__24111\
        );

    \I__3510\ : InMux
    port map (
            O => \N__24119\,
            I => \N__24108\
        );

    \I__3509\ : LocalMux
    port map (
            O => \N__24116\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__3508\ : Odrv4
    port map (
            O => \N__24111\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__3507\ : LocalMux
    port map (
            O => \N__24108\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__3506\ : CascadeMux
    port map (
            O => \N__24101\,
            I => \N__24097\
        );

    \I__3505\ : InMux
    port map (
            O => \N__24100\,
            I => \N__24094\
        );

    \I__3504\ : InMux
    port map (
            O => \N__24097\,
            I => \N__24091\
        );

    \I__3503\ : LocalMux
    port map (
            O => \N__24094\,
            I => \N__24088\
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__24091\,
            I => \N__24085\
        );

    \I__3501\ : Span4Mux_h
    port map (
            O => \N__24088\,
            I => \N__24080\
        );

    \I__3500\ : Span4Mux_h
    port map (
            O => \N__24085\,
            I => \N__24080\
        );

    \I__3499\ : Odrv4
    port map (
            O => \N__24080\,
            I => \current_shift_inst.control_inputZ0Z_10\
        );

    \I__3498\ : InMux
    port map (
            O => \N__24077\,
            I => \N__24074\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__24074\,
            I => \N__24071\
        );

    \I__3496\ : Odrv12
    port map (
            O => \N__24071\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\
        );

    \I__3495\ : InMux
    port map (
            O => \N__24068\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\
        );

    \I__3494\ : InMux
    port map (
            O => \N__24065\,
            I => \N__24060\
        );

    \I__3493\ : CascadeMux
    port map (
            O => \N__24064\,
            I => \N__24057\
        );

    \I__3492\ : InMux
    port map (
            O => \N__24063\,
            I => \N__24054\
        );

    \I__3491\ : LocalMux
    port map (
            O => \N__24060\,
            I => \N__24051\
        );

    \I__3490\ : InMux
    port map (
            O => \N__24057\,
            I => \N__24047\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__24054\,
            I => \N__24042\
        );

    \I__3488\ : Span4Mux_h
    port map (
            O => \N__24051\,
            I => \N__24042\
        );

    \I__3487\ : InMux
    port map (
            O => \N__24050\,
            I => \N__24039\
        );

    \I__3486\ : LocalMux
    port map (
            O => \N__24047\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__3485\ : Odrv4
    port map (
            O => \N__24042\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__24039\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__3483\ : InMux
    port map (
            O => \N__24032\,
            I => \N__24028\
        );

    \I__3482\ : CascadeMux
    port map (
            O => \N__24031\,
            I => \N__24025\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__24028\,
            I => \N__24022\
        );

    \I__3480\ : InMux
    port map (
            O => \N__24025\,
            I => \N__24019\
        );

    \I__3479\ : Span4Mux_v
    port map (
            O => \N__24022\,
            I => \N__24016\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__24019\,
            I => \N__24013\
        );

    \I__3477\ : Span4Mux_v
    port map (
            O => \N__24016\,
            I => \N__24010\
        );

    \I__3476\ : Span4Mux_h
    port map (
            O => \N__24013\,
            I => \N__24007\
        );

    \I__3475\ : Odrv4
    port map (
            O => \N__24010\,
            I => \current_shift_inst.control_inputZ0Z_11\
        );

    \I__3474\ : Odrv4
    port map (
            O => \N__24007\,
            I => \current_shift_inst.control_inputZ0Z_11\
        );

    \I__3473\ : InMux
    port map (
            O => \N__24002\,
            I => \N__23999\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__23999\,
            I => \N__23996\
        );

    \I__3471\ : Odrv12
    port map (
            O => \N__23996\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\
        );

    \I__3470\ : InMux
    port map (
            O => \N__23993\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\
        );

    \I__3469\ : InMux
    port map (
            O => \N__23990\,
            I => \N__23985\
        );

    \I__3468\ : InMux
    port map (
            O => \N__23989\,
            I => \N__23982\
        );

    \I__3467\ : InMux
    port map (
            O => \N__23988\,
            I => \N__23978\
        );

    \I__3466\ : LocalMux
    port map (
            O => \N__23985\,
            I => \N__23975\
        );

    \I__3465\ : LocalMux
    port map (
            O => \N__23982\,
            I => \N__23972\
        );

    \I__3464\ : InMux
    port map (
            O => \N__23981\,
            I => \N__23969\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__23978\,
            I => \N__23964\
        );

    \I__3462\ : Span4Mux_h
    port map (
            O => \N__23975\,
            I => \N__23964\
        );

    \I__3461\ : Odrv12
    port map (
            O => \N__23972\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__23969\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__3459\ : Odrv4
    port map (
            O => \N__23964\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__3458\ : CascadeMux
    port map (
            O => \N__23957\,
            I => \N__23953\
        );

    \I__3457\ : InMux
    port map (
            O => \N__23956\,
            I => \N__23950\
        );

    \I__3456\ : InMux
    port map (
            O => \N__23953\,
            I => \N__23947\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__23950\,
            I => \N__23944\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__23947\,
            I => \N__23941\
        );

    \I__3453\ : Span4Mux_h
    port map (
            O => \N__23944\,
            I => \N__23938\
        );

    \I__3452\ : Span4Mux_h
    port map (
            O => \N__23941\,
            I => \N__23935\
        );

    \I__3451\ : Odrv4
    port map (
            O => \N__23938\,
            I => \current_shift_inst.control_inputZ0Z_12\
        );

    \I__3450\ : Odrv4
    port map (
            O => \N__23935\,
            I => \current_shift_inst.control_inputZ0Z_12\
        );

    \I__3449\ : CascadeMux
    port map (
            O => \N__23930\,
            I => \N__23927\
        );

    \I__3448\ : InMux
    port map (
            O => \N__23927\,
            I => \N__23924\
        );

    \I__3447\ : LocalMux
    port map (
            O => \N__23924\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\
        );

    \I__3446\ : InMux
    port map (
            O => \N__23921\,
            I => \N__23918\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__23918\,
            I => \N__23915\
        );

    \I__3444\ : Odrv4
    port map (
            O => \N__23915\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0\
        );

    \I__3443\ : CascadeMux
    port map (
            O => \N__23912\,
            I => \N__23908\
        );

    \I__3442\ : InMux
    port map (
            O => \N__23911\,
            I => \N__23905\
        );

    \I__3441\ : InMux
    port map (
            O => \N__23908\,
            I => \N__23902\
        );

    \I__3440\ : LocalMux
    port map (
            O => \N__23905\,
            I => \N__23899\
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__23902\,
            I => \N__23896\
        );

    \I__3438\ : Span4Mux_h
    port map (
            O => \N__23899\,
            I => \N__23891\
        );

    \I__3437\ : Span4Mux_h
    port map (
            O => \N__23896\,
            I => \N__23891\
        );

    \I__3436\ : Odrv4
    port map (
            O => \N__23891\,
            I => \current_shift_inst.control_inputZ0Z_0\
        );

    \I__3435\ : InMux
    port map (
            O => \N__23888\,
            I => \N__23885\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__23885\,
            I => \N__23882\
        );

    \I__3433\ : Span4Mux_h
    port map (
            O => \N__23882\,
            I => \N__23877\
        );

    \I__3432\ : InMux
    port map (
            O => \N__23881\,
            I => \N__23874\
        );

    \I__3431\ : InMux
    port map (
            O => \N__23880\,
            I => \N__23871\
        );

    \I__3430\ : Odrv4
    port map (
            O => \N__23877\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_0\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__23874\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_0\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__23871\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_0\
        );

    \I__3427\ : InMux
    port map (
            O => \N__23864\,
            I => \N__23860\
        );

    \I__3426\ : CascadeMux
    port map (
            O => \N__23863\,
            I => \N__23857\
        );

    \I__3425\ : LocalMux
    port map (
            O => \N__23860\,
            I => \N__23854\
        );

    \I__3424\ : InMux
    port map (
            O => \N__23857\,
            I => \N__23851\
        );

    \I__3423\ : Span4Mux_h
    port map (
            O => \N__23854\,
            I => \N__23848\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__23851\,
            I => \N__23845\
        );

    \I__3421\ : Span4Mux_v
    port map (
            O => \N__23848\,
            I => \N__23842\
        );

    \I__3420\ : Span4Mux_h
    port map (
            O => \N__23845\,
            I => \N__23839\
        );

    \I__3419\ : Odrv4
    port map (
            O => \N__23842\,
            I => \current_shift_inst.control_inputZ0Z_1\
        );

    \I__3418\ : Odrv4
    port map (
            O => \N__23839\,
            I => \current_shift_inst.control_inputZ0Z_1\
        );

    \I__3417\ : InMux
    port map (
            O => \N__23834\,
            I => \N__23831\
        );

    \I__3416\ : LocalMux
    port map (
            O => \N__23831\,
            I => \N__23826\
        );

    \I__3415\ : InMux
    port map (
            O => \N__23830\,
            I => \N__23823\
        );

    \I__3414\ : InMux
    port map (
            O => \N__23829\,
            I => \N__23820\
        );

    \I__3413\ : Span4Mux_h
    port map (
            O => \N__23826\,
            I => \N__23815\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__23823\,
            I => \N__23815\
        );

    \I__3411\ : LocalMux
    port map (
            O => \N__23820\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__3410\ : Odrv4
    port map (
            O => \N__23815\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__3409\ : InMux
    port map (
            O => \N__23810\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_0\
        );

    \I__3408\ : CascadeMux
    port map (
            O => \N__23807\,
            I => \N__23803\
        );

    \I__3407\ : InMux
    port map (
            O => \N__23806\,
            I => \N__23800\
        );

    \I__3406\ : InMux
    port map (
            O => \N__23803\,
            I => \N__23797\
        );

    \I__3405\ : LocalMux
    port map (
            O => \N__23800\,
            I => \N__23794\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__23797\,
            I => \N__23791\
        );

    \I__3403\ : Span4Mux_h
    port map (
            O => \N__23794\,
            I => \N__23786\
        );

    \I__3402\ : Span4Mux_h
    port map (
            O => \N__23791\,
            I => \N__23786\
        );

    \I__3401\ : Odrv4
    port map (
            O => \N__23786\,
            I => \current_shift_inst.control_inputZ0Z_2\
        );

    \I__3400\ : InMux
    port map (
            O => \N__23783\,
            I => \N__23780\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__23780\,
            I => \N__23775\
        );

    \I__3398\ : InMux
    port map (
            O => \N__23779\,
            I => \N__23772\
        );

    \I__3397\ : InMux
    port map (
            O => \N__23778\,
            I => \N__23769\
        );

    \I__3396\ : Span4Mux_h
    port map (
            O => \N__23775\,
            I => \N__23762\
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__23772\,
            I => \N__23762\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__23769\,
            I => \N__23762\
        );

    \I__3393\ : Odrv4
    port map (
            O => \N__23762\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__3392\ : InMux
    port map (
            O => \N__23759\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\
        );

    \I__3391\ : InMux
    port map (
            O => \N__23756\,
            I => \N__23750\
        );

    \I__3390\ : InMux
    port map (
            O => \N__23755\,
            I => \N__23743\
        );

    \I__3389\ : InMux
    port map (
            O => \N__23754\,
            I => \N__23743\
        );

    \I__3388\ : InMux
    port map (
            O => \N__23753\,
            I => \N__23743\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__23750\,
            I => \N__23738\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__23743\,
            I => \N__23738\
        );

    \I__3385\ : Odrv4
    port map (
            O => \N__23738\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__3384\ : CascadeMux
    port map (
            O => \N__23735\,
            I => \N__23731\
        );

    \I__3383\ : InMux
    port map (
            O => \N__23734\,
            I => \N__23728\
        );

    \I__3382\ : InMux
    port map (
            O => \N__23731\,
            I => \N__23725\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__23728\,
            I => \N__23722\
        );

    \I__3380\ : LocalMux
    port map (
            O => \N__23725\,
            I => \N__23719\
        );

    \I__3379\ : Span4Mux_h
    port map (
            O => \N__23722\,
            I => \N__23714\
        );

    \I__3378\ : Span4Mux_h
    port map (
            O => \N__23719\,
            I => \N__23714\
        );

    \I__3377\ : Odrv4
    port map (
            O => \N__23714\,
            I => \current_shift_inst.control_inputZ0Z_3\
        );

    \I__3376\ : InMux
    port map (
            O => \N__23711\,
            I => \N__23705\
        );

    \I__3375\ : InMux
    port map (
            O => \N__23710\,
            I => \N__23700\
        );

    \I__3374\ : InMux
    port map (
            O => \N__23709\,
            I => \N__23700\
        );

    \I__3373\ : InMux
    port map (
            O => \N__23708\,
            I => \N__23697\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__23705\,
            I => \N__23692\
        );

    \I__3371\ : LocalMux
    port map (
            O => \N__23700\,
            I => \N__23692\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__23697\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__3369\ : Odrv12
    port map (
            O => \N__23692\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__3368\ : InMux
    port map (
            O => \N__23687\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\
        );

    \I__3367\ : CEMux
    port map (
            O => \N__23684\,
            I => \N__23680\
        );

    \I__3366\ : CEMux
    port map (
            O => \N__23683\,
            I => \N__23668\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__23680\,
            I => \N__23665\
        );

    \I__3364\ : CEMux
    port map (
            O => \N__23679\,
            I => \N__23662\
        );

    \I__3363\ : CEMux
    port map (
            O => \N__23678\,
            I => \N__23659\
        );

    \I__3362\ : CEMux
    port map (
            O => \N__23677\,
            I => \N__23656\
        );

    \I__3361\ : CEMux
    port map (
            O => \N__23676\,
            I => \N__23653\
        );

    \I__3360\ : CEMux
    port map (
            O => \N__23675\,
            I => \N__23650\
        );

    \I__3359\ : CEMux
    port map (
            O => \N__23674\,
            I => \N__23645\
        );

    \I__3358\ : CEMux
    port map (
            O => \N__23673\,
            I => \N__23642\
        );

    \I__3357\ : CEMux
    port map (
            O => \N__23672\,
            I => \N__23638\
        );

    \I__3356\ : CEMux
    port map (
            O => \N__23671\,
            I => \N__23632\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__23668\,
            I => \N__23628\
        );

    \I__3354\ : Span4Mux_h
    port map (
            O => \N__23665\,
            I => \N__23623\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__23662\,
            I => \N__23623\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__23659\,
            I => \N__23616\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__23656\,
            I => \N__23616\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__23653\,
            I => \N__23616\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__23650\,
            I => \N__23613\
        );

    \I__3348\ : CEMux
    port map (
            O => \N__23649\,
            I => \N__23610\
        );

    \I__3347\ : CEMux
    port map (
            O => \N__23648\,
            I => \N__23607\
        );

    \I__3346\ : LocalMux
    port map (
            O => \N__23645\,
            I => \N__23604\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__23642\,
            I => \N__23601\
        );

    \I__3344\ : CEMux
    port map (
            O => \N__23641\,
            I => \N__23598\
        );

    \I__3343\ : LocalMux
    port map (
            O => \N__23638\,
            I => \N__23595\
        );

    \I__3342\ : CEMux
    port map (
            O => \N__23637\,
            I => \N__23592\
        );

    \I__3341\ : CEMux
    port map (
            O => \N__23636\,
            I => \N__23589\
        );

    \I__3340\ : CEMux
    port map (
            O => \N__23635\,
            I => \N__23586\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__23632\,
            I => \N__23582\
        );

    \I__3338\ : CEMux
    port map (
            O => \N__23631\,
            I => \N__23579\
        );

    \I__3337\ : Span4Mux_v
    port map (
            O => \N__23628\,
            I => \N__23573\
        );

    \I__3336\ : Span4Mux_v
    port map (
            O => \N__23623\,
            I => \N__23573\
        );

    \I__3335\ : Span4Mux_v
    port map (
            O => \N__23616\,
            I => \N__23566\
        );

    \I__3334\ : Span4Mux_v
    port map (
            O => \N__23613\,
            I => \N__23566\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__23610\,
            I => \N__23566\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__23607\,
            I => \N__23563\
        );

    \I__3331\ : Span4Mux_v
    port map (
            O => \N__23604\,
            I => \N__23560\
        );

    \I__3330\ : Span4Mux_v
    port map (
            O => \N__23601\,
            I => \N__23555\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__23598\,
            I => \N__23555\
        );

    \I__3328\ : Span4Mux_h
    port map (
            O => \N__23595\,
            I => \N__23552\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__23592\,
            I => \N__23545\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__23589\,
            I => \N__23545\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__23586\,
            I => \N__23545\
        );

    \I__3324\ : CEMux
    port map (
            O => \N__23585\,
            I => \N__23542\
        );

    \I__3323\ : Sp12to4
    port map (
            O => \N__23582\,
            I => \N__23537\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__23579\,
            I => \N__23537\
        );

    \I__3321\ : CEMux
    port map (
            O => \N__23578\,
            I => \N__23534\
        );

    \I__3320\ : Span4Mux_v
    port map (
            O => \N__23573\,
            I => \N__23531\
        );

    \I__3319\ : Span4Mux_v
    port map (
            O => \N__23566\,
            I => \N__23526\
        );

    \I__3318\ : Span4Mux_h
    port map (
            O => \N__23563\,
            I => \N__23526\
        );

    \I__3317\ : Span4Mux_h
    port map (
            O => \N__23560\,
            I => \N__23517\
        );

    \I__3316\ : Span4Mux_v
    port map (
            O => \N__23555\,
            I => \N__23517\
        );

    \I__3315\ : Span4Mux_h
    port map (
            O => \N__23552\,
            I => \N__23517\
        );

    \I__3314\ : Span4Mux_v
    port map (
            O => \N__23545\,
            I => \N__23517\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__23542\,
            I => \N__23514\
        );

    \I__3312\ : Span12Mux_v
    port map (
            O => \N__23537\,
            I => \N__23509\
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__23534\,
            I => \N__23509\
        );

    \I__3310\ : Odrv4
    port map (
            O => \N__23531\,
            I => \N_702_g\
        );

    \I__3309\ : Odrv4
    port map (
            O => \N__23526\,
            I => \N_702_g\
        );

    \I__3308\ : Odrv4
    port map (
            O => \N__23517\,
            I => \N_702_g\
        );

    \I__3307\ : Odrv12
    port map (
            O => \N__23514\,
            I => \N_702_g\
        );

    \I__3306\ : Odrv12
    port map (
            O => \N__23509\,
            I => \N_702_g\
        );

    \I__3305\ : CascadeMux
    port map (
            O => \N__23498\,
            I => \N__23494\
        );

    \I__3304\ : InMux
    port map (
            O => \N__23497\,
            I => \N__23490\
        );

    \I__3303\ : InMux
    port map (
            O => \N__23494\,
            I => \N__23486\
        );

    \I__3302\ : InMux
    port map (
            O => \N__23493\,
            I => \N__23483\
        );

    \I__3301\ : LocalMux
    port map (
            O => \N__23490\,
            I => \N__23480\
        );

    \I__3300\ : InMux
    port map (
            O => \N__23489\,
            I => \N__23477\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__23486\,
            I => \N__23468\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__23483\,
            I => \N__23468\
        );

    \I__3297\ : Span4Mux_h
    port map (
            O => \N__23480\,
            I => \N__23468\
        );

    \I__3296\ : LocalMux
    port map (
            O => \N__23477\,
            I => \N__23468\
        );

    \I__3295\ : Span4Mux_h
    port map (
            O => \N__23468\,
            I => \N__23465\
        );

    \I__3294\ : Odrv4
    port map (
            O => \N__23465\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__3293\ : CascadeMux
    port map (
            O => \N__23462\,
            I => \N__23458\
        );

    \I__3292\ : InMux
    port map (
            O => \N__23461\,
            I => \N__23455\
        );

    \I__3291\ : InMux
    port map (
            O => \N__23458\,
            I => \N__23452\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__23455\,
            I => \N__23449\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__23452\,
            I => \N__23446\
        );

    \I__3288\ : Span4Mux_h
    port map (
            O => \N__23449\,
            I => \N__23441\
        );

    \I__3287\ : Span4Mux_h
    port map (
            O => \N__23446\,
            I => \N__23441\
        );

    \I__3286\ : Odrv4
    port map (
            O => \N__23441\,
            I => \current_shift_inst.control_inputZ0Z_4\
        );

    \I__3285\ : CascadeMux
    port map (
            O => \N__23438\,
            I => \N__23435\
        );

    \I__3284\ : InMux
    port map (
            O => \N__23435\,
            I => \N__23432\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__23432\,
            I => \N__23429\
        );

    \I__3282\ : Span4Mux_h
    port map (
            O => \N__23429\,
            I => \N__23426\
        );

    \I__3281\ : Odrv4
    port map (
            O => \N__23426\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\
        );

    \I__3280\ : InMux
    port map (
            O => \N__23423\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\
        );

    \I__3279\ : CascadeMux
    port map (
            O => \N__23420\,
            I => \N__23417\
        );

    \I__3278\ : InMux
    port map (
            O => \N__23417\,
            I => \N__23414\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__23414\,
            I => \N__23411\
        );

    \I__3276\ : Odrv4
    port map (
            O => \N__23411\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\
        );

    \I__3275\ : CascadeMux
    port map (
            O => \N__23408\,
            I => \N__23405\
        );

    \I__3274\ : InMux
    port map (
            O => \N__23405\,
            I => \N__23402\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__23402\,
            I => \N__23399\
        );

    \I__3272\ : Odrv4
    port map (
            O => \N__23399\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\
        );

    \I__3271\ : CascadeMux
    port map (
            O => \N__23396\,
            I => \N__23393\
        );

    \I__3270\ : InMux
    port map (
            O => \N__23393\,
            I => \N__23390\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__23390\,
            I => \N__23387\
        );

    \I__3268\ : Span4Mux_h
    port map (
            O => \N__23387\,
            I => \N__23384\
        );

    \I__3267\ : Odrv4
    port map (
            O => \N__23384\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\
        );

    \I__3266\ : CascadeMux
    port map (
            O => \N__23381\,
            I => \N__23378\
        );

    \I__3265\ : InMux
    port map (
            O => \N__23378\,
            I => \N__23375\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__23375\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_0\
        );

    \I__3263\ : CascadeMux
    port map (
            O => \N__23372\,
            I => \N__23369\
        );

    \I__3262\ : InMux
    port map (
            O => \N__23369\,
            I => \N__23366\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__23366\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\
        );

    \I__3260\ : CascadeMux
    port map (
            O => \N__23363\,
            I => \N__23360\
        );

    \I__3259\ : InMux
    port map (
            O => \N__23360\,
            I => \N__23357\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__23357\,
            I => \N__23354\
        );

    \I__3257\ : Odrv4
    port map (
            O => \N__23354\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\
        );

    \I__3256\ : CascadeMux
    port map (
            O => \N__23351\,
            I => \N__23348\
        );

    \I__3255\ : InMux
    port map (
            O => \N__23348\,
            I => \N__23345\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__23345\,
            I => \N__23342\
        );

    \I__3253\ : Odrv4
    port map (
            O => \N__23342\,
            I => \pwm_generator_inst.thresholdZ0Z_6\
        );

    \I__3252\ : InMux
    port map (
            O => \N__23339\,
            I => \N__23336\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__23336\,
            I => \pwm_generator_inst.counter_i_6\
        );

    \I__3250\ : InMux
    port map (
            O => \N__23333\,
            I => \N__23330\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__23330\,
            I => \N__23327\
        );

    \I__3248\ : Odrv12
    port map (
            O => \N__23327\,
            I => \pwm_generator_inst.thresholdZ0Z_7\
        );

    \I__3247\ : CascadeMux
    port map (
            O => \N__23324\,
            I => \N__23321\
        );

    \I__3246\ : InMux
    port map (
            O => \N__23321\,
            I => \N__23318\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__23318\,
            I => \pwm_generator_inst.counter_i_7\
        );

    \I__3244\ : CascadeMux
    port map (
            O => \N__23315\,
            I => \N__23312\
        );

    \I__3243\ : InMux
    port map (
            O => \N__23312\,
            I => \N__23309\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__23309\,
            I => \N__23306\
        );

    \I__3241\ : Span4Mux_h
    port map (
            O => \N__23306\,
            I => \N__23303\
        );

    \I__3240\ : Odrv4
    port map (
            O => \N__23303\,
            I => \pwm_generator_inst.thresholdZ0Z_8\
        );

    \I__3239\ : InMux
    port map (
            O => \N__23300\,
            I => \N__23297\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__23297\,
            I => \pwm_generator_inst.counter_i_8\
        );

    \I__3237\ : CascadeMux
    port map (
            O => \N__23294\,
            I => \N__23291\
        );

    \I__3236\ : InMux
    port map (
            O => \N__23291\,
            I => \N__23288\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__23288\,
            I => \N__23285\
        );

    \I__3234\ : Span4Mux_h
    port map (
            O => \N__23285\,
            I => \N__23282\
        );

    \I__3233\ : Odrv4
    port map (
            O => \N__23282\,
            I => \pwm_generator_inst.thresholdZ0Z_9\
        );

    \I__3232\ : InMux
    port map (
            O => \N__23279\,
            I => \N__23276\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__23276\,
            I => \pwm_generator_inst.counter_i_9\
        );

    \I__3230\ : InMux
    port map (
            O => \N__23273\,
            I => \pwm_generator_inst.un14_counter_cry_9\
        );

    \I__3229\ : IoInMux
    port map (
            O => \N__23270\,
            I => \N__23267\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__23267\,
            I => \N__23264\
        );

    \I__3227\ : Span4Mux_s3_v
    port map (
            O => \N__23264\,
            I => \N__23261\
        );

    \I__3226\ : Span4Mux_v
    port map (
            O => \N__23261\,
            I => \N__23258\
        );

    \I__3225\ : Span4Mux_h
    port map (
            O => \N__23258\,
            I => \N__23255\
        );

    \I__3224\ : Span4Mux_h
    port map (
            O => \N__23255\,
            I => \N__23252\
        );

    \I__3223\ : Span4Mux_h
    port map (
            O => \N__23252\,
            I => \N__23249\
        );

    \I__3222\ : Odrv4
    port map (
            O => \N__23249\,
            I => pwm_output_c
        );

    \I__3221\ : InMux
    port map (
            O => \N__23246\,
            I => \N__23243\
        );

    \I__3220\ : LocalMux
    port map (
            O => \N__23243\,
            I => \il_min_comp2_D1\
        );

    \I__3219\ : InMux
    port map (
            O => \N__23240\,
            I => \N__23237\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__23237\,
            I => \N__23234\
        );

    \I__3217\ : Span4Mux_h
    port map (
            O => \N__23234\,
            I => \N__23231\
        );

    \I__3216\ : Span4Mux_v
    port map (
            O => \N__23231\,
            I => \N__23228\
        );

    \I__3215\ : Odrv4
    port map (
            O => \N__23228\,
            I => il_max_comp1_c
        );

    \I__3214\ : CascadeMux
    port map (
            O => \N__23225\,
            I => \N__23222\
        );

    \I__3213\ : InMux
    port map (
            O => \N__23222\,
            I => \N__23219\
        );

    \I__3212\ : LocalMux
    port map (
            O => \N__23219\,
            I => \pwm_generator_inst.thresholdZ0Z_0\
        );

    \I__3211\ : InMux
    port map (
            O => \N__23216\,
            I => \N__23213\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__23213\,
            I => \pwm_generator_inst.counter_i_0\
        );

    \I__3209\ : InMux
    port map (
            O => \N__23210\,
            I => \N__23207\
        );

    \I__3208\ : LocalMux
    port map (
            O => \N__23207\,
            I => \N__23204\
        );

    \I__3207\ : Odrv4
    port map (
            O => \N__23204\,
            I => \pwm_generator_inst.thresholdZ0Z_1\
        );

    \I__3206\ : CascadeMux
    port map (
            O => \N__23201\,
            I => \N__23198\
        );

    \I__3205\ : InMux
    port map (
            O => \N__23198\,
            I => \N__23195\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__23195\,
            I => \pwm_generator_inst.counter_i_1\
        );

    \I__3203\ : CascadeMux
    port map (
            O => \N__23192\,
            I => \N__23189\
        );

    \I__3202\ : InMux
    port map (
            O => \N__23189\,
            I => \N__23186\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__23186\,
            I => \N__23183\
        );

    \I__3200\ : Odrv12
    port map (
            O => \N__23183\,
            I => \pwm_generator_inst.thresholdZ0Z_2\
        );

    \I__3199\ : InMux
    port map (
            O => \N__23180\,
            I => \N__23177\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__23177\,
            I => \pwm_generator_inst.counter_i_2\
        );

    \I__3197\ : InMux
    port map (
            O => \N__23174\,
            I => \N__23171\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__23171\,
            I => \pwm_generator_inst.thresholdZ0Z_3\
        );

    \I__3195\ : CascadeMux
    port map (
            O => \N__23168\,
            I => \N__23165\
        );

    \I__3194\ : InMux
    port map (
            O => \N__23165\,
            I => \N__23162\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__23162\,
            I => \pwm_generator_inst.counter_i_3\
        );

    \I__3192\ : InMux
    port map (
            O => \N__23159\,
            I => \N__23156\
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__23156\,
            I => \N__23153\
        );

    \I__3190\ : Span4Mux_h
    port map (
            O => \N__23153\,
            I => \N__23150\
        );

    \I__3189\ : Odrv4
    port map (
            O => \N__23150\,
            I => \pwm_generator_inst.thresholdZ0Z_4\
        );

    \I__3188\ : CascadeMux
    port map (
            O => \N__23147\,
            I => \N__23144\
        );

    \I__3187\ : InMux
    port map (
            O => \N__23144\,
            I => \N__23141\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__23141\,
            I => \N__23138\
        );

    \I__3185\ : Odrv4
    port map (
            O => \N__23138\,
            I => \pwm_generator_inst.counter_i_4\
        );

    \I__3184\ : CascadeMux
    port map (
            O => \N__23135\,
            I => \N__23132\
        );

    \I__3183\ : InMux
    port map (
            O => \N__23132\,
            I => \N__23129\
        );

    \I__3182\ : LocalMux
    port map (
            O => \N__23129\,
            I => \N__23126\
        );

    \I__3181\ : Odrv4
    port map (
            O => \N__23126\,
            I => \pwm_generator_inst.thresholdZ0Z_5\
        );

    \I__3180\ : InMux
    port map (
            O => \N__23123\,
            I => \N__23120\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__23120\,
            I => \pwm_generator_inst.counter_i_5\
        );

    \I__3178\ : InMux
    port map (
            O => \N__23117\,
            I => \N__23114\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__23114\,
            I => \current_shift_inst.control_input_1_axb_18\
        );

    \I__3176\ : InMux
    port map (
            O => \N__23111\,
            I => \current_shift_inst.un38_control_input_0_cry_23\
        );

    \I__3175\ : InMux
    port map (
            O => \N__23108\,
            I => \N__23105\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__23105\,
            I => \current_shift_inst.control_input_1_axb_19\
        );

    \I__3173\ : InMux
    port map (
            O => \N__23102\,
            I => \current_shift_inst.un38_control_input_0_cry_24\
        );

    \I__3172\ : InMux
    port map (
            O => \N__23099\,
            I => \N__23096\
        );

    \I__3171\ : LocalMux
    port map (
            O => \N__23096\,
            I => \current_shift_inst.control_input_1_axb_20\
        );

    \I__3170\ : InMux
    port map (
            O => \N__23093\,
            I => \current_shift_inst.un38_control_input_0_cry_25\
        );

    \I__3169\ : InMux
    port map (
            O => \N__23090\,
            I => \N__23087\
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__23087\,
            I => \current_shift_inst.control_input_1_axb_21\
        );

    \I__3167\ : InMux
    port map (
            O => \N__23084\,
            I => \current_shift_inst.un38_control_input_0_cry_26\
        );

    \I__3166\ : InMux
    port map (
            O => \N__23081\,
            I => \N__23078\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__23078\,
            I => \current_shift_inst.control_input_1_axb_22\
        );

    \I__3164\ : InMux
    port map (
            O => \N__23075\,
            I => \current_shift_inst.un38_control_input_0_cry_27\
        );

    \I__3163\ : InMux
    port map (
            O => \N__23072\,
            I => \N__23069\
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__23069\,
            I => \current_shift_inst.control_input_1_axb_23\
        );

    \I__3161\ : InMux
    port map (
            O => \N__23066\,
            I => \current_shift_inst.un38_control_input_0_cry_28\
        );

    \I__3160\ : InMux
    port map (
            O => \N__23063\,
            I => \N__23060\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__23060\,
            I => \current_shift_inst.control_input_1_axb_24\
        );

    \I__3158\ : InMux
    port map (
            O => \N__23057\,
            I => \current_shift_inst.un38_control_input_0_cry_29\
        );

    \I__3157\ : CascadeMux
    port map (
            O => \N__23054\,
            I => \N__23051\
        );

    \I__3156\ : InMux
    port map (
            O => \N__23051\,
            I => \N__23048\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__23048\,
            I => \current_shift_inst.control_input_1_cry_24_THRU_CO\
        );

    \I__3154\ : InMux
    port map (
            O => \N__23045\,
            I => \bfn_8_21_0_\
        );

    \I__3153\ : CEMux
    port map (
            O => \N__23042\,
            I => \N__23039\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__23039\,
            I => \N__23034\
        );

    \I__3151\ : CEMux
    port map (
            O => \N__23038\,
            I => \N__23031\
        );

    \I__3150\ : CEMux
    port map (
            O => \N__23037\,
            I => \N__23028\
        );

    \I__3149\ : Span4Mux_h
    port map (
            O => \N__23034\,
            I => \N__23021\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__23031\,
            I => \N__23021\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__23028\,
            I => \N__23018\
        );

    \I__3146\ : CEMux
    port map (
            O => \N__23027\,
            I => \N__23015\
        );

    \I__3145\ : CEMux
    port map (
            O => \N__23026\,
            I => \N__23012\
        );

    \I__3144\ : Span4Mux_v
    port map (
            O => \N__23021\,
            I => \N__23005\
        );

    \I__3143\ : Span4Mux_v
    port map (
            O => \N__23018\,
            I => \N__23005\
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__23015\,
            I => \N__23005\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__23012\,
            I => \N__23002\
        );

    \I__3140\ : Span4Mux_v
    port map (
            O => \N__23005\,
            I => \N__22999\
        );

    \I__3139\ : Span12Mux_v
    port map (
            O => \N__23002\,
            I => \N__22996\
        );

    \I__3138\ : Span4Mux_v
    port map (
            O => \N__22999\,
            I => \N__22993\
        );

    \I__3137\ : Odrv12
    port map (
            O => \N__22996\,
            I => \current_shift_inst.phase_valid_RNISLORZ0Z2\
        );

    \I__3136\ : Odrv4
    port map (
            O => \N__22993\,
            I => \current_shift_inst.phase_valid_RNISLORZ0Z2\
        );

    \I__3135\ : InMux
    port map (
            O => \N__22988\,
            I => \N__22985\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__22985\,
            I => \current_shift_inst.control_input_1_axb_9\
        );

    \I__3133\ : InMux
    port map (
            O => \N__22982\,
            I => \bfn_8_19_0_\
        );

    \I__3132\ : InMux
    port map (
            O => \N__22979\,
            I => \N__22976\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__22976\,
            I => \current_shift_inst.control_input_1_axb_10\
        );

    \I__3130\ : InMux
    port map (
            O => \N__22973\,
            I => \current_shift_inst.un38_control_input_0_cry_15\
        );

    \I__3129\ : InMux
    port map (
            O => \N__22970\,
            I => \N__22967\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__22967\,
            I => \current_shift_inst.control_input_1_axb_11\
        );

    \I__3127\ : InMux
    port map (
            O => \N__22964\,
            I => \current_shift_inst.un38_control_input_0_cry_16\
        );

    \I__3126\ : CascadeMux
    port map (
            O => \N__22961\,
            I => \N__22958\
        );

    \I__3125\ : InMux
    port map (
            O => \N__22958\,
            I => \N__22955\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__22955\,
            I => \N__22952\
        );

    \I__3123\ : Odrv4
    port map (
            O => \N__22952\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIH6661_17\
        );

    \I__3122\ : InMux
    port map (
            O => \N__22949\,
            I => \N__22946\
        );

    \I__3121\ : LocalMux
    port map (
            O => \N__22946\,
            I => \current_shift_inst.control_input_1_axb_12\
        );

    \I__3120\ : InMux
    port map (
            O => \N__22943\,
            I => \current_shift_inst.un38_control_input_0_cry_17\
        );

    \I__3119\ : CascadeMux
    port map (
            O => \N__22940\,
            I => \N__22937\
        );

    \I__3118\ : InMux
    port map (
            O => \N__22937\,
            I => \N__22934\
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__22934\,
            I => \N__22931\
        );

    \I__3116\ : Odrv12
    port map (
            O => \N__22931\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIAL3J_18\
        );

    \I__3115\ : InMux
    port map (
            O => \N__22928\,
            I => \N__22925\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__22925\,
            I => \current_shift_inst.control_input_1_axb_13\
        );

    \I__3113\ : InMux
    port map (
            O => \N__22922\,
            I => \current_shift_inst.un38_control_input_0_cry_18\
        );

    \I__3112\ : CascadeMux
    port map (
            O => \N__22919\,
            I => \N__22916\
        );

    \I__3111\ : InMux
    port map (
            O => \N__22916\,
            I => \N__22913\
        );

    \I__3110\ : LocalMux
    port map (
            O => \N__22913\,
            I => \N__22910\
        );

    \I__3109\ : Odrv4
    port map (
            O => \N__22910\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI4H5J_19\
        );

    \I__3108\ : InMux
    port map (
            O => \N__22907\,
            I => \N__22904\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__22904\,
            I => \current_shift_inst.control_input_1_axb_14\
        );

    \I__3106\ : InMux
    port map (
            O => \N__22901\,
            I => \current_shift_inst.un38_control_input_0_cry_19\
        );

    \I__3105\ : InMux
    port map (
            O => \N__22898\,
            I => \N__22895\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__22895\,
            I => \current_shift_inst.control_input_1_axb_15\
        );

    \I__3103\ : InMux
    port map (
            O => \N__22892\,
            I => \current_shift_inst.un38_control_input_0_cry_20\
        );

    \I__3102\ : InMux
    port map (
            O => \N__22889\,
            I => \N__22886\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__22886\,
            I => \current_shift_inst.control_input_1_axb_16\
        );

    \I__3100\ : InMux
    port map (
            O => \N__22883\,
            I => \current_shift_inst.un38_control_input_0_cry_21\
        );

    \I__3099\ : InMux
    port map (
            O => \N__22880\,
            I => \N__22877\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__22877\,
            I => \current_shift_inst.control_input_1_axb_17\
        );

    \I__3097\ : InMux
    port map (
            O => \N__22874\,
            I => \bfn_8_20_0_\
        );

    \I__3096\ : InMux
    port map (
            O => \N__22871\,
            I => \N__22868\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__22868\,
            I => \current_shift_inst.control_input_1_axb_1\
        );

    \I__3094\ : InMux
    port map (
            O => \N__22865\,
            I => \bfn_8_18_0_\
        );

    \I__3093\ : InMux
    port map (
            O => \N__22862\,
            I => \N__22859\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__22859\,
            I => \current_shift_inst.control_input_1_axb_2\
        );

    \I__3091\ : InMux
    port map (
            O => \N__22856\,
            I => \current_shift_inst.un38_control_input_0_cry_7\
        );

    \I__3090\ : InMux
    port map (
            O => \N__22853\,
            I => \N__22850\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__22850\,
            I => \current_shift_inst.control_input_1_axb_3\
        );

    \I__3088\ : InMux
    port map (
            O => \N__22847\,
            I => \current_shift_inst.un38_control_input_0_cry_8\
        );

    \I__3087\ : InMux
    port map (
            O => \N__22844\,
            I => \N__22841\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__22841\,
            I => \current_shift_inst.control_input_1_axb_4\
        );

    \I__3085\ : InMux
    port map (
            O => \N__22838\,
            I => \current_shift_inst.un38_control_input_0_cry_9\
        );

    \I__3084\ : InMux
    port map (
            O => \N__22835\,
            I => \N__22832\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__22832\,
            I => \current_shift_inst.control_input_1_axb_5\
        );

    \I__3082\ : InMux
    port map (
            O => \N__22829\,
            I => \current_shift_inst.un38_control_input_0_cry_10\
        );

    \I__3081\ : InMux
    port map (
            O => \N__22826\,
            I => \N__22823\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__22823\,
            I => \current_shift_inst.control_input_1_axb_6\
        );

    \I__3079\ : InMux
    port map (
            O => \N__22820\,
            I => \current_shift_inst.un38_control_input_0_cry_11\
        );

    \I__3078\ : InMux
    port map (
            O => \N__22817\,
            I => \N__22814\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__22814\,
            I => \current_shift_inst.control_input_1_axb_7\
        );

    \I__3076\ : InMux
    port map (
            O => \N__22811\,
            I => \current_shift_inst.un38_control_input_0_cry_12\
        );

    \I__3075\ : CascadeMux
    port map (
            O => \N__22808\,
            I => \N__22805\
        );

    \I__3074\ : InMux
    port map (
            O => \N__22805\,
            I => \N__22802\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__22802\,
            I => \N__22799\
        );

    \I__3072\ : Odrv4
    port map (
            O => \N__22799\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIR0UI_13\
        );

    \I__3071\ : InMux
    port map (
            O => \N__22796\,
            I => \N__22793\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__22793\,
            I => \current_shift_inst.control_input_1_axb_8\
        );

    \I__3069\ : InMux
    port map (
            O => \N__22790\,
            I => \current_shift_inst.un38_control_input_0_cry_13\
        );

    \I__3068\ : InMux
    port map (
            O => \N__22787\,
            I => \N__22784\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__22784\,
            I => \current_shift_inst.z_i_0_31\
        );

    \I__3066\ : CascadeMux
    port map (
            O => \N__22781\,
            I => \N__22778\
        );

    \I__3065\ : InMux
    port map (
            O => \N__22778\,
            I => \N__22775\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__22775\,
            I => \current_shift_inst.un38_control_input_0_cry_3_c_invZ0\
        );

    \I__3063\ : InMux
    port map (
            O => \N__22772\,
            I => \N__22769\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__22769\,
            I => \current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0\
        );

    \I__3061\ : CascadeMux
    port map (
            O => \N__22766\,
            I => \N__22763\
        );

    \I__3060\ : InMux
    port map (
            O => \N__22763\,
            I => \N__22760\
        );

    \I__3059\ : LocalMux
    port map (
            O => \N__22760\,
            I => \current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0Z_0\
        );

    \I__3058\ : InMux
    port map (
            O => \N__22757\,
            I => \N__22754\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__22754\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIVQKU1_5\
        );

    \I__3056\ : InMux
    port map (
            O => \N__22751\,
            I => \N__22748\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__22748\,
            I => \current_shift_inst.control_input_1_axb_0\
        );

    \I__3054\ : InMux
    port map (
            O => \N__22745\,
            I => \current_shift_inst.un38_control_input_0_cry_5\
        );

    \I__3053\ : InMux
    port map (
            O => \N__22742\,
            I => \N__22727\
        );

    \I__3052\ : InMux
    port map (
            O => \N__22741\,
            I => \N__22727\
        );

    \I__3051\ : InMux
    port map (
            O => \N__22740\,
            I => \N__22714\
        );

    \I__3050\ : InMux
    port map (
            O => \N__22739\,
            I => \N__22714\
        );

    \I__3049\ : InMux
    port map (
            O => \N__22738\,
            I => \N__22699\
        );

    \I__3048\ : InMux
    port map (
            O => \N__22737\,
            I => \N__22699\
        );

    \I__3047\ : InMux
    port map (
            O => \N__22736\,
            I => \N__22699\
        );

    \I__3046\ : InMux
    port map (
            O => \N__22735\,
            I => \N__22699\
        );

    \I__3045\ : InMux
    port map (
            O => \N__22734\,
            I => \N__22699\
        );

    \I__3044\ : InMux
    port map (
            O => \N__22733\,
            I => \N__22699\
        );

    \I__3043\ : InMux
    port map (
            O => \N__22732\,
            I => \N__22699\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__22727\,
            I => \N__22696\
        );

    \I__3041\ : InMux
    port map (
            O => \N__22726\,
            I => \N__22691\
        );

    \I__3040\ : InMux
    port map (
            O => \N__22725\,
            I => \N__22691\
        );

    \I__3039\ : InMux
    port map (
            O => \N__22724\,
            I => \N__22669\
        );

    \I__3038\ : InMux
    port map (
            O => \N__22723\,
            I => \N__22669\
        );

    \I__3037\ : InMux
    port map (
            O => \N__22722\,
            I => \N__22669\
        );

    \I__3036\ : InMux
    port map (
            O => \N__22721\,
            I => \N__22669\
        );

    \I__3035\ : InMux
    port map (
            O => \N__22720\,
            I => \N__22669\
        );

    \I__3034\ : InMux
    port map (
            O => \N__22719\,
            I => \N__22669\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__22714\,
            I => \N__22666\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__22699\,
            I => \N__22663\
        );

    \I__3031\ : Span4Mux_v
    port map (
            O => \N__22696\,
            I => \N__22658\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__22691\,
            I => \N__22658\
        );

    \I__3029\ : InMux
    port map (
            O => \N__22690\,
            I => \N__22653\
        );

    \I__3028\ : InMux
    port map (
            O => \N__22689\,
            I => \N__22653\
        );

    \I__3027\ : InMux
    port map (
            O => \N__22688\,
            I => \N__22638\
        );

    \I__3026\ : InMux
    port map (
            O => \N__22687\,
            I => \N__22638\
        );

    \I__3025\ : InMux
    port map (
            O => \N__22686\,
            I => \N__22638\
        );

    \I__3024\ : InMux
    port map (
            O => \N__22685\,
            I => \N__22638\
        );

    \I__3023\ : InMux
    port map (
            O => \N__22684\,
            I => \N__22638\
        );

    \I__3022\ : InMux
    port map (
            O => \N__22683\,
            I => \N__22638\
        );

    \I__3021\ : InMux
    port map (
            O => \N__22682\,
            I => \N__22638\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__22669\,
            I => \current_shift_inst.PI_CTRL.N_76\
        );

    \I__3019\ : Odrv4
    port map (
            O => \N__22666\,
            I => \current_shift_inst.PI_CTRL.N_76\
        );

    \I__3018\ : Odrv4
    port map (
            O => \N__22663\,
            I => \current_shift_inst.PI_CTRL.N_76\
        );

    \I__3017\ : Odrv4
    port map (
            O => \N__22658\,
            I => \current_shift_inst.PI_CTRL.N_76\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__22653\,
            I => \current_shift_inst.PI_CTRL.N_76\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__22638\,
            I => \current_shift_inst.PI_CTRL.N_76\
        );

    \I__3014\ : CascadeMux
    port map (
            O => \N__22625\,
            I => \N__22616\
        );

    \I__3013\ : CascadeMux
    port map (
            O => \N__22624\,
            I => \N__22605\
        );

    \I__3012\ : CascadeMux
    port map (
            O => \N__22623\,
            I => \N__22601\
        );

    \I__3011\ : CascadeMux
    port map (
            O => \N__22622\,
            I => \N__22598\
        );

    \I__3010\ : CascadeMux
    port map (
            O => \N__22621\,
            I => \N__22595\
        );

    \I__3009\ : CascadeMux
    port map (
            O => \N__22620\,
            I => \N__22592\
        );

    \I__3008\ : InMux
    port map (
            O => \N__22619\,
            I => \N__22584\
        );

    \I__3007\ : InMux
    port map (
            O => \N__22616\,
            I => \N__22584\
        );

    \I__3006\ : InMux
    port map (
            O => \N__22615\,
            I => \N__22581\
        );

    \I__3005\ : InMux
    port map (
            O => \N__22614\,
            I => \N__22578\
        );

    \I__3004\ : CascadeMux
    port map (
            O => \N__22613\,
            I => \N__22571\
        );

    \I__3003\ : CascadeMux
    port map (
            O => \N__22612\,
            I => \N__22568\
        );

    \I__3002\ : CascadeMux
    port map (
            O => \N__22611\,
            I => \N__22565\
        );

    \I__3001\ : CascadeMux
    port map (
            O => \N__22610\,
            I => \N__22562\
        );

    \I__3000\ : CascadeMux
    port map (
            O => \N__22609\,
            I => \N__22559\
        );

    \I__2999\ : CascadeMux
    port map (
            O => \N__22608\,
            I => \N__22556\
        );

    \I__2998\ : InMux
    port map (
            O => \N__22605\,
            I => \N__22546\
        );

    \I__2997\ : InMux
    port map (
            O => \N__22604\,
            I => \N__22546\
        );

    \I__2996\ : InMux
    port map (
            O => \N__22601\,
            I => \N__22531\
        );

    \I__2995\ : InMux
    port map (
            O => \N__22598\,
            I => \N__22531\
        );

    \I__2994\ : InMux
    port map (
            O => \N__22595\,
            I => \N__22531\
        );

    \I__2993\ : InMux
    port map (
            O => \N__22592\,
            I => \N__22531\
        );

    \I__2992\ : InMux
    port map (
            O => \N__22591\,
            I => \N__22531\
        );

    \I__2991\ : InMux
    port map (
            O => \N__22590\,
            I => \N__22531\
        );

    \I__2990\ : InMux
    port map (
            O => \N__22589\,
            I => \N__22531\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__22584\,
            I => \N__22528\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__22581\,
            I => \N__22523\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__22578\,
            I => \N__22523\
        );

    \I__2986\ : InMux
    port map (
            O => \N__22577\,
            I => \N__22510\
        );

    \I__2985\ : InMux
    port map (
            O => \N__22576\,
            I => \N__22510\
        );

    \I__2984\ : InMux
    port map (
            O => \N__22575\,
            I => \N__22510\
        );

    \I__2983\ : InMux
    port map (
            O => \N__22574\,
            I => \N__22510\
        );

    \I__2982\ : InMux
    port map (
            O => \N__22571\,
            I => \N__22510\
        );

    \I__2981\ : InMux
    port map (
            O => \N__22568\,
            I => \N__22510\
        );

    \I__2980\ : InMux
    port map (
            O => \N__22565\,
            I => \N__22495\
        );

    \I__2979\ : InMux
    port map (
            O => \N__22562\,
            I => \N__22495\
        );

    \I__2978\ : InMux
    port map (
            O => \N__22559\,
            I => \N__22495\
        );

    \I__2977\ : InMux
    port map (
            O => \N__22556\,
            I => \N__22495\
        );

    \I__2976\ : InMux
    port map (
            O => \N__22555\,
            I => \N__22495\
        );

    \I__2975\ : InMux
    port map (
            O => \N__22554\,
            I => \N__22495\
        );

    \I__2974\ : InMux
    port map (
            O => \N__22553\,
            I => \N__22495\
        );

    \I__2973\ : InMux
    port map (
            O => \N__22552\,
            I => \N__22490\
        );

    \I__2972\ : InMux
    port map (
            O => \N__22551\,
            I => \N__22490\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__22546\,
            I => \N__22487\
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__22531\,
            I => \N__22484\
        );

    \I__2969\ : Span4Mux_h
    port map (
            O => \N__22528\,
            I => \N__22479\
        );

    \I__2968\ : Span4Mux_v
    port map (
            O => \N__22523\,
            I => \N__22479\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__22510\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__22495\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__22490\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__2964\ : Odrv4
    port map (
            O => \N__22487\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__2963\ : Odrv4
    port map (
            O => \N__22484\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__2962\ : Odrv4
    port map (
            O => \N__22479\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__2961\ : CascadeMux
    port map (
            O => \N__22466\,
            I => \N__22462\
        );

    \I__2960\ : CascadeMux
    port map (
            O => \N__22465\,
            I => \N__22459\
        );

    \I__2959\ : InMux
    port map (
            O => \N__22462\,
            I => \N__22456\
        );

    \I__2958\ : InMux
    port map (
            O => \N__22459\,
            I => \N__22453\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__22456\,
            I => \current_shift_inst.PI_CTRL.N_47_16\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__22453\,
            I => \current_shift_inst.PI_CTRL.N_47_16\
        );

    \I__2955\ : InMux
    port map (
            O => \N__22448\,
            I => \N__22444\
        );

    \I__2954\ : InMux
    port map (
            O => \N__22447\,
            I => \N__22441\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__22444\,
            I => \N__22436\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__22441\,
            I => \N__22436\
        );

    \I__2951\ : Odrv4
    port map (
            O => \N__22436\,
            I => \current_shift_inst.PI_CTRL.N_46_16\
        );

    \I__2950\ : InMux
    port map (
            O => \N__22433\,
            I => \N__22430\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__22430\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_16\
        );

    \I__2948\ : InMux
    port map (
            O => \N__22427\,
            I => \N__22424\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__22424\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_17\
        );

    \I__2946\ : InMux
    port map (
            O => \N__22421\,
            I => \N__22418\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__22418\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_18\
        );

    \I__2944\ : InMux
    port map (
            O => \N__22415\,
            I => \N__22412\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__22412\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_19\
        );

    \I__2942\ : InMux
    port map (
            O => \N__22409\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__2941\ : InMux
    port map (
            O => \N__22406\,
            I => \N__22403\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__22403\,
            I => \current_shift_inst.PI_CTRL.un1_enablelt3_0\
        );

    \I__2939\ : CascadeMux
    port map (
            O => \N__22400\,
            I => \N__22397\
        );

    \I__2938\ : InMux
    port map (
            O => \N__22397\,
            I => \N__22394\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__22394\,
            I => \N__22391\
        );

    \I__2936\ : Odrv4
    port map (
            O => \N__22391\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\
        );

    \I__2935\ : InMux
    port map (
            O => \N__22388\,
            I => \N__22385\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__22385\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\
        );

    \I__2933\ : InMux
    port map (
            O => \N__22382\,
            I => \N__22379\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__22379\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\
        );

    \I__2931\ : InMux
    port map (
            O => \N__22376\,
            I => \N__22373\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__22373\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\
        );

    \I__2929\ : InMux
    port map (
            O => \N__22370\,
            I => \N__22367\
        );

    \I__2928\ : LocalMux
    port map (
            O => \N__22367\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\
        );

    \I__2927\ : InMux
    port map (
            O => \N__22364\,
            I => \N__22361\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__22361\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\
        );

    \I__2925\ : InMux
    port map (
            O => \N__22358\,
            I => \N__22355\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__22355\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\
        );

    \I__2923\ : InMux
    port map (
            O => \N__22352\,
            I => \N__22349\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__22349\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\
        );

    \I__2921\ : InMux
    port map (
            O => \N__22346\,
            I => \N__22343\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__22343\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\
        );

    \I__2919\ : CascadeMux
    port map (
            O => \N__22340\,
            I => \N__22337\
        );

    \I__2918\ : InMux
    port map (
            O => \N__22337\,
            I => \N__22334\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__22334\,
            I => \N__22331\
        );

    \I__2916\ : Span4Mux_h
    port map (
            O => \N__22331\,
            I => \N__22328\
        );

    \I__2915\ : Span4Mux_h
    port map (
            O => \N__22328\,
            I => \N__22325\
        );

    \I__2914\ : Odrv4
    port map (
            O => \N__22325\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\
        );

    \I__2913\ : InMux
    port map (
            O => \N__22322\,
            I => \N__22319\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__22319\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\
        );

    \I__2911\ : CascadeMux
    port map (
            O => \N__22316\,
            I => \N__22313\
        );

    \I__2910\ : InMux
    port map (
            O => \N__22313\,
            I => \N__22310\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__22310\,
            I => \N__22307\
        );

    \I__2908\ : Span4Mux_v
    port map (
            O => \N__22307\,
            I => \N__22304\
        );

    \I__2907\ : Span4Mux_h
    port map (
            O => \N__22304\,
            I => \N__22301\
        );

    \I__2906\ : Odrv4
    port map (
            O => \N__22301\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\
        );

    \I__2905\ : InMux
    port map (
            O => \N__22298\,
            I => \N__22295\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__22295\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\
        );

    \I__2903\ : CascadeMux
    port map (
            O => \N__22292\,
            I => \N__22289\
        );

    \I__2902\ : InMux
    port map (
            O => \N__22289\,
            I => \N__22286\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__22286\,
            I => \N__22283\
        );

    \I__2900\ : Span4Mux_h
    port map (
            O => \N__22283\,
            I => \N__22280\
        );

    \I__2899\ : Span4Mux_h
    port map (
            O => \N__22280\,
            I => \N__22277\
        );

    \I__2898\ : Odrv4
    port map (
            O => \N__22277\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\
        );

    \I__2897\ : InMux
    port map (
            O => \N__22274\,
            I => \N__22271\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__22271\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\
        );

    \I__2895\ : InMux
    port map (
            O => \N__22268\,
            I => \N__22265\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__22265\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\
        );

    \I__2893\ : InMux
    port map (
            O => \N__22262\,
            I => \N__22259\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__22259\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\
        );

    \I__2891\ : CascadeMux
    port map (
            O => \N__22256\,
            I => \N__22253\
        );

    \I__2890\ : InMux
    port map (
            O => \N__22253\,
            I => \N__22250\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__22250\,
            I => \N__22247\
        );

    \I__2888\ : Span4Mux_h
    port map (
            O => \N__22247\,
            I => \N__22244\
        );

    \I__2887\ : Span4Mux_h
    port map (
            O => \N__22244\,
            I => \N__22241\
        );

    \I__2886\ : Odrv4
    port map (
            O => \N__22241\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ1Z_6\
        );

    \I__2885\ : InMux
    port map (
            O => \N__22238\,
            I => \N__22235\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__22235\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\
        );

    \I__2883\ : InMux
    port map (
            O => \N__22232\,
            I => \N__22229\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__22229\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\
        );

    \I__2881\ : InMux
    port map (
            O => \N__22226\,
            I => \current_shift_inst.control_input_1_cry_24\
        );

    \I__2880\ : InMux
    port map (
            O => \N__22223\,
            I => \N__22220\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__22220\,
            I => \N__22217\
        );

    \I__2878\ : Span12Mux_h
    port map (
            O => \N__22217\,
            I => \N__22214\
        );

    \I__2877\ : Odrv12
    port map (
            O => \N__22214\,
            I => il_min_comp2_c
        );

    \I__2876\ : InMux
    port map (
            O => \N__22211\,
            I => \N__22208\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__22208\,
            I => \N__22205\
        );

    \I__2874\ : Span4Mux_v
    port map (
            O => \N__22205\,
            I => \N__22202\
        );

    \I__2873\ : Span4Mux_h
    port map (
            O => \N__22202\,
            I => \N__22199\
        );

    \I__2872\ : Odrv4
    port map (
            O => \N__22199\,
            I => il_max_comp2_c
        );

    \I__2871\ : InMux
    port map (
            O => \N__22196\,
            I => \N__22193\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__22193\,
            I => \N__22190\
        );

    \I__2869\ : Span4Mux_v
    port map (
            O => \N__22190\,
            I => \N__22187\
        );

    \I__2868\ : Odrv4
    port map (
            O => \N__22187\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_0\
        );

    \I__2867\ : InMux
    port map (
            O => \N__22184\,
            I => \N__22181\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__22181\,
            I => \N__22178\
        );

    \I__2865\ : Span4Mux_h
    port map (
            O => \N__22178\,
            I => \N__22175\
        );

    \I__2864\ : Odrv4
    port map (
            O => \N__22175\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_6\
        );

    \I__2863\ : InMux
    port map (
            O => \N__22172\,
            I => \N__22169\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__22169\,
            I => \N__22166\
        );

    \I__2861\ : Odrv12
    port map (
            O => \N__22166\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_3\
        );

    \I__2860\ : InMux
    port map (
            O => \N__22163\,
            I => \N__22160\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__22160\,
            I => \N__22157\
        );

    \I__2858\ : Odrv12
    port map (
            O => \N__22157\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_5\
        );

    \I__2857\ : InMux
    port map (
            O => \N__22154\,
            I => \bfn_7_19_0_\
        );

    \I__2856\ : InMux
    port map (
            O => \N__22151\,
            I => \current_shift_inst.control_input_1_cry_16\
        );

    \I__2855\ : InMux
    port map (
            O => \N__22148\,
            I => \current_shift_inst.control_input_1_cry_17\
        );

    \I__2854\ : InMux
    port map (
            O => \N__22145\,
            I => \current_shift_inst.control_input_1_cry_18\
        );

    \I__2853\ : InMux
    port map (
            O => \N__22142\,
            I => \current_shift_inst.control_input_1_cry_19\
        );

    \I__2852\ : InMux
    port map (
            O => \N__22139\,
            I => \current_shift_inst.control_input_1_cry_20\
        );

    \I__2851\ : InMux
    port map (
            O => \N__22136\,
            I => \current_shift_inst.control_input_1_cry_21\
        );

    \I__2850\ : InMux
    port map (
            O => \N__22133\,
            I => \current_shift_inst.control_input_1_cry_22\
        );

    \I__2849\ : InMux
    port map (
            O => \N__22130\,
            I => \bfn_7_20_0_\
        );

    \I__2848\ : InMux
    port map (
            O => \N__22127\,
            I => \current_shift_inst.control_input_1_cry_6\
        );

    \I__2847\ : InMux
    port map (
            O => \N__22124\,
            I => \bfn_7_18_0_\
        );

    \I__2846\ : InMux
    port map (
            O => \N__22121\,
            I => \current_shift_inst.control_input_1_cry_8\
        );

    \I__2845\ : InMux
    port map (
            O => \N__22118\,
            I => \current_shift_inst.control_input_1_cry_9\
        );

    \I__2844\ : InMux
    port map (
            O => \N__22115\,
            I => \current_shift_inst.control_input_1_cry_10\
        );

    \I__2843\ : InMux
    port map (
            O => \N__22112\,
            I => \current_shift_inst.control_input_1_cry_11\
        );

    \I__2842\ : InMux
    port map (
            O => \N__22109\,
            I => \current_shift_inst.control_input_1_cry_12\
        );

    \I__2841\ : InMux
    port map (
            O => \N__22106\,
            I => \current_shift_inst.control_input_1_cry_13\
        );

    \I__2840\ : InMux
    port map (
            O => \N__22103\,
            I => \current_shift_inst.control_input_1_cry_14\
        );

    \I__2839\ : InMux
    port map (
            O => \N__22100\,
            I => \current_shift_inst.control_input_1_cry_0\
        );

    \I__2838\ : InMux
    port map (
            O => \N__22097\,
            I => \current_shift_inst.control_input_1_cry_1\
        );

    \I__2837\ : InMux
    port map (
            O => \N__22094\,
            I => \current_shift_inst.control_input_1_cry_2\
        );

    \I__2836\ : InMux
    port map (
            O => \N__22091\,
            I => \current_shift_inst.control_input_1_cry_3\
        );

    \I__2835\ : InMux
    port map (
            O => \N__22088\,
            I => \current_shift_inst.control_input_1_cry_4\
        );

    \I__2834\ : InMux
    port map (
            O => \N__22085\,
            I => \current_shift_inst.control_input_1_cry_5\
        );

    \I__2833\ : InMux
    port map (
            O => \N__22082\,
            I => \N__22079\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__22079\,
            I => \N__22076\
        );

    \I__2831\ : Odrv4
    port map (
            O => \N__22076\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31\
        );

    \I__2830\ : InMux
    port map (
            O => \N__22073\,
            I => \N__22070\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__22070\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31\
        );

    \I__2828\ : CascadeMux
    port map (
            O => \N__22067\,
            I => \N__22064\
        );

    \I__2827\ : InMux
    port map (
            O => \N__22064\,
            I => \N__22061\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__22061\,
            I => \N__22058\
        );

    \I__2825\ : Span4Mux_v
    port map (
            O => \N__22058\,
            I => \N__22055\
        );

    \I__2824\ : Odrv4
    port map (
            O => \N__22055\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\
        );

    \I__2823\ : CascadeMux
    port map (
            O => \N__22052\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_\
        );

    \I__2822\ : InMux
    port map (
            O => \N__22049\,
            I => \N__22046\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__22046\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_3\
        );

    \I__2820\ : CascadeMux
    port map (
            O => \N__22043\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_2_cascade_\
        );

    \I__2819\ : InMux
    port map (
            O => \N__22040\,
            I => \N__22037\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__22037\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_2\
        );

    \I__2817\ : InMux
    port map (
            O => \N__22034\,
            I => \N__22028\
        );

    \I__2816\ : InMux
    port map (
            O => \N__22033\,
            I => \N__22028\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__22028\,
            I => \N__22025\
        );

    \I__2814\ : Span4Mux_v
    port map (
            O => \N__22025\,
            I => \N__22022\
        );

    \I__2813\ : Odrv4
    port map (
            O => \N__22022\,
            I => \current_shift_inst.PI_CTRL.N_47_21\
        );

    \I__2812\ : InMux
    port map (
            O => \N__22019\,
            I => \N__22015\
        );

    \I__2811\ : InMux
    port map (
            O => \N__22018\,
            I => \N__22012\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__22015\,
            I => \current_shift_inst.PI_CTRL.N_43\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__22012\,
            I => \current_shift_inst.PI_CTRL.N_43\
        );

    \I__2808\ : CascadeMux
    port map (
            O => \N__22007\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31_cascade_\
        );

    \I__2807\ : InMux
    port map (
            O => \N__22004\,
            I => \N__22001\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__22001\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31\
        );

    \I__2805\ : InMux
    port map (
            O => \N__21998\,
            I => \N__21995\
        );

    \I__2804\ : LocalMux
    port map (
            O => \N__21995\,
            I => \current_shift_inst.PI_CTRL.N_46_21\
        );

    \I__2803\ : CascadeMux
    port map (
            O => \N__21992\,
            I => \current_shift_inst.PI_CTRL.N_46_21_cascade_\
        );

    \I__2802\ : InMux
    port map (
            O => \N__21989\,
            I => \N__21985\
        );

    \I__2801\ : InMux
    port map (
            O => \N__21988\,
            I => \N__21982\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__21985\,
            I => \current_shift_inst.PI_CTRL.N_44\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__21982\,
            I => \current_shift_inst.PI_CTRL.N_44\
        );

    \I__2798\ : InMux
    port map (
            O => \N__21977\,
            I => \N__21974\
        );

    \I__2797\ : LocalMux
    port map (
            O => \N__21974\,
            I => \N__21971\
        );

    \I__2796\ : Span4Mux_h
    port map (
            O => \N__21971\,
            I => \N__21968\
        );

    \I__2795\ : Odrv4
    port map (
            O => \N__21968\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_1\
        );

    \I__2794\ : InMux
    port map (
            O => \N__21965\,
            I => \N__21962\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__21962\,
            I => \N__21959\
        );

    \I__2792\ : Odrv4
    port map (
            O => \N__21959\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_4\
        );

    \I__2791\ : InMux
    port map (
            O => \N__21956\,
            I => \N__21953\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__21953\,
            I => \N__21950\
        );

    \I__2789\ : Span4Mux_v
    port map (
            O => \N__21950\,
            I => \N__21947\
        );

    \I__2788\ : Span4Mux_h
    port map (
            O => \N__21947\,
            I => \N__21944\
        );

    \I__2787\ : Odrv4
    port map (
            O => \N__21944\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_9\
        );

    \I__2786\ : CascadeMux
    port map (
            O => \N__21941\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\
        );

    \I__2785\ : InMux
    port map (
            O => \N__21938\,
            I => \N__21935\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__21935\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_18\
        );

    \I__2783\ : CascadeMux
    port map (
            O => \N__21932\,
            I => \N__21929\
        );

    \I__2782\ : InMux
    port map (
            O => \N__21929\,
            I => \N__21926\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__21926\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_23\
        );

    \I__2780\ : CascadeMux
    port map (
            O => \N__21923\,
            I => \N__21920\
        );

    \I__2779\ : InMux
    port map (
            O => \N__21920\,
            I => \N__21917\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__21917\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_22\
        );

    \I__2777\ : InMux
    port map (
            O => \N__21914\,
            I => \N__21911\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__21911\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_24\
        );

    \I__2775\ : CascadeMux
    port map (
            O => \N__21908\,
            I => \N__21901\
        );

    \I__2774\ : CascadeMux
    port map (
            O => \N__21907\,
            I => \N__21897\
        );

    \I__2773\ : CascadeMux
    port map (
            O => \N__21906\,
            I => \N__21893\
        );

    \I__2772\ : InMux
    port map (
            O => \N__21905\,
            I => \N__21878\
        );

    \I__2771\ : InMux
    port map (
            O => \N__21904\,
            I => \N__21878\
        );

    \I__2770\ : InMux
    port map (
            O => \N__21901\,
            I => \N__21878\
        );

    \I__2769\ : InMux
    port map (
            O => \N__21900\,
            I => \N__21878\
        );

    \I__2768\ : InMux
    port map (
            O => \N__21897\,
            I => \N__21878\
        );

    \I__2767\ : InMux
    port map (
            O => \N__21896\,
            I => \N__21878\
        );

    \I__2766\ : InMux
    port map (
            O => \N__21893\,
            I => \N__21878\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__21878\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_25\
        );

    \I__2764\ : InMux
    port map (
            O => \N__21875\,
            I => \N__21872\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__21872\,
            I => \N__21866\
        );

    \I__2762\ : InMux
    port map (
            O => \N__21871\,
            I => \N__21859\
        );

    \I__2761\ : InMux
    port map (
            O => \N__21870\,
            I => \N__21859\
        );

    \I__2760\ : InMux
    port map (
            O => \N__21869\,
            I => \N__21859\
        );

    \I__2759\ : Odrv4
    port map (
            O => \N__21866\,
            I => clk_10khz_i
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__21859\,
            I => clk_10khz_i
        );

    \I__2757\ : InMux
    port map (
            O => \N__21854\,
            I => \N__21851\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__21851\,
            I => \N__21848\
        );

    \I__2755\ : Odrv4
    port map (
            O => \N__21848\,
            I => \clk_10khz_RNIIENAZ0Z2\
        );

    \I__2754\ : InMux
    port map (
            O => \N__21845\,
            I => \N__21842\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__21842\,
            I => \N__21839\
        );

    \I__2752\ : Odrv12
    port map (
            O => \N__21839\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_7\
        );

    \I__2751\ : InMux
    port map (
            O => \N__21836\,
            I => \N__21833\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__21833\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\
        );

    \I__2749\ : InMux
    port map (
            O => \N__21830\,
            I => \N__21827\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__21827\,
            I => \N__21824\
        );

    \I__2747\ : Odrv4
    port map (
            O => \N__21824\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_20\
        );

    \I__2746\ : CascadeMux
    port map (
            O => \N__21821\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_10_31_cascade_\
        );

    \I__2745\ : InMux
    port map (
            O => \N__21818\,
            I => \N__21815\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__21815\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_11_31\
        );

    \I__2743\ : InMux
    port map (
            O => \N__21812\,
            I => \N__21809\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__21809\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_9_31\
        );

    \I__2741\ : InMux
    port map (
            O => \N__21806\,
            I => \N__21803\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__21803\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_8_31\
        );

    \I__2739\ : CascadeMux
    port map (
            O => \N__21800\,
            I => \N__21797\
        );

    \I__2738\ : InMux
    port map (
            O => \N__21797\,
            I => \N__21794\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__21794\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_16\
        );

    \I__2736\ : InMux
    port map (
            O => \N__21791\,
            I => \N__21788\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__21788\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_21\
        );

    \I__2734\ : CascadeMux
    port map (
            O => \N__21785\,
            I => \N__21782\
        );

    \I__2733\ : InMux
    port map (
            O => \N__21782\,
            I => \N__21779\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__21779\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\
        );

    \I__2731\ : CascadeMux
    port map (
            O => \N__21776\,
            I => \N__21773\
        );

    \I__2730\ : InMux
    port map (
            O => \N__21773\,
            I => \N__21770\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__21770\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\
        );

    \I__2728\ : CascadeMux
    port map (
            O => \N__21767\,
            I => \N__21764\
        );

    \I__2727\ : InMux
    port map (
            O => \N__21764\,
            I => \N__21761\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__21761\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\
        );

    \I__2725\ : CascadeMux
    port map (
            O => \N__21758\,
            I => \N__21755\
        );

    \I__2724\ : InMux
    port map (
            O => \N__21755\,
            I => \N__21752\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__21752\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\
        );

    \I__2722\ : InMux
    port map (
            O => \N__21749\,
            I => \N__21746\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__21746\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_15\
        );

    \I__2720\ : CascadeMux
    port map (
            O => \N__21743\,
            I => \N__21740\
        );

    \I__2719\ : InMux
    port map (
            O => \N__21740\,
            I => \N__21737\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__21737\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_19\
        );

    \I__2717\ : CascadeMux
    port map (
            O => \N__21734\,
            I => \N__21731\
        );

    \I__2716\ : InMux
    port map (
            O => \N__21731\,
            I => \N__21728\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__21728\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\
        );

    \I__2714\ : InMux
    port map (
            O => \N__21725\,
            I => \N__21722\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__21722\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\
        );

    \I__2712\ : InMux
    port map (
            O => \N__21719\,
            I => \N__21716\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__21716\,
            I => \N__21708\
        );

    \I__2710\ : InMux
    port map (
            O => \N__21715\,
            I => \N__21705\
        );

    \I__2709\ : InMux
    port map (
            O => \N__21714\,
            I => \N__21702\
        );

    \I__2708\ : InMux
    port map (
            O => \N__21713\,
            I => \N__21697\
        );

    \I__2707\ : InMux
    port map (
            O => \N__21712\,
            I => \N__21697\
        );

    \I__2706\ : InMux
    port map (
            O => \N__21711\,
            I => \N__21694\
        );

    \I__2705\ : Span4Mux_v
    port map (
            O => \N__21708\,
            I => \N__21685\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__21705\,
            I => \N__21685\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__21702\,
            I => \N__21685\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__21697\,
            I => \N__21685\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__21694\,
            I => un2_counter_8
        );

    \I__2700\ : Odrv4
    port map (
            O => \N__21685\,
            I => un2_counter_8
        );

    \I__2699\ : InMux
    port map (
            O => \N__21680\,
            I => \N__21677\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__21677\,
            I => \counter_RNO_0Z0Z_10\
        );

    \I__2697\ : CascadeMux
    port map (
            O => \N__21674\,
            I => \N__21671\
        );

    \I__2696\ : InMux
    port map (
            O => \N__21671\,
            I => \N__21668\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__21668\,
            I => \N__21662\
        );

    \I__2694\ : InMux
    port map (
            O => \N__21667\,
            I => \N__21659\
        );

    \I__2693\ : CascadeMux
    port map (
            O => \N__21666\,
            I => \N__21656\
        );

    \I__2692\ : CascadeMux
    port map (
            O => \N__21665\,
            I => \N__21652\
        );

    \I__2691\ : Span4Mux_h
    port map (
            O => \N__21662\,
            I => \N__21649\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__21659\,
            I => \N__21646\
        );

    \I__2689\ : InMux
    port map (
            O => \N__21656\,
            I => \N__21643\
        );

    \I__2688\ : InMux
    port map (
            O => \N__21655\,
            I => \N__21638\
        );

    \I__2687\ : InMux
    port map (
            O => \N__21652\,
            I => \N__21638\
        );

    \I__2686\ : Odrv4
    port map (
            O => \N__21649\,
            I => un2_counter_9
        );

    \I__2685\ : Odrv4
    port map (
            O => \N__21646\,
            I => un2_counter_9
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__21643\,
            I => un2_counter_9
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__21638\,
            I => un2_counter_9
        );

    \I__2682\ : CascadeMux
    port map (
            O => \N__21629\,
            I => \N__21625\
        );

    \I__2681\ : InMux
    port map (
            O => \N__21628\,
            I => \N__21622\
        );

    \I__2680\ : InMux
    port map (
            O => \N__21625\,
            I => \N__21616\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__21622\,
            I => \N__21613\
        );

    \I__2678\ : InMux
    port map (
            O => \N__21621\,
            I => \N__21608\
        );

    \I__2677\ : InMux
    port map (
            O => \N__21620\,
            I => \N__21608\
        );

    \I__2676\ : InMux
    port map (
            O => \N__21619\,
            I => \N__21605\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__21616\,
            I => \N__21598\
        );

    \I__2674\ : Span4Mux_v
    port map (
            O => \N__21613\,
            I => \N__21598\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__21608\,
            I => \N__21598\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__21605\,
            I => un2_counter_7
        );

    \I__2671\ : Odrv4
    port map (
            O => \N__21598\,
            I => un2_counter_7
        );

    \I__2670\ : InMux
    port map (
            O => \N__21593\,
            I => \N__21589\
        );

    \I__2669\ : InMux
    port map (
            O => \N__21592\,
            I => \N__21586\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__21589\,
            I => \counterZ0Z_10\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__21586\,
            I => \counterZ0Z_10\
        );

    \I__2666\ : InMux
    port map (
            O => \N__21581\,
            I => \N__21578\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__21578\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_8\
        );

    \I__2664\ : CascadeMux
    port map (
            O => \N__21575\,
            I => \N__21572\
        );

    \I__2663\ : InMux
    port map (
            O => \N__21572\,
            I => \N__21569\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__21569\,
            I => \N__21566\
        );

    \I__2661\ : Span4Mux_v
    port map (
            O => \N__21566\,
            I => \N__21563\
        );

    \I__2660\ : Odrv4
    port map (
            O => \N__21563\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\
        );

    \I__2659\ : InMux
    port map (
            O => \N__21560\,
            I => \N__21557\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__21557\,
            I => \N__21554\
        );

    \I__2657\ : Odrv4
    port map (
            O => \N__21554\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\
        );

    \I__2656\ : CascadeMux
    port map (
            O => \N__21551\,
            I => \N__21548\
        );

    \I__2655\ : InMux
    port map (
            O => \N__21548\,
            I => \N__21545\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__21545\,
            I => \N__21542\
        );

    \I__2653\ : Odrv4
    port map (
            O => \N__21542\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\
        );

    \I__2652\ : CascadeMux
    port map (
            O => \N__21539\,
            I => \N__21536\
        );

    \I__2651\ : InMux
    port map (
            O => \N__21536\,
            I => \N__21533\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__21533\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\
        );

    \I__2649\ : CascadeMux
    port map (
            O => \N__21530\,
            I => \N__21527\
        );

    \I__2648\ : InMux
    port map (
            O => \N__21527\,
            I => \N__21524\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__21524\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\
        );

    \I__2646\ : CascadeMux
    port map (
            O => \N__21521\,
            I => \N__21518\
        );

    \I__2645\ : InMux
    port map (
            O => \N__21518\,
            I => \N__21515\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__21515\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\
        );

    \I__2643\ : CascadeMux
    port map (
            O => \N__21512\,
            I => \N__21509\
        );

    \I__2642\ : InMux
    port map (
            O => \N__21509\,
            I => \N__21506\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__21506\,
            I => \N__21503\
        );

    \I__2640\ : Span4Mux_v
    port map (
            O => \N__21503\,
            I => \N__21500\
        );

    \I__2639\ : Odrv4
    port map (
            O => \N__21500\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_17\
        );

    \I__2638\ : CascadeMux
    port map (
            O => \N__21497\,
            I => \N__21494\
        );

    \I__2637\ : InMux
    port map (
            O => \N__21494\,
            I => \N__21491\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__21491\,
            I => \N__21488\
        );

    \I__2635\ : Odrv12
    port map (
            O => \N__21488\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\
        );

    \I__2634\ : InMux
    port map (
            O => \N__21485\,
            I => \N__21482\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__21482\,
            I => \counter_RNO_0Z0Z_7\
        );

    \I__2632\ : InMux
    port map (
            O => \N__21479\,
            I => \N__21475\
        );

    \I__2631\ : InMux
    port map (
            O => \N__21478\,
            I => \N__21472\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__21475\,
            I => \counterZ0Z_7\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__21472\,
            I => \counterZ0Z_7\
        );

    \I__2628\ : CascadeMux
    port map (
            O => \N__21467\,
            I => \N__21462\
        );

    \I__2627\ : InMux
    port map (
            O => \N__21466\,
            I => \N__21459\
        );

    \I__2626\ : InMux
    port map (
            O => \N__21465\,
            I => \N__21456\
        );

    \I__2625\ : InMux
    port map (
            O => \N__21462\,
            I => \N__21453\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__21459\,
            I => \N__21448\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__21456\,
            I => \N__21448\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__21453\,
            I => \counterZ0Z_1\
        );

    \I__2621\ : Odrv4
    port map (
            O => \N__21448\,
            I => \counterZ0Z_1\
        );

    \I__2620\ : InMux
    port map (
            O => \N__21443\,
            I => \N__21439\
        );

    \I__2619\ : InMux
    port map (
            O => \N__21442\,
            I => \N__21436\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__21439\,
            I => \counterZ0Z_2\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__21436\,
            I => \counterZ0Z_2\
        );

    \I__2616\ : CascadeMux
    port map (
            O => \N__21431\,
            I => \un2_counter_5_cascade_\
        );

    \I__2615\ : InMux
    port map (
            O => \N__21428\,
            I => \N__21422\
        );

    \I__2614\ : InMux
    port map (
            O => \N__21427\,
            I => \N__21417\
        );

    \I__2613\ : InMux
    port map (
            O => \N__21426\,
            I => \N__21417\
        );

    \I__2612\ : InMux
    port map (
            O => \N__21425\,
            I => \N__21414\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__21422\,
            I => \N__21411\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__21417\,
            I => \counterZ0Z_0\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__21414\,
            I => \counterZ0Z_0\
        );

    \I__2608\ : Odrv4
    port map (
            O => \N__21411\,
            I => \counterZ0Z_0\
        );

    \I__2607\ : CascadeMux
    port map (
            O => \N__21404\,
            I => \un2_counter_9_cascade_\
        );

    \I__2606\ : CascadeMux
    port map (
            O => \N__21401\,
            I => \clk_10khz_RNIIENAZ0Z2_cascade_\
        );

    \I__2605\ : InMux
    port map (
            O => \N__21398\,
            I => \N__21395\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__21395\,
            I => \N__21392\
        );

    \I__2603\ : Odrv4
    port map (
            O => \N__21392\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_2\
        );

    \I__2602\ : InMux
    port map (
            O => \N__21389\,
            I => \N__21385\
        );

    \I__2601\ : InMux
    port map (
            O => \N__21388\,
            I => \N__21382\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__21385\,
            I => \N__21377\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__21382\,
            I => \N__21377\
        );

    \I__2598\ : Odrv4
    port map (
            O => \N__21377\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\
        );

    \I__2597\ : InMux
    port map (
            O => \N__21374\,
            I => \bfn_4_16_0_\
        );

    \I__2596\ : InMux
    port map (
            O => \N__21371\,
            I => \N__21365\
        );

    \I__2595\ : InMux
    port map (
            O => \N__21370\,
            I => \N__21365\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__21365\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\
        );

    \I__2593\ : InMux
    port map (
            O => \N__21362\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\
        );

    \I__2592\ : InMux
    port map (
            O => \N__21359\,
            I => \N__21355\
        );

    \I__2591\ : CascadeMux
    port map (
            O => \N__21358\,
            I => \N__21352\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__21355\,
            I => \N__21349\
        );

    \I__2589\ : InMux
    port map (
            O => \N__21352\,
            I => \N__21346\
        );

    \I__2588\ : Span4Mux_v
    port map (
            O => \N__21349\,
            I => \N__21343\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__21346\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\
        );

    \I__2586\ : Odrv4
    port map (
            O => \N__21343\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\
        );

    \I__2585\ : InMux
    port map (
            O => \N__21338\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\
        );

    \I__2584\ : InMux
    port map (
            O => \N__21335\,
            I => \N__21331\
        );

    \I__2583\ : InMux
    port map (
            O => \N__21334\,
            I => \N__21328\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__21331\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__21328\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__2580\ : InMux
    port map (
            O => \N__21323\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\
        );

    \I__2579\ : InMux
    port map (
            O => \N__21320\,
            I => \N__21316\
        );

    \I__2578\ : InMux
    port map (
            O => \N__21319\,
            I => \N__21313\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__21316\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__21313\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__2575\ : InMux
    port map (
            O => \N__21308\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\
        );

    \I__2574\ : InMux
    port map (
            O => \N__21305\,
            I => \N__21301\
        );

    \I__2573\ : InMux
    port map (
            O => \N__21304\,
            I => \N__21298\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__21301\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__21298\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__2570\ : InMux
    port map (
            O => \N__21293\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\
        );

    \I__2569\ : CascadeMux
    port map (
            O => \N__21290\,
            I => \N__21286\
        );

    \I__2568\ : InMux
    port map (
            O => \N__21289\,
            I => \N__21283\
        );

    \I__2567\ : InMux
    port map (
            O => \N__21286\,
            I => \N__21280\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__21283\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__21280\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__2564\ : InMux
    port map (
            O => \N__21275\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\
        );

    \I__2563\ : InMux
    port map (
            O => \N__21272\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\
        );

    \I__2562\ : InMux
    port map (
            O => \N__21269\,
            I => \N__21262\
        );

    \I__2561\ : CascadeMux
    port map (
            O => \N__21268\,
            I => \N__21259\
        );

    \I__2560\ : CascadeMux
    port map (
            O => \N__21267\,
            I => \N__21254\
        );

    \I__2559\ : CascadeMux
    port map (
            O => \N__21266\,
            I => \N__21250\
        );

    \I__2558\ : CascadeMux
    port map (
            O => \N__21265\,
            I => \N__21247\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__21262\,
            I => \N__21242\
        );

    \I__2556\ : InMux
    port map (
            O => \N__21259\,
            I => \N__21237\
        );

    \I__2555\ : InMux
    port map (
            O => \N__21258\,
            I => \N__21237\
        );

    \I__2554\ : InMux
    port map (
            O => \N__21257\,
            I => \N__21226\
        );

    \I__2553\ : InMux
    port map (
            O => \N__21254\,
            I => \N__21226\
        );

    \I__2552\ : InMux
    port map (
            O => \N__21253\,
            I => \N__21226\
        );

    \I__2551\ : InMux
    port map (
            O => \N__21250\,
            I => \N__21226\
        );

    \I__2550\ : InMux
    port map (
            O => \N__21247\,
            I => \N__21226\
        );

    \I__2549\ : InMux
    port map (
            O => \N__21246\,
            I => \N__21223\
        );

    \I__2548\ : InMux
    port map (
            O => \N__21245\,
            I => \N__21220\
        );

    \I__2547\ : Span4Mux_h
    port map (
            O => \N__21242\,
            I => \N__21217\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__21237\,
            I => \N__21214\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__21226\,
            I => \N__21207\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__21223\,
            I => \N__21207\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__21220\,
            I => \N__21207\
        );

    \I__2542\ : Span4Mux_v
    port map (
            O => \N__21217\,
            I => \N__21204\
        );

    \I__2541\ : Span4Mux_v
    port map (
            O => \N__21214\,
            I => \N__21201\
        );

    \I__2540\ : Span12Mux_v
    port map (
            O => \N__21207\,
            I => \N__21198\
        );

    \I__2539\ : Span4Mux_v
    port map (
            O => \N__21204\,
            I => \N__21195\
        );

    \I__2538\ : Span4Mux_v
    port map (
            O => \N__21201\,
            I => \N__21192\
        );

    \I__2537\ : Odrv12
    port map (
            O => \N__21198\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__2536\ : Odrv4
    port map (
            O => \N__21195\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__2535\ : Odrv4
    port map (
            O => \N__21192\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__2534\ : InMux
    port map (
            O => \N__21185\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\
        );

    \I__2533\ : CascadeMux
    port map (
            O => \N__21182\,
            I => \N__21179\
        );

    \I__2532\ : InMux
    port map (
            O => \N__21179\,
            I => \N__21173\
        );

    \I__2531\ : InMux
    port map (
            O => \N__21178\,
            I => \N__21173\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__21173\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__2529\ : InMux
    port map (
            O => \N__21170\,
            I => \bfn_4_15_0_\
        );

    \I__2528\ : InMux
    port map (
            O => \N__21167\,
            I => \N__21161\
        );

    \I__2527\ : InMux
    port map (
            O => \N__21166\,
            I => \N__21161\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__21161\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__2525\ : InMux
    port map (
            O => \N__21158\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\
        );

    \I__2524\ : CascadeMux
    port map (
            O => \N__21155\,
            I => \N__21151\
        );

    \I__2523\ : InMux
    port map (
            O => \N__21154\,
            I => \N__21146\
        );

    \I__2522\ : InMux
    port map (
            O => \N__21151\,
            I => \N__21146\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__21146\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__2520\ : InMux
    port map (
            O => \N__21143\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\
        );

    \I__2519\ : CascadeMux
    port map (
            O => \N__21140\,
            I => \N__21137\
        );

    \I__2518\ : InMux
    port map (
            O => \N__21137\,
            I => \N__21133\
        );

    \I__2517\ : InMux
    port map (
            O => \N__21136\,
            I => \N__21130\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__21133\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__21130\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__2514\ : InMux
    port map (
            O => \N__21125\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\
        );

    \I__2513\ : InMux
    port map (
            O => \N__21122\,
            I => \N__21118\
        );

    \I__2512\ : InMux
    port map (
            O => \N__21121\,
            I => \N__21115\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__21118\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__21115\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__2509\ : InMux
    port map (
            O => \N__21110\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\
        );

    \I__2508\ : InMux
    port map (
            O => \N__21107\,
            I => \N__21101\
        );

    \I__2507\ : InMux
    port map (
            O => \N__21106\,
            I => \N__21101\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__21101\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__2505\ : InMux
    port map (
            O => \N__21098\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\
        );

    \I__2504\ : CascadeMux
    port map (
            O => \N__21095\,
            I => \N__21091\
        );

    \I__2503\ : CascadeMux
    port map (
            O => \N__21094\,
            I => \N__21088\
        );

    \I__2502\ : InMux
    port map (
            O => \N__21091\,
            I => \N__21083\
        );

    \I__2501\ : InMux
    port map (
            O => \N__21088\,
            I => \N__21083\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__21083\,
            I => \N__21080\
        );

    \I__2499\ : Odrv4
    port map (
            O => \N__21080\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__2498\ : InMux
    port map (
            O => \N__21077\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\
        );

    \I__2497\ : InMux
    port map (
            O => \N__21074\,
            I => \N__21068\
        );

    \I__2496\ : InMux
    port map (
            O => \N__21073\,
            I => \N__21068\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__21068\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\
        );

    \I__2494\ : InMux
    port map (
            O => \N__21065\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\
        );

    \I__2493\ : InMux
    port map (
            O => \N__21062\,
            I => \N__21058\
        );

    \I__2492\ : InMux
    port map (
            O => \N__21061\,
            I => \N__21054\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__21058\,
            I => \N__21051\
        );

    \I__2490\ : InMux
    port map (
            O => \N__21057\,
            I => \N__21048\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__21054\,
            I => \N__21045\
        );

    \I__2488\ : Span12Mux_v
    port map (
            O => \N__21051\,
            I => \N__21042\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__21048\,
            I => \N__21037\
        );

    \I__2486\ : Span4Mux_h
    port map (
            O => \N__21045\,
            I => \N__21037\
        );

    \I__2485\ : Odrv12
    port map (
            O => \N__21042\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__2484\ : Odrv4
    port map (
            O => \N__21037\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__2483\ : InMux
    port map (
            O => \N__21032\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\
        );

    \I__2482\ : InMux
    port map (
            O => \N__21029\,
            I => \N__21026\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__21026\,
            I => \N__21021\
        );

    \I__2480\ : CascadeMux
    port map (
            O => \N__21025\,
            I => \N__21018\
        );

    \I__2479\ : InMux
    port map (
            O => \N__21024\,
            I => \N__21015\
        );

    \I__2478\ : Span4Mux_v
    port map (
            O => \N__21021\,
            I => \N__21012\
        );

    \I__2477\ : InMux
    port map (
            O => \N__21018\,
            I => \N__21009\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__21015\,
            I => \N__21006\
        );

    \I__2475\ : Span4Mux_v
    port map (
            O => \N__21012\,
            I => \N__21001\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__21009\,
            I => \N__21001\
        );

    \I__2473\ : Span4Mux_h
    port map (
            O => \N__21006\,
            I => \N__20998\
        );

    \I__2472\ : Span4Mux_h
    port map (
            O => \N__21001\,
            I => \N__20995\
        );

    \I__2471\ : Odrv4
    port map (
            O => \N__20998\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__2470\ : Odrv4
    port map (
            O => \N__20995\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__2469\ : InMux
    port map (
            O => \N__20990\,
            I => \bfn_4_14_0_\
        );

    \I__2468\ : InMux
    port map (
            O => \N__20987\,
            I => \N__20984\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__20984\,
            I => \N__20981\
        );

    \I__2466\ : Span4Mux_v
    port map (
            O => \N__20981\,
            I => \N__20977\
        );

    \I__2465\ : InMux
    port map (
            O => \N__20980\,
            I => \N__20973\
        );

    \I__2464\ : Span4Mux_v
    port map (
            O => \N__20977\,
            I => \N__20970\
        );

    \I__2463\ : InMux
    port map (
            O => \N__20976\,
            I => \N__20967\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__20973\,
            I => \N__20964\
        );

    \I__2461\ : Span4Mux_h
    port map (
            O => \N__20970\,
            I => \N__20961\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__20967\,
            I => \N__20956\
        );

    \I__2459\ : Span4Mux_h
    port map (
            O => \N__20964\,
            I => \N__20956\
        );

    \I__2458\ : Odrv4
    port map (
            O => \N__20961\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__2457\ : Odrv4
    port map (
            O => \N__20956\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__2456\ : InMux
    port map (
            O => \N__20951\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\
        );

    \I__2455\ : InMux
    port map (
            O => \N__20948\,
            I => \N__20942\
        );

    \I__2454\ : InMux
    port map (
            O => \N__20947\,
            I => \N__20942\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__20942\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\
        );

    \I__2452\ : InMux
    port map (
            O => \N__20939\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\
        );

    \I__2451\ : InMux
    port map (
            O => \N__20936\,
            I => \N__20930\
        );

    \I__2450\ : InMux
    port map (
            O => \N__20935\,
            I => \N__20930\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__20930\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\
        );

    \I__2448\ : InMux
    port map (
            O => \N__20927\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\
        );

    \I__2447\ : InMux
    port map (
            O => \N__20924\,
            I => \N__20921\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__20921\,
            I => \N__20917\
        );

    \I__2445\ : InMux
    port map (
            O => \N__20920\,
            I => \N__20914\
        );

    \I__2444\ : Odrv4
    port map (
            O => \N__20917\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__20914\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__2442\ : InMux
    port map (
            O => \N__20909\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\
        );

    \I__2441\ : InMux
    port map (
            O => \N__20906\,
            I => \N__20900\
        );

    \I__2440\ : InMux
    port map (
            O => \N__20905\,
            I => \N__20900\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__20900\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__2438\ : InMux
    port map (
            O => \N__20897\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\
        );

    \I__2437\ : CascadeMux
    port map (
            O => \N__20894\,
            I => \N__20891\
        );

    \I__2436\ : InMux
    port map (
            O => \N__20891\,
            I => \N__20888\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__20888\,
            I => \N__20884\
        );

    \I__2434\ : InMux
    port map (
            O => \N__20887\,
            I => \N__20881\
        );

    \I__2433\ : Odrv4
    port map (
            O => \N__20884\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__20881\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__2431\ : InMux
    port map (
            O => \N__20876\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\
        );

    \I__2430\ : InMux
    port map (
            O => \N__20873\,
            I => \N__20869\
        );

    \I__2429\ : InMux
    port map (
            O => \N__20872\,
            I => \N__20866\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__20869\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__20866\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__2426\ : CascadeMux
    port map (
            O => \N__20861\,
            I => \N__20851\
        );

    \I__2425\ : CascadeMux
    port map (
            O => \N__20860\,
            I => \N__20848\
        );

    \I__2424\ : CascadeMux
    port map (
            O => \N__20859\,
            I => \N__20843\
        );

    \I__2423\ : CascadeMux
    port map (
            O => \N__20858\,
            I => \N__20840\
        );

    \I__2422\ : InMux
    port map (
            O => \N__20857\,
            I => \N__20833\
        );

    \I__2421\ : InMux
    port map (
            O => \N__20856\,
            I => \N__20833\
        );

    \I__2420\ : InMux
    port map (
            O => \N__20855\,
            I => \N__20833\
        );

    \I__2419\ : InMux
    port map (
            O => \N__20854\,
            I => \N__20830\
        );

    \I__2418\ : InMux
    port map (
            O => \N__20851\,
            I => \N__20825\
        );

    \I__2417\ : InMux
    port map (
            O => \N__20848\,
            I => \N__20825\
        );

    \I__2416\ : InMux
    port map (
            O => \N__20847\,
            I => \N__20820\
        );

    \I__2415\ : InMux
    port map (
            O => \N__20846\,
            I => \N__20820\
        );

    \I__2414\ : InMux
    port map (
            O => \N__20843\,
            I => \N__20815\
        );

    \I__2413\ : InMux
    port map (
            O => \N__20840\,
            I => \N__20815\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__20833\,
            I => \N__20812\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__20830\,
            I => \N__20808\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__20825\,
            I => \N__20803\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__20820\,
            I => \N__20803\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__20815\,
            I => \N__20798\
        );

    \I__2407\ : Span4Mux_v
    port map (
            O => \N__20812\,
            I => \N__20798\
        );

    \I__2406\ : InMux
    port map (
            O => \N__20811\,
            I => \N__20795\
        );

    \I__2405\ : Span4Mux_v
    port map (
            O => \N__20808\,
            I => \N__20792\
        );

    \I__2404\ : Span12Mux_h
    port map (
            O => \N__20803\,
            I => \N__20789\
        );

    \I__2403\ : Span4Mux_h
    port map (
            O => \N__20798\,
            I => \N__20784\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__20795\,
            I => \N__20784\
        );

    \I__2401\ : Odrv4
    port map (
            O => \N__20792\,
            I => pwm_duty_input_6
        );

    \I__2400\ : Odrv12
    port map (
            O => \N__20789\,
            I => pwm_duty_input_6
        );

    \I__2399\ : Odrv4
    port map (
            O => \N__20784\,
            I => pwm_duty_input_6
        );

    \I__2398\ : InMux
    port map (
            O => \N__20777\,
            I => \N__20763\
        );

    \I__2397\ : InMux
    port map (
            O => \N__20776\,
            I => \N__20763\
        );

    \I__2396\ : InMux
    port map (
            O => \N__20775\,
            I => \N__20754\
        );

    \I__2395\ : InMux
    port map (
            O => \N__20774\,
            I => \N__20754\
        );

    \I__2394\ : InMux
    port map (
            O => \N__20773\,
            I => \N__20754\
        );

    \I__2393\ : InMux
    port map (
            O => \N__20772\,
            I => \N__20754\
        );

    \I__2392\ : InMux
    port map (
            O => \N__20771\,
            I => \N__20747\
        );

    \I__2391\ : InMux
    port map (
            O => \N__20770\,
            I => \N__20747\
        );

    \I__2390\ : InMux
    port map (
            O => \N__20769\,
            I => \N__20747\
        );

    \I__2389\ : InMux
    port map (
            O => \N__20768\,
            I => \N__20744\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__20763\,
            I => \N__20737\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__20754\,
            I => \N__20737\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__20747\,
            I => \N__20737\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__20744\,
            I => \N__20734\
        );

    \I__2384\ : Span4Mux_v
    port map (
            O => \N__20737\,
            I => \N__20731\
        );

    \I__2383\ : Odrv12
    port map (
            O => \N__20734\,
            I => \N_28_mux\
        );

    \I__2382\ : Odrv4
    port map (
            O => \N__20731\,
            I => \N_28_mux\
        );

    \I__2381\ : CascadeMux
    port map (
            O => \N__20726\,
            I => \N__20716\
        );

    \I__2380\ : CascadeMux
    port map (
            O => \N__20725\,
            I => \N__20713\
        );

    \I__2379\ : CascadeMux
    port map (
            O => \N__20724\,
            I => \N__20709\
        );

    \I__2378\ : CascadeMux
    port map (
            O => \N__20723\,
            I => \N__20706\
        );

    \I__2377\ : CascadeMux
    port map (
            O => \N__20722\,
            I => \N__20703\
        );

    \I__2376\ : InMux
    port map (
            O => \N__20721\,
            I => \N__20697\
        );

    \I__2375\ : InMux
    port map (
            O => \N__20720\,
            I => \N__20697\
        );

    \I__2374\ : InMux
    port map (
            O => \N__20719\,
            I => \N__20688\
        );

    \I__2373\ : InMux
    port map (
            O => \N__20716\,
            I => \N__20688\
        );

    \I__2372\ : InMux
    port map (
            O => \N__20713\,
            I => \N__20688\
        );

    \I__2371\ : InMux
    port map (
            O => \N__20712\,
            I => \N__20688\
        );

    \I__2370\ : InMux
    port map (
            O => \N__20709\,
            I => \N__20685\
        );

    \I__2369\ : InMux
    port map (
            O => \N__20706\,
            I => \N__20680\
        );

    \I__2368\ : InMux
    port map (
            O => \N__20703\,
            I => \N__20680\
        );

    \I__2367\ : InMux
    port map (
            O => \N__20702\,
            I => \N__20677\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__20697\,
            I => \N__20668\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__20688\,
            I => \N__20668\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__20685\,
            I => \N__20668\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__20680\,
            I => \N__20668\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__20677\,
            I => \N__20665\
        );

    \I__2361\ : Span4Mux_v
    port map (
            O => \N__20668\,
            I => \N__20662\
        );

    \I__2360\ : Odrv12
    port map (
            O => \N__20665\,
            I => i8_mux
        );

    \I__2359\ : Odrv4
    port map (
            O => \N__20662\,
            I => i8_mux
        );

    \I__2358\ : InMux
    port map (
            O => \N__20657\,
            I => \N__20654\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__20654\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8\
        );

    \I__2356\ : CascadeMux
    port map (
            O => \N__20651\,
            I => \N__20648\
        );

    \I__2355\ : InMux
    port map (
            O => \N__20648\,
            I => \N__20645\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__20645\,
            I => \N__20642\
        );

    \I__2353\ : Span4Mux_h
    port map (
            O => \N__20642\,
            I => \N__20639\
        );

    \I__2352\ : Span4Mux_v
    port map (
            O => \N__20639\,
            I => \N__20636\
        );

    \I__2351\ : Odrv4
    port map (
            O => \N__20636\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\
        );

    \I__2350\ : InMux
    port map (
            O => \N__20633\,
            I => \N__20630\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__20630\,
            I => \N__20627\
        );

    \I__2348\ : Span4Mux_h
    port map (
            O => \N__20627\,
            I => \N__20624\
        );

    \I__2347\ : Span4Mux_v
    port map (
            O => \N__20624\,
            I => \N__20621\
        );

    \I__2346\ : Odrv4
    port map (
            O => \N__20621\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\
        );

    \I__2345\ : InMux
    port map (
            O => \N__20618\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\
        );

    \I__2344\ : CascadeMux
    port map (
            O => \N__20615\,
            I => \N__20612\
        );

    \I__2343\ : InMux
    port map (
            O => \N__20612\,
            I => \N__20609\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__20609\,
            I => \N__20606\
        );

    \I__2341\ : Span4Mux_v
    port map (
            O => \N__20606\,
            I => \N__20603\
        );

    \I__2340\ : Span4Mux_h
    port map (
            O => \N__20603\,
            I => \N__20600\
        );

    \I__2339\ : Odrv4
    port map (
            O => \N__20600\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\
        );

    \I__2338\ : InMux
    port map (
            O => \N__20597\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\
        );

    \I__2337\ : CascadeMux
    port map (
            O => \N__20594\,
            I => \N__20591\
        );

    \I__2336\ : InMux
    port map (
            O => \N__20591\,
            I => \N__20587\
        );

    \I__2335\ : InMux
    port map (
            O => \N__20590\,
            I => \N__20584\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__20587\,
            I => \N__20580\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__20584\,
            I => \N__20577\
        );

    \I__2332\ : InMux
    port map (
            O => \N__20583\,
            I => \N__20574\
        );

    \I__2331\ : Span4Mux_h
    port map (
            O => \N__20580\,
            I => \N__20569\
        );

    \I__2330\ : Span4Mux_h
    port map (
            O => \N__20577\,
            I => \N__20569\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__20574\,
            I => \N__20566\
        );

    \I__2328\ : Span4Mux_v
    port map (
            O => \N__20569\,
            I => \N__20563\
        );

    \I__2327\ : Span4Mux_v
    port map (
            O => \N__20566\,
            I => \N__20560\
        );

    \I__2326\ : Odrv4
    port map (
            O => \N__20563\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__2325\ : Odrv4
    port map (
            O => \N__20560\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__2324\ : InMux
    port map (
            O => \N__20555\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\
        );

    \I__2323\ : CascadeMux
    port map (
            O => \N__20552\,
            I => \N__20549\
        );

    \I__2322\ : InMux
    port map (
            O => \N__20549\,
            I => \N__20545\
        );

    \I__2321\ : InMux
    port map (
            O => \N__20548\,
            I => \N__20542\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__20545\,
            I => \N__20537\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__20542\,
            I => \N__20534\
        );

    \I__2318\ : InMux
    port map (
            O => \N__20541\,
            I => \N__20531\
        );

    \I__2317\ : InMux
    port map (
            O => \N__20540\,
            I => \N__20528\
        );

    \I__2316\ : Span4Mux_v
    port map (
            O => \N__20537\,
            I => \N__20523\
        );

    \I__2315\ : Span4Mux_v
    port map (
            O => \N__20534\,
            I => \N__20523\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__20531\,
            I => \N__20520\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__20528\,
            I => \N__20517\
        );

    \I__2312\ : Span4Mux_v
    port map (
            O => \N__20523\,
            I => \N__20514\
        );

    \I__2311\ : Span4Mux_v
    port map (
            O => \N__20520\,
            I => \N__20509\
        );

    \I__2310\ : Span4Mux_v
    port map (
            O => \N__20517\,
            I => \N__20509\
        );

    \I__2309\ : Odrv4
    port map (
            O => \N__20514\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__2308\ : Odrv4
    port map (
            O => \N__20509\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__2307\ : InMux
    port map (
            O => \N__20504\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\
        );

    \I__2306\ : InMux
    port map (
            O => \N__20501\,
            I => \N__20498\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__20498\,
            I => \N__20495\
        );

    \I__2304\ : Span4Mux_h
    port map (
            O => \N__20495\,
            I => \N__20490\
        );

    \I__2303\ : InMux
    port map (
            O => \N__20494\,
            I => \N__20487\
        );

    \I__2302\ : InMux
    port map (
            O => \N__20493\,
            I => \N__20484\
        );

    \I__2301\ : Span4Mux_v
    port map (
            O => \N__20490\,
            I => \N__20477\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__20487\,
            I => \N__20477\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__20484\,
            I => \N__20477\
        );

    \I__2298\ : Odrv4
    port map (
            O => \N__20477\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__2297\ : InMux
    port map (
            O => \N__20474\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\
        );

    \I__2296\ : InMux
    port map (
            O => \N__20471\,
            I => \N__20468\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__20468\,
            I => \N__20464\
        );

    \I__2294\ : InMux
    port map (
            O => \N__20467\,
            I => \N__20460\
        );

    \I__2293\ : Span4Mux_h
    port map (
            O => \N__20464\,
            I => \N__20457\
        );

    \I__2292\ : InMux
    port map (
            O => \N__20463\,
            I => \N__20454\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__20460\,
            I => \N__20451\
        );

    \I__2290\ : Sp12to4
    port map (
            O => \N__20457\,
            I => \N__20448\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__20454\,
            I => \N__20443\
        );

    \I__2288\ : Span4Mux_h
    port map (
            O => \N__20451\,
            I => \N__20443\
        );

    \I__2287\ : Odrv12
    port map (
            O => \N__20448\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__2286\ : Odrv4
    port map (
            O => \N__20443\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__2285\ : InMux
    port map (
            O => \N__20438\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\
        );

    \I__2284\ : InMux
    port map (
            O => \N__20435\,
            I => un5_counter_cry_9
        );

    \I__2283\ : InMux
    port map (
            O => \N__20432\,
            I => \N__20428\
        );

    \I__2282\ : InMux
    port map (
            O => \N__20431\,
            I => \N__20425\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__20428\,
            I => \counterZ0Z_11\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__20425\,
            I => \counterZ0Z_11\
        );

    \I__2279\ : InMux
    port map (
            O => \N__20420\,
            I => un5_counter_cry_10
        );

    \I__2278\ : InMux
    port map (
            O => \N__20417\,
            I => \N__20413\
        );

    \I__2277\ : InMux
    port map (
            O => \N__20416\,
            I => \N__20410\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__20413\,
            I => \counterZ0Z_12\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__20410\,
            I => \counterZ0Z_12\
        );

    \I__2274\ : InMux
    port map (
            O => \N__20405\,
            I => un5_counter_cry_11
        );

    \I__2273\ : InMux
    port map (
            O => \N__20402\,
            I => \N__20399\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__20399\,
            I => \counter_RNO_0Z0Z_12\
        );

    \I__2271\ : InMux
    port map (
            O => \N__20396\,
            I => \N__20393\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__20393\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0\
        );

    \I__2269\ : InMux
    port map (
            O => \N__20390\,
            I => \N__20387\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__20387\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4\
        );

    \I__2267\ : InMux
    port map (
            O => \N__20384\,
            I => \N__20381\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__20381\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1\
        );

    \I__2265\ : InMux
    port map (
            O => \N__20378\,
            I => \N__20375\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__20375\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3\
        );

    \I__2263\ : InMux
    port map (
            O => \N__20372\,
            I => \N__20369\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__20369\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6\
        );

    \I__2261\ : InMux
    port map (
            O => \N__20366\,
            I => \N__20363\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__20363\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5\
        );

    \I__2259\ : InMux
    port map (
            O => \N__20360\,
            I => un5_counter_cry_1
        );

    \I__2258\ : InMux
    port map (
            O => \N__20357\,
            I => \N__20353\
        );

    \I__2257\ : InMux
    port map (
            O => \N__20356\,
            I => \N__20350\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__20353\,
            I => \counterZ0Z_3\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__20350\,
            I => \counterZ0Z_3\
        );

    \I__2254\ : InMux
    port map (
            O => \N__20345\,
            I => un5_counter_cry_2
        );

    \I__2253\ : InMux
    port map (
            O => \N__20342\,
            I => \N__20338\
        );

    \I__2252\ : InMux
    port map (
            O => \N__20341\,
            I => \N__20335\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__20338\,
            I => \counterZ0Z_4\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__20335\,
            I => \counterZ0Z_4\
        );

    \I__2249\ : InMux
    port map (
            O => \N__20330\,
            I => un5_counter_cry_3
        );

    \I__2248\ : InMux
    port map (
            O => \N__20327\,
            I => \N__20323\
        );

    \I__2247\ : InMux
    port map (
            O => \N__20326\,
            I => \N__20320\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__20323\,
            I => \counterZ0Z_5\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__20320\,
            I => \counterZ0Z_5\
        );

    \I__2244\ : InMux
    port map (
            O => \N__20315\,
            I => un5_counter_cry_4
        );

    \I__2243\ : CascadeMux
    port map (
            O => \N__20312\,
            I => \N__20308\
        );

    \I__2242\ : InMux
    port map (
            O => \N__20311\,
            I => \N__20305\
        );

    \I__2241\ : InMux
    port map (
            O => \N__20308\,
            I => \N__20302\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__20305\,
            I => \counterZ0Z_6\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__20302\,
            I => \counterZ0Z_6\
        );

    \I__2238\ : InMux
    port map (
            O => \N__20297\,
            I => un5_counter_cry_5
        );

    \I__2237\ : InMux
    port map (
            O => \N__20294\,
            I => un5_counter_cry_6
        );

    \I__2236\ : CascadeMux
    port map (
            O => \N__20291\,
            I => \N__20287\
        );

    \I__2235\ : InMux
    port map (
            O => \N__20290\,
            I => \N__20284\
        );

    \I__2234\ : InMux
    port map (
            O => \N__20287\,
            I => \N__20281\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__20284\,
            I => \counterZ0Z_8\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__20281\,
            I => \counterZ0Z_8\
        );

    \I__2231\ : InMux
    port map (
            O => \N__20276\,
            I => un5_counter_cry_7
        );

    \I__2230\ : InMux
    port map (
            O => \N__20273\,
            I => \N__20269\
        );

    \I__2229\ : InMux
    port map (
            O => \N__20272\,
            I => \N__20266\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__20269\,
            I => \counterZ0Z_9\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__20266\,
            I => \counterZ0Z_9\
        );

    \I__2226\ : InMux
    port map (
            O => \N__20261\,
            I => \bfn_4_8_0_\
        );

    \I__2225\ : InMux
    port map (
            O => \N__20258\,
            I => \N__20255\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__20255\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\
        );

    \I__2223\ : CascadeMux
    port map (
            O => \N__20252\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_\
        );

    \I__2222\ : InMux
    port map (
            O => \N__20249\,
            I => \N__20246\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__20246\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9\
        );

    \I__2220\ : InMux
    port map (
            O => \N__20243\,
            I => \N__20240\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__20240\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\
        );

    \I__2218\ : InMux
    port map (
            O => \N__20237\,
            I => \N__20234\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__20234\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\
        );

    \I__2216\ : CascadeMux
    port map (
            O => \N__20231\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_\
        );

    \I__2215\ : InMux
    port map (
            O => \N__20228\,
            I => \N__20225\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__20225\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\
        );

    \I__2213\ : InMux
    port map (
            O => \N__20222\,
            I => \N__20219\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__20219\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\
        );

    \I__2211\ : InMux
    port map (
            O => \N__20216\,
            I => \N__20213\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__20213\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9\
        );

    \I__2209\ : InMux
    port map (
            O => \N__20210\,
            I => \N__20207\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__20207\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\
        );

    \I__2207\ : InMux
    port map (
            O => \N__20204\,
            I => \N__20201\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__20201\,
            I => \N__20198\
        );

    \I__2205\ : Span4Mux_h
    port map (
            O => \N__20198\,
            I => \N__20194\
        );

    \I__2204\ : InMux
    port map (
            O => \N__20197\,
            I => \N__20191\
        );

    \I__2203\ : Odrv4
    port map (
            O => \N__20194\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__20191\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\
        );

    \I__2201\ : InMux
    port map (
            O => \N__20186\,
            I => \N__20183\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__20183\,
            I => \N__20179\
        );

    \I__2199\ : InMux
    port map (
            O => \N__20182\,
            I => \N__20175\
        );

    \I__2198\ : Span4Mux_h
    port map (
            O => \N__20179\,
            I => \N__20172\
        );

    \I__2197\ : InMux
    port map (
            O => \N__20178\,
            I => \N__20169\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__20175\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_14\
        );

    \I__2195\ : Odrv4
    port map (
            O => \N__20172\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_14\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__20169\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_14\
        );

    \I__2193\ : CascadeMux
    port map (
            O => \N__20162\,
            I => \N__20159\
        );

    \I__2192\ : InMux
    port map (
            O => \N__20159\,
            I => \N__20156\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__20156\,
            I => \N__20153\
        );

    \I__2190\ : Odrv4
    port map (
            O => \N__20153\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO\
        );

    \I__2189\ : CascadeMux
    port map (
            O => \N__20150\,
            I => \N__20146\
        );

    \I__2188\ : InMux
    port map (
            O => \N__20149\,
            I => \N__20143\
        );

    \I__2187\ : InMux
    port map (
            O => \N__20146\,
            I => \N__20140\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__20143\,
            I => \N__20127\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__20140\,
            I => \N__20127\
        );

    \I__2184\ : InMux
    port map (
            O => \N__20139\,
            I => \N__20122\
        );

    \I__2183\ : InMux
    port map (
            O => \N__20138\,
            I => \N__20122\
        );

    \I__2182\ : InMux
    port map (
            O => \N__20137\,
            I => \N__20111\
        );

    \I__2181\ : InMux
    port map (
            O => \N__20136\,
            I => \N__20111\
        );

    \I__2180\ : InMux
    port map (
            O => \N__20135\,
            I => \N__20111\
        );

    \I__2179\ : InMux
    port map (
            O => \N__20134\,
            I => \N__20111\
        );

    \I__2178\ : InMux
    port map (
            O => \N__20133\,
            I => \N__20111\
        );

    \I__2177\ : InMux
    port map (
            O => \N__20132\,
            I => \N__20108\
        );

    \I__2176\ : Span4Mux_v
    port map (
            O => \N__20127\,
            I => \N__20105\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__20122\,
            I => \N__20102\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__20111\,
            I => \N__20098\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__20108\,
            I => \N__20095\
        );

    \I__2172\ : Span4Mux_v
    port map (
            O => \N__20105\,
            I => \N__20091\
        );

    \I__2171\ : Span4Mux_h
    port map (
            O => \N__20102\,
            I => \N__20088\
        );

    \I__2170\ : InMux
    port map (
            O => \N__20101\,
            I => \N__20085\
        );

    \I__2169\ : Span4Mux_v
    port map (
            O => \N__20098\,
            I => \N__20080\
        );

    \I__2168\ : Span4Mux_v
    port map (
            O => \N__20095\,
            I => \N__20080\
        );

    \I__2167\ : InMux
    port map (
            O => \N__20094\,
            I => \N__20077\
        );

    \I__2166\ : Odrv4
    port map (
            O => \N__20091\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2165\ : Odrv4
    port map (
            O => \N__20088\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__20085\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2163\ : Odrv4
    port map (
            O => \N__20080\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__20077\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2161\ : InMux
    port map (
            O => \N__20066\,
            I => \N__20063\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__20063\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_4\
        );

    \I__2159\ : CascadeMux
    port map (
            O => \N__20060\,
            I => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\
        );

    \I__2158\ : InMux
    port map (
            O => \N__20057\,
            I => \N__20052\
        );

    \I__2157\ : InMux
    port map (
            O => \N__20056\,
            I => \N__20049\
        );

    \I__2156\ : InMux
    port map (
            O => \N__20055\,
            I => \N__20046\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__20052\,
            I => \N__20043\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__20049\,
            I => \N__20038\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__20046\,
            I => \N__20038\
        );

    \I__2152\ : Span4Mux_v
    port map (
            O => \N__20043\,
            I => \N__20035\
        );

    \I__2151\ : Span4Mux_v
    port map (
            O => \N__20038\,
            I => \N__20032\
        );

    \I__2150\ : Odrv4
    port map (
            O => \N__20035\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__2149\ : Odrv4
    port map (
            O => \N__20032\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__2148\ : CascadeMux
    port map (
            O => \N__20027\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_9_9_cascade_\
        );

    \I__2147\ : CascadeMux
    port map (
            O => \N__20024\,
            I => \N__20021\
        );

    \I__2146\ : InMux
    port map (
            O => \N__20021\,
            I => \N__20018\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__20018\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\
        );

    \I__2144\ : InMux
    port map (
            O => \N__20015\,
            I => \N__20012\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__20012\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\
        );

    \I__2142\ : CascadeMux
    port map (
            O => \N__20009\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9_cascade_\
        );

    \I__2141\ : InMux
    port map (
            O => \N__20006\,
            I => \N__19997\
        );

    \I__2140\ : InMux
    port map (
            O => \N__20005\,
            I => \N__19986\
        );

    \I__2139\ : InMux
    port map (
            O => \N__20004\,
            I => \N__19986\
        );

    \I__2138\ : InMux
    port map (
            O => \N__20003\,
            I => \N__19986\
        );

    \I__2137\ : InMux
    port map (
            O => \N__20002\,
            I => \N__19986\
        );

    \I__2136\ : InMux
    port map (
            O => \N__20001\,
            I => \N__19986\
        );

    \I__2135\ : InMux
    port map (
            O => \N__20000\,
            I => \N__19983\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__19997\,
            I => \N__19978\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__19986\,
            I => \N__19978\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__19983\,
            I => \N__19975\
        );

    \I__2131\ : Span12Mux_v
    port map (
            O => \N__19978\,
            I => \N__19972\
        );

    \I__2130\ : Span12Mux_s7_v
    port map (
            O => \N__19975\,
            I => \N__19969\
        );

    \I__2129\ : Odrv12
    port map (
            O => \N__19972\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__2128\ : Odrv12
    port map (
            O => \N__19969\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__2127\ : InMux
    port map (
            O => \N__19964\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_3\
        );

    \I__2126\ : InMux
    port map (
            O => \N__19961\,
            I => \N__19958\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__19958\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_5\
        );

    \I__2124\ : InMux
    port map (
            O => \N__19955\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_4\
        );

    \I__2123\ : InMux
    port map (
            O => \N__19952\,
            I => \N__19949\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__19949\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_6\
        );

    \I__2121\ : InMux
    port map (
            O => \N__19946\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_5\
        );

    \I__2120\ : InMux
    port map (
            O => \N__19943\,
            I => \N__19940\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__19940\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_7\
        );

    \I__2118\ : InMux
    port map (
            O => \N__19937\,
            I => \N__19934\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__19934\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7\
        );

    \I__2116\ : InMux
    port map (
            O => \N__19931\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_6\
        );

    \I__2115\ : CascadeMux
    port map (
            O => \N__19928\,
            I => \N__19925\
        );

    \I__2114\ : InMux
    port map (
            O => \N__19925\,
            I => \N__19922\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__19922\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_8\
        );

    \I__2112\ : InMux
    port map (
            O => \N__19919\,
            I => \bfn_3_10_0_\
        );

    \I__2111\ : InMux
    port map (
            O => \N__19916\,
            I => \N__19913\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__19913\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO\
        );

    \I__2109\ : CascadeMux
    port map (
            O => \N__19910\,
            I => \N__19907\
        );

    \I__2108\ : InMux
    port map (
            O => \N__19907\,
            I => \N__19904\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__19904\,
            I => \N__19901\
        );

    \I__2106\ : Odrv12
    port map (
            O => \N__19901\,
            I => \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9\
        );

    \I__2105\ : InMux
    port map (
            O => \N__19898\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_8\
        );

    \I__2104\ : CascadeMux
    port map (
            O => \N__19895\,
            I => \N__19892\
        );

    \I__2103\ : InMux
    port map (
            O => \N__19892\,
            I => \N__19889\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__19889\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9\
        );

    \I__2101\ : InMux
    port map (
            O => \N__19886\,
            I => \N__19883\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__19883\,
            I => \N__19879\
        );

    \I__2099\ : InMux
    port map (
            O => \N__19882\,
            I => \N__19876\
        );

    \I__2098\ : Span4Mux_s3_h
    port map (
            O => \N__19879\,
            I => \N__19873\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__19876\,
            I => \N__19870\
        );

    \I__2096\ : Odrv4
    port map (
            O => \N__19873\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__2095\ : Odrv12
    port map (
            O => \N__19870\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__2094\ : InMux
    port map (
            O => \N__19865\,
            I => \N__19862\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__19862\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4\
        );

    \I__2092\ : CascadeMux
    port map (
            O => \N__19859\,
            I => \un2_counter_7_cascade_\
        );

    \I__2091\ : InMux
    port map (
            O => \N__19856\,
            I => \N__19853\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__19853\,
            I => \N__19850\
        );

    \I__2089\ : Span4Mux_h
    port map (
            O => \N__19850\,
            I => \N__19847\
        );

    \I__2088\ : Odrv4
    port map (
            O => \N__19847\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_0\
        );

    \I__2087\ : CascadeMux
    port map (
            O => \N__19844\,
            I => \N__19841\
        );

    \I__2086\ : InMux
    port map (
            O => \N__19841\,
            I => \N__19838\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__19838\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_1\
        );

    \I__2084\ : InMux
    port map (
            O => \N__19835\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_0\
        );

    \I__2083\ : InMux
    port map (
            O => \N__19832\,
            I => \N__19829\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__19829\,
            I => \N__19826\
        );

    \I__2081\ : Span4Mux_v
    port map (
            O => \N__19826\,
            I => \N__19823\
        );

    \I__2080\ : Odrv4
    port map (
            O => \N__19823\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_2\
        );

    \I__2079\ : InMux
    port map (
            O => \N__19820\,
            I => \N__19817\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__19817\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2\
        );

    \I__2077\ : InMux
    port map (
            O => \N__19814\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_1\
        );

    \I__2076\ : InMux
    port map (
            O => \N__19811\,
            I => \N__19808\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__19808\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_3\
        );

    \I__2074\ : InMux
    port map (
            O => \N__19805\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_2\
        );

    \I__2073\ : InMux
    port map (
            O => \N__19802\,
            I => \N__19799\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__19799\,
            I => \N__19796\
        );

    \I__2071\ : Span4Mux_v
    port map (
            O => \N__19796\,
            I => \N__19792\
        );

    \I__2070\ : InMux
    port map (
            O => \N__19795\,
            I => \N__19789\
        );

    \I__2069\ : Odrv4
    port map (
            O => \N__19792\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__19789\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\
        );

    \I__2067\ : InMux
    port map (
            O => \N__19784\,
            I => \N__19781\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__19781\,
            I => \N__19776\
        );

    \I__2065\ : CascadeMux
    port map (
            O => \N__19780\,
            I => \N__19773\
        );

    \I__2064\ : InMux
    port map (
            O => \N__19779\,
            I => \N__19770\
        );

    \I__2063\ : Span4Mux_v
    port map (
            O => \N__19776\,
            I => \N__19767\
        );

    \I__2062\ : InMux
    port map (
            O => \N__19773\,
            I => \N__19764\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__19770\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_12\
        );

    \I__2060\ : Odrv4
    port map (
            O => \N__19767\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_12\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__19764\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_12\
        );

    \I__2058\ : CascadeMux
    port map (
            O => \N__19757\,
            I => \N__19754\
        );

    \I__2057\ : InMux
    port map (
            O => \N__19754\,
            I => \N__19751\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__19751\,
            I => \N__19748\
        );

    \I__2055\ : Span4Mux_v
    port map (
            O => \N__19748\,
            I => \N__19745\
        );

    \I__2054\ : Odrv4
    port map (
            O => \N__19745\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO\
        );

    \I__2053\ : CascadeMux
    port map (
            O => \N__19742\,
            I => \current_shift_inst.PI_CTRL.N_98_cascade_\
        );

    \I__2052\ : InMux
    port map (
            O => \N__19739\,
            I => \N__19727\
        );

    \I__2051\ : InMux
    port map (
            O => \N__19738\,
            I => \N__19727\
        );

    \I__2050\ : InMux
    port map (
            O => \N__19737\,
            I => \N__19727\
        );

    \I__2049\ : InMux
    port map (
            O => \N__19736\,
            I => \N__19727\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__19727\,
            I => \N__19723\
        );

    \I__2047\ : InMux
    port map (
            O => \N__19726\,
            I => \N__19720\
        );

    \I__2046\ : Odrv4
    port map (
            O => \N__19723\,
            I => \current_shift_inst.PI_CTRL.N_96\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__19720\,
            I => \current_shift_inst.PI_CTRL.N_96\
        );

    \I__2044\ : CascadeMux
    port map (
            O => \N__19715\,
            I => \N__19709\
        );

    \I__2043\ : CascadeMux
    port map (
            O => \N__19714\,
            I => \N__19705\
        );

    \I__2042\ : InMux
    port map (
            O => \N__19713\,
            I => \N__19700\
        );

    \I__2041\ : InMux
    port map (
            O => \N__19712\,
            I => \N__19697\
        );

    \I__2040\ : InMux
    port map (
            O => \N__19709\,
            I => \N__19686\
        );

    \I__2039\ : InMux
    port map (
            O => \N__19708\,
            I => \N__19686\
        );

    \I__2038\ : InMux
    port map (
            O => \N__19705\,
            I => \N__19686\
        );

    \I__2037\ : InMux
    port map (
            O => \N__19704\,
            I => \N__19686\
        );

    \I__2036\ : InMux
    port map (
            O => \N__19703\,
            I => \N__19686\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__19700\,
            I => \N__19682\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__19697\,
            I => \N__19676\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__19686\,
            I => \N__19676\
        );

    \I__2032\ : InMux
    port map (
            O => \N__19685\,
            I => \N__19673\
        );

    \I__2031\ : Span4Mux_v
    port map (
            O => \N__19682\,
            I => \N__19670\
        );

    \I__2030\ : InMux
    port map (
            O => \N__19681\,
            I => \N__19667\
        );

    \I__2029\ : Span4Mux_v
    port map (
            O => \N__19676\,
            I => \N__19662\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__19673\,
            I => \N__19662\
        );

    \I__2027\ : Span4Mux_v
    port map (
            O => \N__19670\,
            I => \N__19659\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__19667\,
            I => \N__19654\
        );

    \I__2025\ : Sp12to4
    port map (
            O => \N__19662\,
            I => \N__19654\
        );

    \I__2024\ : Odrv4
    port map (
            O => \N__19659\,
            I => \current_shift_inst.PI_CTRL.N_178\
        );

    \I__2023\ : Odrv12
    port map (
            O => \N__19654\,
            I => \current_shift_inst.PI_CTRL.N_178\
        );

    \I__2022\ : InMux
    port map (
            O => \N__19649\,
            I => \N__19646\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__19646\,
            I => \N__19643\
        );

    \I__2020\ : Odrv4
    port map (
            O => \N__19643\,
            I => \current_shift_inst.PI_CTRL.N_91\
        );

    \I__2019\ : CascadeMux
    port map (
            O => \N__19640\,
            I => \N__19637\
        );

    \I__2018\ : InMux
    port map (
            O => \N__19637\,
            I => \N__19634\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__19634\,
            I => \N__19631\
        );

    \I__2016\ : Odrv4
    port map (
            O => \N__19631\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO\
        );

    \I__2015\ : CascadeMux
    port map (
            O => \N__19628\,
            I => \N__19624\
        );

    \I__2014\ : InMux
    port map (
            O => \N__19627\,
            I => \N__19621\
        );

    \I__2013\ : InMux
    port map (
            O => \N__19624\,
            I => \N__19618\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__19621\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_18\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__19618\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_18\
        );

    \I__2010\ : InMux
    port map (
            O => \N__19613\,
            I => \N__19610\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__19610\,
            I => \N__19606\
        );

    \I__2008\ : InMux
    port map (
            O => \N__19609\,
            I => \N__19603\
        );

    \I__2007\ : Odrv4
    port map (
            O => \N__19606\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__19603\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\
        );

    \I__2005\ : CascadeMux
    port map (
            O => \N__19598\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_18_cascade_\
        );

    \I__2004\ : InMux
    port map (
            O => \N__19595\,
            I => \N__19592\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__19592\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO\
        );

    \I__2002\ : InMux
    port map (
            O => \N__19589\,
            I => \N__19585\
        );

    \I__2001\ : InMux
    port map (
            O => \N__19588\,
            I => \N__19582\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__19585\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__19582\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\
        );

    \I__1998\ : CascadeMux
    port map (
            O => \N__19577\,
            I => \N__19574\
        );

    \I__1997\ : InMux
    port map (
            O => \N__19574\,
            I => \N__19571\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__19571\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO\
        );

    \I__1995\ : InMux
    port map (
            O => \N__19568\,
            I => \N__19563\
        );

    \I__1994\ : InMux
    port map (
            O => \N__19567\,
            I => \N__19558\
        );

    \I__1993\ : InMux
    port map (
            O => \N__19566\,
            I => \N__19558\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__19563\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_16\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__19558\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_16\
        );

    \I__1990\ : InMux
    port map (
            O => \N__19553\,
            I => \N__19549\
        );

    \I__1989\ : InMux
    port map (
            O => \N__19552\,
            I => \N__19546\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__19549\,
            I => \N__19543\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__19546\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\
        );

    \I__1986\ : Odrv4
    port map (
            O => \N__19543\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\
        );

    \I__1985\ : InMux
    port map (
            O => \N__19538\,
            I => \N__19533\
        );

    \I__1984\ : InMux
    port map (
            O => \N__19537\,
            I => \N__19530\
        );

    \I__1983\ : InMux
    port map (
            O => \N__19536\,
            I => \N__19527\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__19533\,
            I => \N__19522\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__19530\,
            I => \N__19522\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__19527\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_13\
        );

    \I__1979\ : Odrv12
    port map (
            O => \N__19522\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_13\
        );

    \I__1978\ : InMux
    port map (
            O => \N__19517\,
            I => \N__19514\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__19514\,
            I => \N__19511\
        );

    \I__1976\ : Span4Mux_h
    port map (
            O => \N__19511\,
            I => \N__19507\
        );

    \I__1975\ : InMux
    port map (
            O => \N__19510\,
            I => \N__19504\
        );

    \I__1974\ : Span4Mux_v
    port map (
            O => \N__19507\,
            I => \N__19501\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__19504\,
            I => \N__19498\
        );

    \I__1972\ : Odrv4
    port map (
            O => \N__19501\,
            I => \pwm_generator_inst.O_10\
        );

    \I__1971\ : Odrv4
    port map (
            O => \N__19498\,
            I => \pwm_generator_inst.O_10\
        );

    \I__1970\ : InMux
    port map (
            O => \N__19493\,
            I => \N__19490\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__19490\,
            I => \N__19486\
        );

    \I__1968\ : InMux
    port map (
            O => \N__19489\,
            I => \N__19482\
        );

    \I__1967\ : Span4Mux_v
    port map (
            O => \N__19486\,
            I => \N__19479\
        );

    \I__1966\ : InMux
    port map (
            O => \N__19485\,
            I => \N__19476\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__19482\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_10\
        );

    \I__1964\ : Odrv4
    port map (
            O => \N__19479\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_10\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__19476\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_10\
        );

    \I__1962\ : CascadeMux
    port map (
            O => \N__19469\,
            I => \N__19466\
        );

    \I__1961\ : InMux
    port map (
            O => \N__19466\,
            I => \N__19463\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__19463\,
            I => \N__19460\
        );

    \I__1959\ : Span4Mux_v
    port map (
            O => \N__19460\,
            I => \N__19457\
        );

    \I__1958\ : Odrv4
    port map (
            O => \N__19457\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO\
        );

    \I__1957\ : InMux
    port map (
            O => \N__19454\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_16\
        );

    \I__1956\ : InMux
    port map (
            O => \N__19451\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_17\
        );

    \I__1955\ : InMux
    port map (
            O => \N__19448\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_18\
        );

    \I__1954\ : InMux
    port map (
            O => \N__19445\,
            I => \N__19440\
        );

    \I__1953\ : InMux
    port map (
            O => \N__19444\,
            I => \N__19437\
        );

    \I__1952\ : InMux
    port map (
            O => \N__19443\,
            I => \N__19434\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__19440\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_15\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__19437\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_15\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__19434\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_15\
        );

    \I__1948\ : InMux
    port map (
            O => \N__19427\,
            I => \N__19423\
        );

    \I__1947\ : InMux
    port map (
            O => \N__19426\,
            I => \N__19420\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__19423\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__19420\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\
        );

    \I__1944\ : CascadeMux
    port map (
            O => \N__19415\,
            I => \N__19412\
        );

    \I__1943\ : InMux
    port map (
            O => \N__19412\,
            I => \N__19409\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__19409\,
            I => \N__19406\
        );

    \I__1941\ : Odrv4
    port map (
            O => \N__19406\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO\
        );

    \I__1940\ : InMux
    port map (
            O => \N__19403\,
            I => \N__19400\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__19400\,
            I => \N__19396\
        );

    \I__1938\ : InMux
    port map (
            O => \N__19399\,
            I => \N__19393\
        );

    \I__1937\ : Odrv4
    port map (
            O => \N__19396\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_17\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__19393\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_17\
        );

    \I__1935\ : InMux
    port map (
            O => \N__19388\,
            I => \N__19384\
        );

    \I__1934\ : InMux
    port map (
            O => \N__19387\,
            I => \N__19381\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__19384\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__19381\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\
        );

    \I__1931\ : CascadeMux
    port map (
            O => \N__19376\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_\
        );

    \I__1930\ : InMux
    port map (
            O => \N__19373\,
            I => \N__19370\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__19370\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO\
        );

    \I__1928\ : InMux
    port map (
            O => \N__19367\,
            I => \N__19364\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__19364\,
            I => \N__19361\
        );

    \I__1926\ : Span4Mux_h
    port map (
            O => \N__19361\,
            I => \N__19358\
        );

    \I__1925\ : Odrv4
    port map (
            O => \N__19358\,
            I => \pwm_generator_inst.O_8\
        );

    \I__1924\ : InMux
    port map (
            O => \N__19355\,
            I => \N__19352\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__19352\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_8\
        );

    \I__1922\ : InMux
    port map (
            O => \N__19349\,
            I => \N__19346\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__19346\,
            I => \N__19343\
        );

    \I__1920\ : Span4Mux_h
    port map (
            O => \N__19343\,
            I => \N__19340\
        );

    \I__1919\ : Odrv4
    port map (
            O => \N__19340\,
            I => \pwm_generator_inst.O_9\
        );

    \I__1918\ : InMux
    port map (
            O => \N__19337\,
            I => \N__19334\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__19334\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_9\
        );

    \I__1916\ : InMux
    port map (
            O => \N__19331\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_9\
        );

    \I__1915\ : InMux
    port map (
            O => \N__19328\,
            I => \N__19325\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__19325\,
            I => \N__19321\
        );

    \I__1913\ : InMux
    port map (
            O => \N__19324\,
            I => \N__19318\
        );

    \I__1912\ : Span4Mux_v
    port map (
            O => \N__19321\,
            I => \N__19315\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__19318\,
            I => \N__19312\
        );

    \I__1910\ : Odrv4
    port map (
            O => \N__19315\,
            I => \pwm_generator_inst.un3_threshold_acc\
        );

    \I__1909\ : Odrv4
    port map (
            O => \N__19312\,
            I => \pwm_generator_inst.un3_threshold_acc\
        );

    \I__1908\ : InMux
    port map (
            O => \N__19307\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_10\
        );

    \I__1907\ : InMux
    port map (
            O => \N__19304\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_11\
        );

    \I__1906\ : InMux
    port map (
            O => \N__19301\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_12\
        );

    \I__1905\ : InMux
    port map (
            O => \N__19298\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_13\
        );

    \I__1904\ : InMux
    port map (
            O => \N__19295\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_14\
        );

    \I__1903\ : InMux
    port map (
            O => \N__19292\,
            I => \bfn_2_9_0_\
        );

    \I__1902\ : InMux
    port map (
            O => \N__19289\,
            I => \N__19286\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__19286\,
            I => \N__19283\
        );

    \I__1900\ : Span4Mux_h
    port map (
            O => \N__19283\,
            I => \N__19280\
        );

    \I__1899\ : Odrv4
    port map (
            O => \N__19280\,
            I => \pwm_generator_inst.O_0\
        );

    \I__1898\ : InMux
    port map (
            O => \N__19277\,
            I => \N__19274\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__19274\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_0\
        );

    \I__1896\ : InMux
    port map (
            O => \N__19271\,
            I => \N__19268\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__19268\,
            I => \N__19265\
        );

    \I__1894\ : Span4Mux_h
    port map (
            O => \N__19265\,
            I => \N__19262\
        );

    \I__1893\ : Odrv4
    port map (
            O => \N__19262\,
            I => \pwm_generator_inst.O_1\
        );

    \I__1892\ : InMux
    port map (
            O => \N__19259\,
            I => \N__19256\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__19256\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_1\
        );

    \I__1890\ : InMux
    port map (
            O => \N__19253\,
            I => \N__19250\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__19250\,
            I => \N__19247\
        );

    \I__1888\ : Span4Mux_v
    port map (
            O => \N__19247\,
            I => \N__19244\
        );

    \I__1887\ : Odrv4
    port map (
            O => \N__19244\,
            I => \pwm_generator_inst.O_2\
        );

    \I__1886\ : InMux
    port map (
            O => \N__19241\,
            I => \N__19238\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__19238\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_2\
        );

    \I__1884\ : InMux
    port map (
            O => \N__19235\,
            I => \N__19232\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__19232\,
            I => \N__19229\
        );

    \I__1882\ : Span4Mux_v
    port map (
            O => \N__19229\,
            I => \N__19226\
        );

    \I__1881\ : Odrv4
    port map (
            O => \N__19226\,
            I => \pwm_generator_inst.O_3\
        );

    \I__1880\ : InMux
    port map (
            O => \N__19223\,
            I => \N__19220\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__19220\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_3\
        );

    \I__1878\ : InMux
    port map (
            O => \N__19217\,
            I => \N__19214\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__19214\,
            I => \N__19211\
        );

    \I__1876\ : Span4Mux_h
    port map (
            O => \N__19211\,
            I => \N__19208\
        );

    \I__1875\ : Odrv4
    port map (
            O => \N__19208\,
            I => \pwm_generator_inst.O_4\
        );

    \I__1874\ : InMux
    port map (
            O => \N__19205\,
            I => \N__19202\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__19202\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_4\
        );

    \I__1872\ : InMux
    port map (
            O => \N__19199\,
            I => \N__19196\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__19196\,
            I => \N__19193\
        );

    \I__1870\ : Span4Mux_h
    port map (
            O => \N__19193\,
            I => \N__19190\
        );

    \I__1869\ : Odrv4
    port map (
            O => \N__19190\,
            I => \pwm_generator_inst.O_5\
        );

    \I__1868\ : InMux
    port map (
            O => \N__19187\,
            I => \N__19184\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__19184\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_5\
        );

    \I__1866\ : InMux
    port map (
            O => \N__19181\,
            I => \N__19178\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__19178\,
            I => \N__19175\
        );

    \I__1864\ : Span4Mux_h
    port map (
            O => \N__19175\,
            I => \N__19172\
        );

    \I__1863\ : Odrv4
    port map (
            O => \N__19172\,
            I => \pwm_generator_inst.O_6\
        );

    \I__1862\ : InMux
    port map (
            O => \N__19169\,
            I => \N__19166\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__19166\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_6\
        );

    \I__1860\ : InMux
    port map (
            O => \N__19163\,
            I => \N__19160\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__19160\,
            I => \N__19157\
        );

    \I__1858\ : Span4Mux_h
    port map (
            O => \N__19157\,
            I => \N__19154\
        );

    \I__1857\ : Odrv4
    port map (
            O => \N__19154\,
            I => \pwm_generator_inst.O_7\
        );

    \I__1856\ : InMux
    port map (
            O => \N__19151\,
            I => \N__19148\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__19148\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_7\
        );

    \I__1854\ : InMux
    port map (
            O => \N__19145\,
            I => \N__19142\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__19142\,
            I => un7_start_stop
        );

    \I__1852\ : InMux
    port map (
            O => \N__19139\,
            I => \N__19134\
        );

    \I__1851\ : InMux
    port map (
            O => \N__19138\,
            I => \N__19129\
        );

    \I__1850\ : InMux
    port map (
            O => \N__19137\,
            I => \N__19129\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__19134\,
            I => \N__19126\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__19129\,
            I => pwm_duty_input_5
        );

    \I__1847\ : Odrv4
    port map (
            O => \N__19126\,
            I => pwm_duty_input_5
        );

    \I__1846\ : CascadeMux
    port map (
            O => \N__19121\,
            I => \N__19117\
        );

    \I__1845\ : InMux
    port map (
            O => \N__19120\,
            I => \N__19113\
        );

    \I__1844\ : InMux
    port map (
            O => \N__19117\,
            I => \N__19108\
        );

    \I__1843\ : InMux
    port map (
            O => \N__19116\,
            I => \N__19108\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__19113\,
            I => \N__19105\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__19108\,
            I => pwm_duty_input_9
        );

    \I__1840\ : Odrv4
    port map (
            O => \N__19105\,
            I => pwm_duty_input_9
        );

    \I__1839\ : InMux
    port map (
            O => \N__19100\,
            I => \N__19096\
        );

    \I__1838\ : CascadeMux
    port map (
            O => \N__19099\,
            I => \N__19092\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__19096\,
            I => \N__19089\
        );

    \I__1836\ : InMux
    port map (
            O => \N__19095\,
            I => \N__19086\
        );

    \I__1835\ : InMux
    port map (
            O => \N__19092\,
            I => \N__19083\
        );

    \I__1834\ : Span4Mux_v
    port map (
            O => \N__19089\,
            I => \N__19080\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__19086\,
            I => pwm_duty_input_8
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__19083\,
            I => pwm_duty_input_8
        );

    \I__1831\ : Odrv4
    port map (
            O => \N__19080\,
            I => pwm_duty_input_8
        );

    \I__1830\ : CascadeMux
    port map (
            O => \N__19073\,
            I => \N__19070\
        );

    \I__1829\ : InMux
    port map (
            O => \N__19070\,
            I => \N__19067\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__19067\,
            I => \current_shift_inst.PI_CTRL.m7_2\
        );

    \I__1827\ : InMux
    port map (
            O => \N__19064\,
            I => \N__19059\
        );

    \I__1826\ : InMux
    port map (
            O => \N__19063\,
            I => \N__19056\
        );

    \I__1825\ : InMux
    port map (
            O => \N__19062\,
            I => \N__19053\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__19059\,
            I => \N__19050\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__19056\,
            I => pwm_duty_input_7
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__19053\,
            I => pwm_duty_input_7
        );

    \I__1821\ : Odrv4
    port map (
            O => \N__19050\,
            I => pwm_duty_input_7
        );

    \I__1820\ : InMux
    port map (
            O => \N__19043\,
            I => \N__19040\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__19040\,
            I => \N__19037\
        );

    \I__1818\ : Odrv4
    port map (
            O => \N__19037\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\
        );

    \I__1817\ : CascadeMux
    port map (
            O => \N__19034\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3_cascade_\
        );

    \I__1816\ : CascadeMux
    port map (
            O => \N__19031\,
            I => \N__19027\
        );

    \I__1815\ : InMux
    port map (
            O => \N__19030\,
            I => \N__19019\
        );

    \I__1814\ : InMux
    port map (
            O => \N__19027\,
            I => \N__19019\
        );

    \I__1813\ : InMux
    port map (
            O => \N__19026\,
            I => \N__19019\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__19019\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_3\
        );

    \I__1811\ : InMux
    port map (
            O => \N__19016\,
            I => \N__19012\
        );

    \I__1810\ : InMux
    port map (
            O => \N__19015\,
            I => \N__19009\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__19012\,
            I => pwm_duty_input_1
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__19009\,
            I => pwm_duty_input_1
        );

    \I__1807\ : InMux
    port map (
            O => \N__19004\,
            I => \N__18999\
        );

    \I__1806\ : InMux
    port map (
            O => \N__19003\,
            I => \N__18996\
        );

    \I__1805\ : InMux
    port map (
            O => \N__19002\,
            I => \N__18993\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__18999\,
            I => pwm_duty_input_3
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__18996\,
            I => pwm_duty_input_3
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__18993\,
            I => pwm_duty_input_3
        );

    \I__1801\ : CascadeMux
    port map (
            O => \N__18986\,
            I => \N__18983\
        );

    \I__1800\ : InMux
    port map (
            O => \N__18983\,
            I => \N__18979\
        );

    \I__1799\ : InMux
    port map (
            O => \N__18982\,
            I => \N__18976\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__18979\,
            I => pwm_duty_input_0
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__18976\,
            I => pwm_duty_input_0
        );

    \I__1796\ : InMux
    port map (
            O => \N__18971\,
            I => \N__18967\
        );

    \I__1795\ : InMux
    port map (
            O => \N__18970\,
            I => \N__18964\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__18967\,
            I => pwm_duty_input_2
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__18964\,
            I => pwm_duty_input_2
        );

    \I__1792\ : InMux
    port map (
            O => \N__18959\,
            I => \N__18956\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__18956\,
            I => \current_shift_inst.PI_CTRL.m14_2\
        );

    \I__1790\ : InMux
    port map (
            O => \N__18953\,
            I => \N__18932\
        );

    \I__1789\ : InMux
    port map (
            O => \N__18952\,
            I => \N__18932\
        );

    \I__1788\ : InMux
    port map (
            O => \N__18951\,
            I => \N__18915\
        );

    \I__1787\ : InMux
    port map (
            O => \N__18950\,
            I => \N__18915\
        );

    \I__1786\ : InMux
    port map (
            O => \N__18949\,
            I => \N__18915\
        );

    \I__1785\ : InMux
    port map (
            O => \N__18948\,
            I => \N__18915\
        );

    \I__1784\ : InMux
    port map (
            O => \N__18947\,
            I => \N__18915\
        );

    \I__1783\ : InMux
    port map (
            O => \N__18946\,
            I => \N__18915\
        );

    \I__1782\ : InMux
    port map (
            O => \N__18945\,
            I => \N__18915\
        );

    \I__1781\ : InMux
    port map (
            O => \N__18944\,
            I => \N__18915\
        );

    \I__1780\ : InMux
    port map (
            O => \N__18943\,
            I => \N__18900\
        );

    \I__1779\ : InMux
    port map (
            O => \N__18942\,
            I => \N__18900\
        );

    \I__1778\ : InMux
    port map (
            O => \N__18941\,
            I => \N__18900\
        );

    \I__1777\ : InMux
    port map (
            O => \N__18940\,
            I => \N__18900\
        );

    \I__1776\ : InMux
    port map (
            O => \N__18939\,
            I => \N__18900\
        );

    \I__1775\ : InMux
    port map (
            O => \N__18938\,
            I => \N__18900\
        );

    \I__1774\ : InMux
    port map (
            O => \N__18937\,
            I => \N__18900\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__18932\,
            I => \N__18897\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__18915\,
            I => \N__18892\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__18900\,
            I => \N__18892\
        );

    \I__1770\ : Span4Mux_h
    port map (
            O => \N__18897\,
            I => \N__18880\
        );

    \I__1769\ : Span4Mux_v
    port map (
            O => \N__18892\,
            I => \N__18880\
        );

    \I__1768\ : InMux
    port map (
            O => \N__18891\,
            I => \N__18875\
        );

    \I__1767\ : InMux
    port map (
            O => \N__18890\,
            I => \N__18875\
        );

    \I__1766\ : InMux
    port map (
            O => \N__18889\,
            I => \N__18868\
        );

    \I__1765\ : InMux
    port map (
            O => \N__18888\,
            I => \N__18868\
        );

    \I__1764\ : InMux
    port map (
            O => \N__18887\,
            I => \N__18868\
        );

    \I__1763\ : InMux
    port map (
            O => \N__18886\,
            I => \N__18863\
        );

    \I__1762\ : InMux
    port map (
            O => \N__18885\,
            I => \N__18863\
        );

    \I__1761\ : Span4Mux_v
    port map (
            O => \N__18880\,
            I => \N__18856\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__18875\,
            I => \N__18856\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__18868\,
            I => \N__18856\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__18863\,
            I => pwm_duty_input_10
        );

    \I__1757\ : Odrv4
    port map (
            O => \N__18856\,
            I => pwm_duty_input_10
        );

    \I__1756\ : CascadeMux
    port map (
            O => \N__18851\,
            I => \current_shift_inst.PI_CTRL.N_19_cascade_\
        );

    \I__1755\ : InMux
    port map (
            O => \N__18848\,
            I => \N__18843\
        );

    \I__1754\ : InMux
    port map (
            O => \N__18847\,
            I => \N__18840\
        );

    \I__1753\ : InMux
    port map (
            O => \N__18846\,
            I => \N__18837\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__18843\,
            I => pwm_duty_input_4
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__18840\,
            I => pwm_duty_input_4
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__18837\,
            I => pwm_duty_input_4
        );

    \I__1749\ : CascadeMux
    port map (
            O => \N__18830\,
            I => \N__18827\
        );

    \I__1748\ : InMux
    port map (
            O => \N__18827\,
            I => \N__18824\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__18824\,
            I => \N__18821\
        );

    \I__1746\ : Span4Mux_v
    port map (
            O => \N__18821\,
            I => \N__18818\
        );

    \I__1745\ : Odrv4
    port map (
            O => \N__18818\,
            I => \pwm_generator_inst.un2_threshold_acc_2_10\
        );

    \I__1744\ : InMux
    port map (
            O => \N__18815\,
            I => \N__18812\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__18812\,
            I => \N__18809\
        );

    \I__1742\ : Odrv4
    port map (
            O => \N__18809\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0\
        );

    \I__1741\ : InMux
    port map (
            O => \N__18806\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\
        );

    \I__1740\ : InMux
    port map (
            O => \N__18803\,
            I => \N__18800\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__18800\,
            I => \N__18797\
        );

    \I__1738\ : Span4Mux_v
    port map (
            O => \N__18797\,
            I => \N__18794\
        );

    \I__1737\ : Odrv4
    port map (
            O => \N__18794\,
            I => \pwm_generator_inst.un2_threshold_acc_2_11\
        );

    \I__1736\ : CascadeMux
    port map (
            O => \N__18791\,
            I => \N__18788\
        );

    \I__1735\ : InMux
    port map (
            O => \N__18788\,
            I => \N__18785\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__18785\,
            I => \N__18782\
        );

    \I__1733\ : Odrv4
    port map (
            O => \N__18782\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0\
        );

    \I__1732\ : InMux
    port map (
            O => \N__18779\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\
        );

    \I__1731\ : CascadeMux
    port map (
            O => \N__18776\,
            I => \N__18773\
        );

    \I__1730\ : InMux
    port map (
            O => \N__18773\,
            I => \N__18770\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__18770\,
            I => \N__18767\
        );

    \I__1728\ : Span4Mux_h
    port map (
            O => \N__18767\,
            I => \N__18764\
        );

    \I__1727\ : Odrv4
    port map (
            O => \N__18764\,
            I => \pwm_generator_inst.un2_threshold_acc_2_12\
        );

    \I__1726\ : InMux
    port map (
            O => \N__18761\,
            I => \N__18758\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__18758\,
            I => \N__18755\
        );

    \I__1724\ : Odrv4
    port map (
            O => \N__18755\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0\
        );

    \I__1723\ : InMux
    port map (
            O => \N__18752\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\
        );

    \I__1722\ : InMux
    port map (
            O => \N__18749\,
            I => \N__18746\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__18746\,
            I => \N__18743\
        );

    \I__1720\ : Span4Mux_v
    port map (
            O => \N__18743\,
            I => \N__18740\
        );

    \I__1719\ : Odrv4
    port map (
            O => \N__18740\,
            I => \pwm_generator_inst.un2_threshold_acc_2_13\
        );

    \I__1718\ : InMux
    port map (
            O => \N__18737\,
            I => \N__18734\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__18734\,
            I => \N__18731\
        );

    \I__1716\ : Odrv4
    port map (
            O => \N__18731\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0\
        );

    \I__1715\ : InMux
    port map (
            O => \N__18728\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\
        );

    \I__1714\ : CascadeMux
    port map (
            O => \N__18725\,
            I => \N__18722\
        );

    \I__1713\ : InMux
    port map (
            O => \N__18722\,
            I => \N__18719\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__18719\,
            I => \N__18716\
        );

    \I__1711\ : Span4Mux_h
    port map (
            O => \N__18716\,
            I => \N__18713\
        );

    \I__1710\ : Odrv4
    port map (
            O => \N__18713\,
            I => \pwm_generator_inst.un2_threshold_acc_2_14\
        );

    \I__1709\ : InMux
    port map (
            O => \N__18710\,
            I => \N__18707\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__18707\,
            I => \N__18704\
        );

    \I__1707\ : Odrv4
    port map (
            O => \N__18704\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0\
        );

    \I__1706\ : InMux
    port map (
            O => \N__18701\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\
        );

    \I__1705\ : InMux
    port map (
            O => \N__18698\,
            I => \N__18695\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__18695\,
            I => \N__18692\
        );

    \I__1703\ : Odrv4
    port map (
            O => \N__18692\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0\
        );

    \I__1702\ : CascadeMux
    port map (
            O => \N__18689\,
            I => \N__18682\
        );

    \I__1701\ : CascadeMux
    port map (
            O => \N__18688\,
            I => \N__18678\
        );

    \I__1700\ : CascadeMux
    port map (
            O => \N__18687\,
            I => \N__18674\
        );

    \I__1699\ : InMux
    port map (
            O => \N__18686\,
            I => \N__18668\
        );

    \I__1698\ : InMux
    port map (
            O => \N__18685\,
            I => \N__18668\
        );

    \I__1697\ : InMux
    port map (
            O => \N__18682\,
            I => \N__18655\
        );

    \I__1696\ : InMux
    port map (
            O => \N__18681\,
            I => \N__18655\
        );

    \I__1695\ : InMux
    port map (
            O => \N__18678\,
            I => \N__18655\
        );

    \I__1694\ : InMux
    port map (
            O => \N__18677\,
            I => \N__18655\
        );

    \I__1693\ : InMux
    port map (
            O => \N__18674\,
            I => \N__18655\
        );

    \I__1692\ : InMux
    port map (
            O => \N__18673\,
            I => \N__18655\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__18668\,
            I => \N__18650\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__18655\,
            I => \N__18650\
        );

    \I__1689\ : Span4Mux_v
    port map (
            O => \N__18650\,
            I => \N__18647\
        );

    \I__1688\ : Odrv4
    port map (
            O => \N__18647\,
            I => \pwm_generator_inst.un2_threshold_acc_1_25\
        );

    \I__1687\ : InMux
    port map (
            O => \N__18644\,
            I => \N__18641\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__18641\,
            I => \N__18638\
        );

    \I__1685\ : Odrv4
    port map (
            O => \N__18638\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0\
        );

    \I__1684\ : InMux
    port map (
            O => \N__18635\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\
        );

    \I__1683\ : InMux
    port map (
            O => \N__18632\,
            I => \N__18629\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__18629\,
            I => \N__18626\
        );

    \I__1681\ : Odrv4
    port map (
            O => \N__18626\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16\
        );

    \I__1680\ : InMux
    port map (
            O => \N__18623\,
            I => \N__18620\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__18620\,
            I => \N__18617\
        );

    \I__1678\ : Odrv4
    port map (
            O => \N__18617\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO\
        );

    \I__1677\ : InMux
    port map (
            O => \N__18614\,
            I => \bfn_1_14_0_\
        );

    \I__1676\ : InMux
    port map (
            O => \N__18611\,
            I => \N__18608\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__18608\,
            I => \N_110_i_i\
        );

    \I__1674\ : InMux
    port map (
            O => \N__18605\,
            I => \N__18602\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__18602\,
            I => \N__18599\
        );

    \I__1672\ : Span4Mux_v
    port map (
            O => \N__18599\,
            I => \N__18596\
        );

    \I__1671\ : Odrv4
    port map (
            O => \N__18596\,
            I => \pwm_generator_inst.un2_threshold_acc_1_18\
        );

    \I__1670\ : CascadeMux
    port map (
            O => \N__18593\,
            I => \N__18590\
        );

    \I__1669\ : InMux
    port map (
            O => \N__18590\,
            I => \N__18587\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__18587\,
            I => \N__18584\
        );

    \I__1667\ : Span4Mux_v
    port map (
            O => \N__18584\,
            I => \N__18581\
        );

    \I__1666\ : Odrv4
    port map (
            O => \N__18581\,
            I => \pwm_generator_inst.un2_threshold_acc_2_3\
        );

    \I__1665\ : CascadeMux
    port map (
            O => \N__18578\,
            I => \N__18575\
        );

    \I__1664\ : InMux
    port map (
            O => \N__18575\,
            I => \N__18572\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__18572\,
            I => \N__18569\
        );

    \I__1662\ : Odrv4
    port map (
            O => \N__18569\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0\
        );

    \I__1661\ : InMux
    port map (
            O => \N__18566\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\
        );

    \I__1660\ : InMux
    port map (
            O => \N__18563\,
            I => \N__18560\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__18560\,
            I => \N__18557\
        );

    \I__1658\ : Span4Mux_v
    port map (
            O => \N__18557\,
            I => \N__18554\
        );

    \I__1657\ : Odrv4
    port map (
            O => \N__18554\,
            I => \pwm_generator_inst.un2_threshold_acc_1_19\
        );

    \I__1656\ : CascadeMux
    port map (
            O => \N__18551\,
            I => \N__18548\
        );

    \I__1655\ : InMux
    port map (
            O => \N__18548\,
            I => \N__18545\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__18545\,
            I => \N__18542\
        );

    \I__1653\ : Odrv4
    port map (
            O => \N__18542\,
            I => \pwm_generator_inst.un2_threshold_acc_2_4\
        );

    \I__1652\ : InMux
    port map (
            O => \N__18539\,
            I => \N__18536\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__18536\,
            I => \N__18533\
        );

    \I__1650\ : Odrv4
    port map (
            O => \N__18533\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0\
        );

    \I__1649\ : InMux
    port map (
            O => \N__18530\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\
        );

    \I__1648\ : InMux
    port map (
            O => \N__18527\,
            I => \N__18524\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__18524\,
            I => \N__18521\
        );

    \I__1646\ : Span4Mux_v
    port map (
            O => \N__18521\,
            I => \N__18518\
        );

    \I__1645\ : Odrv4
    port map (
            O => \N__18518\,
            I => \pwm_generator_inst.un2_threshold_acc_1_20\
        );

    \I__1644\ : CascadeMux
    port map (
            O => \N__18515\,
            I => \N__18512\
        );

    \I__1643\ : InMux
    port map (
            O => \N__18512\,
            I => \N__18509\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__18509\,
            I => \N__18506\
        );

    \I__1641\ : Span4Mux_h
    port map (
            O => \N__18506\,
            I => \N__18503\
        );

    \I__1640\ : Odrv4
    port map (
            O => \N__18503\,
            I => \pwm_generator_inst.un2_threshold_acc_2_5\
        );

    \I__1639\ : InMux
    port map (
            O => \N__18500\,
            I => \N__18497\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__18497\,
            I => \N__18494\
        );

    \I__1637\ : Odrv4
    port map (
            O => \N__18494\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0\
        );

    \I__1636\ : InMux
    port map (
            O => \N__18491\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\
        );

    \I__1635\ : InMux
    port map (
            O => \N__18488\,
            I => \N__18485\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__18485\,
            I => \N__18482\
        );

    \I__1633\ : Span4Mux_v
    port map (
            O => \N__18482\,
            I => \N__18479\
        );

    \I__1632\ : Odrv4
    port map (
            O => \N__18479\,
            I => \pwm_generator_inst.un2_threshold_acc_1_21\
        );

    \I__1631\ : CascadeMux
    port map (
            O => \N__18476\,
            I => \N__18473\
        );

    \I__1630\ : InMux
    port map (
            O => \N__18473\,
            I => \N__18470\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__18470\,
            I => \N__18467\
        );

    \I__1628\ : Span4Mux_h
    port map (
            O => \N__18467\,
            I => \N__18464\
        );

    \I__1627\ : Odrv4
    port map (
            O => \N__18464\,
            I => \pwm_generator_inst.un2_threshold_acc_2_6\
        );

    \I__1626\ : InMux
    port map (
            O => \N__18461\,
            I => \N__18458\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__18458\,
            I => \N__18455\
        );

    \I__1624\ : Odrv4
    port map (
            O => \N__18455\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0\
        );

    \I__1623\ : InMux
    port map (
            O => \N__18452\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\
        );

    \I__1622\ : InMux
    port map (
            O => \N__18449\,
            I => \N__18446\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__18446\,
            I => \N__18443\
        );

    \I__1620\ : Span4Mux_v
    port map (
            O => \N__18443\,
            I => \N__18440\
        );

    \I__1619\ : Odrv4
    port map (
            O => \N__18440\,
            I => \pwm_generator_inst.un2_threshold_acc_1_22\
        );

    \I__1618\ : CascadeMux
    port map (
            O => \N__18437\,
            I => \N__18434\
        );

    \I__1617\ : InMux
    port map (
            O => \N__18434\,
            I => \N__18431\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__18431\,
            I => \N__18428\
        );

    \I__1615\ : Odrv4
    port map (
            O => \N__18428\,
            I => \pwm_generator_inst.un2_threshold_acc_2_7\
        );

    \I__1614\ : InMux
    port map (
            O => \N__18425\,
            I => \N__18422\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__18422\,
            I => \N__18419\
        );

    \I__1612\ : Odrv4
    port map (
            O => \N__18419\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0\
        );

    \I__1611\ : InMux
    port map (
            O => \N__18416\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\
        );

    \I__1610\ : InMux
    port map (
            O => \N__18413\,
            I => \N__18410\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__18410\,
            I => \N__18407\
        );

    \I__1608\ : Span4Mux_v
    port map (
            O => \N__18407\,
            I => \N__18404\
        );

    \I__1607\ : Odrv4
    port map (
            O => \N__18404\,
            I => \pwm_generator_inst.un2_threshold_acc_1_23\
        );

    \I__1606\ : CascadeMux
    port map (
            O => \N__18401\,
            I => \N__18398\
        );

    \I__1605\ : InMux
    port map (
            O => \N__18398\,
            I => \N__18395\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__18395\,
            I => \N__18392\
        );

    \I__1603\ : Odrv4
    port map (
            O => \N__18392\,
            I => \pwm_generator_inst.un2_threshold_acc_2_8\
        );

    \I__1602\ : CascadeMux
    port map (
            O => \N__18389\,
            I => \N__18386\
        );

    \I__1601\ : InMux
    port map (
            O => \N__18386\,
            I => \N__18383\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__18383\,
            I => \N__18380\
        );

    \I__1599\ : Odrv4
    port map (
            O => \N__18380\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0\
        );

    \I__1598\ : InMux
    port map (
            O => \N__18377\,
            I => \bfn_1_13_0_\
        );

    \I__1597\ : InMux
    port map (
            O => \N__18374\,
            I => \N__18371\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__18371\,
            I => \N__18368\
        );

    \I__1595\ : Span4Mux_v
    port map (
            O => \N__18368\,
            I => \N__18365\
        );

    \I__1594\ : Span4Mux_s1_h
    port map (
            O => \N__18365\,
            I => \N__18362\
        );

    \I__1593\ : Odrv4
    port map (
            O => \N__18362\,
            I => \pwm_generator_inst.un2_threshold_acc_1_24\
        );

    \I__1592\ : CascadeMux
    port map (
            O => \N__18359\,
            I => \N__18356\
        );

    \I__1591\ : InMux
    port map (
            O => \N__18356\,
            I => \N__18353\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__18353\,
            I => \N__18350\
        );

    \I__1589\ : Span4Mux_h
    port map (
            O => \N__18350\,
            I => \N__18347\
        );

    \I__1588\ : Odrv4
    port map (
            O => \N__18347\,
            I => \pwm_generator_inst.un2_threshold_acc_2_9\
        );

    \I__1587\ : InMux
    port map (
            O => \N__18344\,
            I => \N__18341\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__18341\,
            I => \N__18338\
        );

    \I__1585\ : Odrv4
    port map (
            O => \N__18338\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0\
        );

    \I__1584\ : InMux
    port map (
            O => \N__18335\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\
        );

    \I__1583\ : InMux
    port map (
            O => \N__18332\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_19\
        );

    \I__1582\ : InMux
    port map (
            O => \N__18329\,
            I => \N__18326\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__18326\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1_16\
        );

    \I__1580\ : CascadeMux
    port map (
            O => \N__18323\,
            I => \N__18320\
        );

    \I__1579\ : InMux
    port map (
            O => \N__18320\,
            I => \N__18314\
        );

    \I__1578\ : InMux
    port map (
            O => \N__18319\,
            I => \N__18314\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__18314\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1_15\
        );

    \I__1576\ : InMux
    port map (
            O => \N__18311\,
            I => \N__18308\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__18308\,
            I => \N__18305\
        );

    \I__1574\ : Odrv4
    port map (
            O => \N__18305\,
            I => \pwm_generator_inst.un2_threshold_acc_2_0\
        );

    \I__1573\ : CascadeMux
    port map (
            O => \N__18302\,
            I => \N__18299\
        );

    \I__1572\ : InMux
    port map (
            O => \N__18299\,
            I => \N__18296\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__18296\,
            I => \N__18293\
        );

    \I__1570\ : Span4Mux_v
    port map (
            O => \N__18293\,
            I => \N__18290\
        );

    \I__1569\ : Odrv4
    port map (
            O => \N__18290\,
            I => \pwm_generator_inst.un2_threshold_acc_1_15\
        );

    \I__1568\ : InMux
    port map (
            O => \N__18287\,
            I => \N__18284\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__18284\,
            I => \N__18281\
        );

    \I__1566\ : Odrv4
    port map (
            O => \N__18281\,
            I => \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4\
        );

    \I__1565\ : InMux
    port map (
            O => \N__18278\,
            I => \N__18275\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__18275\,
            I => \N__18272\
        );

    \I__1563\ : Span4Mux_v
    port map (
            O => \N__18272\,
            I => \N__18269\
        );

    \I__1562\ : Odrv4
    port map (
            O => \N__18269\,
            I => \pwm_generator_inst.un2_threshold_acc_1_16\
        );

    \I__1561\ : CascadeMux
    port map (
            O => \N__18266\,
            I => \N__18263\
        );

    \I__1560\ : InMux
    port map (
            O => \N__18263\,
            I => \N__18260\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__18260\,
            I => \N__18257\
        );

    \I__1558\ : Odrv4
    port map (
            O => \N__18257\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1\
        );

    \I__1557\ : CascadeMux
    port map (
            O => \N__18254\,
            I => \N__18251\
        );

    \I__1556\ : InMux
    port map (
            O => \N__18251\,
            I => \N__18248\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__18248\,
            I => \N__18245\
        );

    \I__1554\ : Odrv4
    port map (
            O => \N__18245\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0\
        );

    \I__1553\ : InMux
    port map (
            O => \N__18242\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\
        );

    \I__1552\ : InMux
    port map (
            O => \N__18239\,
            I => \N__18236\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__18236\,
            I => \N__18233\
        );

    \I__1550\ : Span4Mux_v
    port map (
            O => \N__18233\,
            I => \N__18230\
        );

    \I__1549\ : Odrv4
    port map (
            O => \N__18230\,
            I => \pwm_generator_inst.un2_threshold_acc_1_17\
        );

    \I__1548\ : CascadeMux
    port map (
            O => \N__18227\,
            I => \N__18224\
        );

    \I__1547\ : InMux
    port map (
            O => \N__18224\,
            I => \N__18221\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__18221\,
            I => \N__18218\
        );

    \I__1545\ : Span4Mux_v
    port map (
            O => \N__18218\,
            I => \N__18215\
        );

    \I__1544\ : Odrv4
    port map (
            O => \N__18215\,
            I => \pwm_generator_inst.un2_threshold_acc_2_2\
        );

    \I__1543\ : InMux
    port map (
            O => \N__18212\,
            I => \N__18209\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__18209\,
            I => \N__18206\
        );

    \I__1541\ : Odrv4
    port map (
            O => \N__18206\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0\
        );

    \I__1540\ : InMux
    port map (
            O => \N__18203\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\
        );

    \I__1539\ : InMux
    port map (
            O => \N__18200\,
            I => \bfn_1_10_0_\
        );

    \I__1538\ : InMux
    port map (
            O => \N__18197\,
            I => \N__18194\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__18194\,
            I => \N__18191\
        );

    \I__1536\ : Odrv4
    port map (
            O => \N__18191\,
            I => \pwm_generator_inst.O_12\
        );

    \I__1535\ : InMux
    port map (
            O => \N__18188\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_0\
        );

    \I__1534\ : InMux
    port map (
            O => \N__18185\,
            I => \N__18182\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__18182\,
            I => \N__18179\
        );

    \I__1532\ : Odrv4
    port map (
            O => \N__18179\,
            I => \pwm_generator_inst.O_13\
        );

    \I__1531\ : InMux
    port map (
            O => \N__18176\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_1\
        );

    \I__1530\ : InMux
    port map (
            O => \N__18173\,
            I => \N__18170\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__18170\,
            I => \N__18167\
        );

    \I__1528\ : Span4Mux_h
    port map (
            O => \N__18167\,
            I => \N__18164\
        );

    \I__1527\ : Odrv4
    port map (
            O => \N__18164\,
            I => \pwm_generator_inst.O_14\
        );

    \I__1526\ : InMux
    port map (
            O => \N__18161\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_2\
        );

    \I__1525\ : InMux
    port map (
            O => \N__18158\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_3\
        );

    \I__1524\ : InMux
    port map (
            O => \N__18155\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_4\
        );

    \I__1523\ : InMux
    port map (
            O => \N__18152\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_5\
        );

    \I__1522\ : InMux
    port map (
            O => \N__18149\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_6\
        );

    \I__1521\ : InMux
    port map (
            O => \N__18146\,
            I => \N__18137\
        );

    \I__1520\ : InMux
    port map (
            O => \N__18145\,
            I => \N__18137\
        );

    \I__1519\ : InMux
    port map (
            O => \N__18144\,
            I => \N__18137\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__18137\,
            I => \N__18134\
        );

    \I__1517\ : Odrv4
    port map (
            O => \N__18134\,
            I => \current_shift_inst.PI_CTRL.N_97\
        );

    \IN_MUX_bfv_8_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_17_0_\
        );

    \IN_MUX_bfv_8_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_0_cry_6\,
            carryinitout => \bfn_8_18_0_\
        );

    \IN_MUX_bfv_8_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_0_cry_14\,
            carryinitout => \bfn_8_19_0_\
        );

    \IN_MUX_bfv_8_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_0_cry_22\,
            carryinitout => \bfn_8_20_0_\
        );

    \IN_MUX_bfv_8_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_0_cry_30\,
            carryinitout => \bfn_8_21_0_\
        );

    \IN_MUX_bfv_4_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_7_0_\
        );

    \IN_MUX_bfv_4_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un5_counter_cry_8,
            carryinitout => \bfn_4_8_0_\
        );

    \IN_MUX_bfv_1_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_9_0_\
        );

    \IN_MUX_bfv_1_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_acc_cry_7\,
            carryinitout => \bfn_1_10_0_\
        );

    \IN_MUX_bfv_1_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_acc_cry_15\,
            carryinitout => \bfn_1_11_0_\
        );

    \IN_MUX_bfv_14_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_22_0_\
        );

    \IN_MUX_bfv_14_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_14_23_0_\
        );

    \IN_MUX_bfv_14_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_14_24_0_\
        );

    \IN_MUX_bfv_15_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_17_0_\
        );

    \IN_MUX_bfv_15_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_15_18_0_\
        );

    \IN_MUX_bfv_15_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_15_19_0_\
        );

    \IN_MUX_bfv_13_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_23_0_\
        );

    \IN_MUX_bfv_13_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_13_24_0_\
        );

    \IN_MUX_bfv_13_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_13_25_0_\
        );

    \IN_MUX_bfv_18_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_17_0_\
        );

    \IN_MUX_bfv_18_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_18_18_0_\
        );

    \IN_MUX_bfv_18_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_18_19_0_\
        );

    \IN_MUX_bfv_8_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_11_0_\
        );

    \IN_MUX_bfv_8_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_8_12_0_\
        );

    \IN_MUX_bfv_8_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_8_13_0_\
        );

    \IN_MUX_bfv_11_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_8_0_\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_11_9_0_\
        );

    \IN_MUX_bfv_11_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_11_10_0_\
        );

    \IN_MUX_bfv_10_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_18_0_\
        );

    \IN_MUX_bfv_10_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.z_5_cry_8\,
            carryinitout => \bfn_10_19_0_\
        );

    \IN_MUX_bfv_10_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.z_5_cry_16\,
            carryinitout => \bfn_10_20_0_\
        );

    \IN_MUX_bfv_10_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.z_5_cry_24\,
            carryinitout => \bfn_10_21_0_\
        );

    \IN_MUX_bfv_1_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_12_0_\
        );

    \IN_MUX_bfv_1_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7\,
            carryinitout => \bfn_1_13_0_\
        );

    \IN_MUX_bfv_1_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15\,
            carryinitout => \bfn_1_14_0_\
        );

    \IN_MUX_bfv_2_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_7_0_\
        );

    \IN_MUX_bfv_2_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_acc_1_cry_7\,
            carryinitout => \bfn_2_8_0_\
        );

    \IN_MUX_bfv_2_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_acc_1_cry_15\,
            carryinitout => \bfn_2_9_0_\
        );

    \IN_MUX_bfv_9_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_8_0_\
        );

    \IN_MUX_bfv_9_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un14_counter_cry_7\,
            carryinitout => \bfn_9_9_0_\
        );

    \IN_MUX_bfv_3_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_9_0_\
        );

    \IN_MUX_bfv_3_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un19_threshold_acc_cry_7\,
            carryinitout => \bfn_3_10_0_\
        );

    \IN_MUX_bfv_10_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_9_0_\
        );

    \IN_MUX_bfv_10_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.counter_cry_7\,
            carryinitout => \bfn_10_10_0_\
        );

    \IN_MUX_bfv_13_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_19_0_\
        );

    \IN_MUX_bfv_13_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8\,
            carryinitout => \bfn_13_20_0_\
        );

    \IN_MUX_bfv_13_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16\,
            carryinitout => \bfn_13_21_0_\
        );

    \IN_MUX_bfv_16_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_19_0_\
        );

    \IN_MUX_bfv_16_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            carryinitout => \bfn_16_20_0_\
        );

    \IN_MUX_bfv_16_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            carryinitout => \bfn_16_21_0_\
        );

    \IN_MUX_bfv_18_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_13_0_\
        );

    \IN_MUX_bfv_18_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_18_14_0_\
        );

    \IN_MUX_bfv_18_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_18_15_0_\
        );

    \IN_MUX_bfv_18_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_18_16_0_\
        );

    \IN_MUX_bfv_17_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_11_0_\
        );

    \IN_MUX_bfv_17_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            carryinitout => \bfn_17_12_0_\
        );

    \IN_MUX_bfv_17_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            carryinitout => \bfn_17_13_0_\
        );

    \IN_MUX_bfv_17_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            carryinitout => \bfn_17_14_0_\
        );

    \IN_MUX_bfv_15_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_7_0_\
        );

    \IN_MUX_bfv_15_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_15_8_0_\
        );

    \IN_MUX_bfv_15_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_15_9_0_\
        );

    \IN_MUX_bfv_15_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_15_10_0_\
        );

    \IN_MUX_bfv_16_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_7_0_\
        );

    \IN_MUX_bfv_16_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            carryinitout => \bfn_16_8_0_\
        );

    \IN_MUX_bfv_16_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            carryinitout => \bfn_16_9_0_\
        );

    \IN_MUX_bfv_16_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            carryinitout => \bfn_16_10_0_\
        );

    \IN_MUX_bfv_10_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_14_0_\
        );

    \IN_MUX_bfv_10_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.z_cry_7\,
            carryinitout => \bfn_10_15_0_\
        );

    \IN_MUX_bfv_10_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.z_cry_15\,
            carryinitout => \bfn_10_16_0_\
        );

    \IN_MUX_bfv_10_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.z_cry_23\,
            carryinitout => \bfn_10_17_0_\
        );

    \IN_MUX_bfv_11_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_14_0_\
        );

    \IN_MUX_bfv_11_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_cry_8\,
            carryinitout => \bfn_11_15_0_\
        );

    \IN_MUX_bfv_11_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_cry_16\,
            carryinitout => \bfn_11_16_0_\
        );

    \IN_MUX_bfv_11_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_cry_24\,
            carryinitout => \bfn_11_17_0_\
        );

    \IN_MUX_bfv_13_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_13_0_\
        );

    \IN_MUX_bfv_13_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_13_14_0_\
        );

    \IN_MUX_bfv_13_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_13_15_0_\
        );

    \IN_MUX_bfv_13_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_13_16_0_\
        );

    \IN_MUX_bfv_15_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_13_0_\
        );

    \IN_MUX_bfv_15_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_7\,
            carryinitout => \bfn_15_14_0_\
        );

    \IN_MUX_bfv_15_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_15\,
            carryinitout => \bfn_15_15_0_\
        );

    \IN_MUX_bfv_15_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_23\,
            carryinitout => \bfn_15_16_0_\
        );

    \IN_MUX_bfv_9_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_21_0_\
        );

    \IN_MUX_bfv_9_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_9_22_0_\
        );

    \IN_MUX_bfv_9_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_9_23_0_\
        );

    \IN_MUX_bfv_9_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_9_24_0_\
        );

    \IN_MUX_bfv_9_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_25_0_\
        );

    \IN_MUX_bfv_9_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_phase.counter_cry_7\,
            carryinitout => \bfn_9_26_0_\
        );

    \IN_MUX_bfv_9_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_phase.counter_cry_15\,
            carryinitout => \bfn_9_27_0_\
        );

    \IN_MUX_bfv_9_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_phase.counter_cry_23\,
            carryinitout => \bfn_9_28_0_\
        );

    \IN_MUX_bfv_7_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_17_0_\
        );

    \IN_MUX_bfv_7_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_1_cry_7\,
            carryinitout => \bfn_7_18_0_\
        );

    \IN_MUX_bfv_7_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_1_cry_15\,
            carryinitout => \bfn_7_19_0_\
        );

    \IN_MUX_bfv_7_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_1_cry_23\,
            carryinitout => \bfn_7_20_0_\
        );

    \IN_MUX_bfv_4_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_13_0_\
        );

    \IN_MUX_bfv_4_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            carryinitout => \bfn_4_14_0_\
        );

    \IN_MUX_bfv_4_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            carryinitout => \bfn_4_15_0_\
        );

    \IN_MUX_bfv_4_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            carryinitout => \bfn_4_16_0_\
        );

    \IN_MUX_bfv_9_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_13_0_\
        );

    \IN_MUX_bfv_9_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\,
            carryinitout => \bfn_9_14_0_\
        );

    \IN_MUX_bfv_9_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\,
            carryinitout => \bfn_9_15_0_\
        );

    \IN_MUX_bfv_9_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\,
            carryinitout => \bfn_9_16_0_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__32273\,
            GLOBALBUFFEROUTPUT => \delay_measurement_inst.delay_hc_timer.N_321_i_g\
        );

    \current_shift_inst.timer_s1.running_RNII51H_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__32414\,
            GLOBALBUFFEROUTPUT => \current_shift_inst.timer_s1.N_187_i_g\
        );

    \current_shift_inst.timer_phase.running_RNIC90O_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__33452\,
            GLOBALBUFFEROUTPUT => \current_shift_inst.timer_phase.N_188_i_g\
        );

    \osc\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b10"
        )
    port map (
            CLKHFPU => \N__28547\,
            CLKHFEN => \N__28548\,
            CLKHF => clk_12mhz
        );

    \rgb_drv\ : SB_RGBA_DRV
    generic map (
            RGB2_CURRENT => "0b111111",
            CURRENT_MODE => "0b0",
            RGB0_CURRENT => "0b111111",
            RGB1_CURRENT => "0b111111"
        )
    port map (
            RGBLEDEN => \N__28528\,
            RGB2PWM => \N__18611\,
            RGB1 => rgb_g_wire,
            CURREN => \N__28656\,
            RGB2 => rgb_b_wire,
            RGB1PWM => \N__19145\,
            RGB0PWM => \N__46780\,
            RGB0 => rgb_r_wire
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_5_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000001110"
        )
    port map (
            in0 => \N__20501\,
            in1 => \N__19703\,
            in2 => \N__21265\,
            in3 => \N__20001\,
            lcout => pwm_duty_input_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47351\,
            ce => \N__23648\,
            sr => \N__46683\
        );

    \current_shift_inst.PI_CTRL.control_out_7_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101100110000"
        )
    port map (
            in0 => \N__20003\,
            in1 => \N__21253\,
            in2 => \N__19714\,
            in3 => \N__21062\,
            lcout => pwm_duty_input_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47351\,
            ce => \N__23648\,
            sr => \N__46683\
        );

    \current_shift_inst.PI_CTRL.control_out_8_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000001110"
        )
    port map (
            in0 => \N__21029\,
            in1 => \N__19708\,
            in2 => \N__21267\,
            in3 => \N__20004\,
            lcout => pwm_duty_input_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47351\,
            ce => \N__23648\,
            sr => \N__46683\
        );

    \current_shift_inst.PI_CTRL.control_out_9_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101100110000"
        )
    port map (
            in0 => \N__20005\,
            in1 => \N__21257\,
            in2 => \N__19715\,
            in3 => \N__20987\,
            lcout => pwm_duty_input_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47351\,
            ce => \N__23648\,
            sr => \N__46683\
        );

    \current_shift_inst.PI_CTRL.control_out_6_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000001110"
        )
    port map (
            in0 => \N__20471\,
            in1 => \N__19704\,
            in2 => \N__21266\,
            in3 => \N__20002\,
            lcout => pwm_duty_input_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47351\,
            ce => \N__23648\,
            sr => \N__46683\
        );

    \current_shift_inst.PI_CTRL.control_out_0_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__18144\,
            in1 => \N__19026\,
            in2 => \N__20651\,
            in3 => \N__19736\,
            lcout => pwm_duty_input_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47350\,
            ce => \N__23672\,
            sr => \N__46693\
        );

    \current_shift_inst.PI_CTRL.control_out_3_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010111110001"
        )
    port map (
            in0 => \N__19739\,
            in1 => \N__19043\,
            in2 => \N__20594\,
            in3 => \N__19712\,
            lcout => pwm_duty_input_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47350\,
            ce => \N__23672\,
            sr => \N__46693\
        );

    \current_shift_inst.PI_CTRL.control_out_4_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000101010101"
        )
    port map (
            in0 => \N__19649\,
            in1 => \N__19886\,
            in2 => \N__20552\,
            in3 => \N__20006\,
            lcout => pwm_duty_input_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47350\,
            ce => \N__23672\,
            sr => \N__46693\
        );

    \current_shift_inst.PI_CTRL.control_out_1_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__19737\,
            in1 => \N__20633\,
            in2 => \N__19031\,
            in3 => \N__18145\,
            lcout => pwm_duty_input_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47350\,
            ce => \N__23672\,
            sr => \N__46693\
        );

    \current_shift_inst.PI_CTRL.control_out_2_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__18146\,
            in1 => \N__19030\,
            in2 => \N__20615\,
            in3 => \N__19738\,
            lcout => pwm_duty_input_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47350\,
            ce => \N__23672\,
            sr => \N__46693\
        );

    \current_shift_inst.PI_CTRL.control_out_10_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21246\,
            lcout => pwm_duty_input_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47349\,
            ce => \N__23578\,
            sr => \N__46703\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__19489\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19510\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__19685\,
            in1 => \N__21245\,
            in2 => \_gnd_net_\,
            in3 => \N__20057\,
            lcout => \current_shift_inst.PI_CTRL.N_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20197\,
            in2 => \_gnd_net_\,
            in3 => \N__20182\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19324\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_9_0_\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18197\,
            in2 => \_gnd_net_\,
            in3 => \N__18188\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_0\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18185\,
            in2 => \_gnd_net_\,
            in3 => \N__18176\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_1\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18173\,
            in2 => \_gnd_net_\,
            in3 => \N__18161\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_2\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18287\,
            in2 => \_gnd_net_\,
            in3 => \N__18158\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_3\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28796\,
            in2 => \N__18254\,
            in3 => \N__18155\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_4\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18212\,
            in2 => \N__28848\,
            in3 => \N__18152\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_5\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28800\,
            in2 => \N__18578\,
            in3 => \N__18149\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_6\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18539\,
            in2 => \_gnd_net_\,
            in3 => \N__18200\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_1_10_0_\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18500\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_8\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18461\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_9\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18425\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_10\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18389\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_11\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18344\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_12\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18815\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_13\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18791\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_14\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18761\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_11_0_\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18737\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_16\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18710\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_17\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18644\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_18\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18332\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__18686\,
            in1 => \N__18319\,
            in2 => \_gnd_net_\,
            in3 => \N__18952\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__18953\,
            in1 => \N__18329\,
            in2 => \N__18323\,
            in3 => \N__18685\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_axb_4_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18311\,
            in2 => \N__18302\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \bfn_1_12_0_\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18278\,
            in2 => \N__18266\,
            in3 => \N__18242\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18239\,
            in2 => \N__18227\,
            in3 => \N__18203\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18605\,
            in2 => \N__18593\,
            in3 => \N__18566\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18563\,
            in2 => \N__18551\,
            in3 => \N__18530\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18527\,
            in2 => \N__18515\,
            in3 => \N__18491\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18488\,
            in2 => \N__18476\,
            in3 => \N__18452\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18449\,
            in2 => \N__18437\,
            in3 => \N__18416\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18413\,
            in2 => \N__18401\,
            in3 => \N__18377\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0\,
            ltout => OPEN,
            carryin => \bfn_1_13_0_\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18374\,
            in2 => \N__18359\,
            in3 => \N__18335\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18673\,
            in2 => \N__18830\,
            in3 => \N__18806\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18803\,
            in2 => \N__18687\,
            in3 => \N__18779\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18677\,
            in2 => \N__18776\,
            in3 => \N__18752\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18749\,
            in2 => \N__18688\,
            in3 => \N__18728\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18681\,
            in2 => \N__18725\,
            in3 => \N__18701\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18698\,
            in2 => \N__18689\,
            in3 => \N__18635\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__18632\,
            in1 => \N__18623\,
            in2 => \_gnd_net_\,
            in3 => \N__18614\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.N_110_i_i_LC_1_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__46778\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34564\,
            lcout => \N_110_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un7_start_stop_LC_1_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__46779\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34568\,
            lcout => un7_start_stop,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNILM9T_5_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19116\,
            in1 => \N__19137\,
            in2 => \N__19099\,
            in3 => \N__19062\,
            lcout => \current_shift_inst.PI_CTRL.m14_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNIDE9T_3_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__19003\,
            in1 => \N__19138\,
            in2 => \N__19121\,
            in3 => \N__18847\,
            lcout => \current_shift_inst.PI_CTRL.m7_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNIVCED1_7_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__19095\,
            in1 => \N__18886\,
            in2 => \N__19073\,
            in3 => \N__19063\,
            lcout => i8_mux,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010001"
        )
    port map (
            in0 => \N__21269\,
            in1 => \N__20548\,
            in2 => \_gnd_net_\,
            in3 => \N__20055\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010000"
        )
    port map (
            in0 => \N__20590\,
            in1 => \N__19681\,
            in2 => \N__19034\,
            in3 => \N__19726\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNIUU8T_0_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__19016\,
            in1 => \N__19004\,
            in2 => \N__18986\,
            in3 => \N__18971\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.N_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNIK2D32_4_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100000"
        )
    port map (
            in0 => \N__18959\,
            in1 => \N__18885\,
            in2 => \N__18851\,
            in3 => \N__18848\,
            lcout => \N_28_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19277\,
            in2 => \_gnd_net_\,
            in3 => \N__19289\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_2_7_0_\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19259\,
            in2 => \_gnd_net_\,
            in3 => \N__19271\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_0\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19241\,
            in2 => \_gnd_net_\,
            in3 => \N__19253\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_1\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19223\,
            in2 => \_gnd_net_\,
            in3 => \N__19235\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_2\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19205\,
            in2 => \_gnd_net_\,
            in3 => \N__19217\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_3\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19187\,
            in2 => \_gnd_net_\,
            in3 => \N__19199\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_4\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19169\,
            in2 => \_gnd_net_\,
            in3 => \N__19181\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_5\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19151\,
            in2 => \_gnd_net_\,
            in3 => \N__19163\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_6\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19355\,
            in2 => \_gnd_net_\,
            in3 => \N__19367\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_8\,
            ltout => OPEN,
            carryin => \bfn_2_8_0_\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19337\,
            in2 => \_gnd_net_\,
            in3 => \N__19349\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_8\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19485\,
            in2 => \_gnd_net_\,
            in3 => \N__19331\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_9\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__20132\,
            in1 => \N__19328\,
            in2 => \_gnd_net_\,
            in3 => \N__19307\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_10\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19780\,
            in3 => \N__19304\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_11\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19537\,
            in2 => \_gnd_net_\,
            in3 => \N__19301\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_12\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20178\,
            in2 => \_gnd_net_\,
            in3 => \N__19298\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_13\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19443\,
            in2 => \_gnd_net_\,
            in3 => \N__19295\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_14\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19566\,
            in2 => \_gnd_net_\,
            in3 => \N__19292\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_2_9_0_\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19399\,
            in2 => \_gnd_net_\,
            in3 => \N__19454\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_16\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19628\,
            in3 => \N__19451\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_17\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19448\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19795\,
            in2 => \_gnd_net_\,
            in3 => \N__19779\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19588\,
            in2 => \_gnd_net_\,
            in3 => \N__19567\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__19445\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19426\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010111001100"
        )
    port map (
            in0 => \N__19444\,
            in1 => \N__19427\,
            in2 => \N__19415\,
            in3 => \N__20135\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__19403\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19387\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_17\,
            ltout => \pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001001110"
        )
    port map (
            in0 => \N__20136\,
            in1 => \N__19388\,
            in2 => \N__19376\,
            in3 => \N__19373\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010111001100"
        )
    port map (
            in0 => \N__19538\,
            in1 => \N__19552\,
            in2 => \N__19640\,
            in3 => \N__20133\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__19609\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19627\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_18\,
            ltout => \pwm_generator_inst.un15_threshold_acc_1_axb_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__19613\,
            in1 => \N__20137\,
            in2 => \N__19598\,
            in3 => \N__19595\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001001110"
        )
    port map (
            in0 => \N__20134\,
            in1 => \N__19589\,
            in2 => \N__19577\,
            in3 => \N__19568\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_9_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000001010000"
        )
    port map (
            in0 => \N__20702\,
            in1 => \N__20768\,
            in2 => \N__19895\,
            in3 => \N__20854\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47339\,
            ce => 'H',
            sr => \N__46719\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__19536\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19553\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__19517\,
            in1 => \N__19493\,
            in2 => \N__19469\,
            in3 => \N__20094\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_2_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__44205\,
            in1 => \N__40328\,
            in2 => \N__34114\,
            in3 => \N__43912\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47330\,
            ce => \N__31224\,
            sr => \N__46727\
        );

    \phase_controller_inst1.stoper_hc.target_time_1_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111010101010"
        )
    port map (
            in0 => \N__44204\,
            in1 => \N__40327\,
            in2 => \N__41276\,
            in3 => \N__43911\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47330\,
            ce => \N__31224\,
            sr => \N__46727\
        );

    \phase_controller_inst1.stoper_hc.target_time_3_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111011101100"
        )
    port map (
            in0 => \N__43913\,
            in1 => \N__44206\,
            in2 => \N__40343\,
            in3 => \N__35522\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47330\,
            ce => \N__31224\,
            sr => \N__46727\
        );

    \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001000000011"
        )
    port map (
            in0 => \N__34169\,
            in1 => \N__40326\,
            in2 => \N__44207\,
            in3 => \N__43910\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ1Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47330\,
            ce => \N__31224\,
            sr => \N__46727\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__19802\,
            in1 => \N__19784\,
            in2 => \N__19757\,
            in3 => \N__20101\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_10_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20258\,
            in1 => \N__20228\,
            in2 => \N__20024\,
            in3 => \N__20222\,
            lcout => \current_shift_inst.PI_CTRL.N_178\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_3_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__20583\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20540\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.N_98_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_3_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__19882\,
            in1 => \N__21258\,
            in2 => \N__19742\,
            in3 => \N__20000\,
            lcout => \current_shift_inst.PI_CTRL.N_96\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_3_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000111"
        )
    port map (
            in0 => \N__20541\,
            in1 => \N__20056\,
            in2 => \N__21268\,
            in3 => \N__19713\,
            lcout => \current_shift_inst.PI_CTRL.N_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_LC_3_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21466\,
            in2 => \_gnd_net_\,
            in3 => \N__21427\,
            lcout => \counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47348\,
            ce => 'H',
            sr => \N__46684\
        );

    \counter_RNIM6001_12_LC_3_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__20431\,
            in1 => \N__20272\,
            in2 => \N__20291\,
            in3 => \N__20416\,
            lcout => un2_counter_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNII76D_3_LC_3_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20326\,
            in1 => \N__20341\,
            in2 => \N__20312\,
            in3 => \N__20356\,
            lcout => un2_counter_7,
            ltout => \un2_counter_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_0_LC_3_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__21667\,
            in1 => \N__21426\,
            in2 => \N__19859\,
            in3 => \N__21714\,
            lcout => \counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47348\,
            ce => 'H',
            sr => \N__46684\
        );

    \pwm_generator_inst.threshold_ACC_7_LC_3_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110101100"
        )
    port map (
            in0 => \N__20777\,
            in1 => \N__20721\,
            in2 => \N__20859\,
            in3 => \N__19937\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47346\,
            ce => 'H',
            sr => \N__46694\
        );

    \counter_12_LC_3_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__20402\,
            in1 => \N__21711\,
            in2 => \N__21674\,
            in3 => \N__21619\,
            lcout => \counterZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47346\,
            ce => 'H',
            sr => \N__46694\
        );

    \pwm_generator_inst.threshold_ACC_2_LC_3_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101001100000000"
        )
    port map (
            in0 => \N__20776\,
            in1 => \N__20720\,
            in2 => \N__20858\,
            in3 => \N__19820\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47346\,
            ce => 'H',
            sr => \N__46694\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_3_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19856\,
            in2 => \N__20150\,
            in3 => \N__20149\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_3_9_0_\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_3_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19844\,
            in3 => \N__19835\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_0\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_3_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19832\,
            in2 => \_gnd_net_\,
            in3 => \N__19814\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_1\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_3_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19811\,
            in2 => \_gnd_net_\,
            in3 => \N__19805\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_2\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_3_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20066\,
            in2 => \_gnd_net_\,
            in3 => \N__19964\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_3\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_3_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19961\,
            in2 => \_gnd_net_\,
            in3 => \N__19955\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_4\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_3_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19952\,
            in2 => \_gnd_net_\,
            in3 => \N__19946\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_5\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_3_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19943\,
            in2 => \_gnd_net_\,
            in3 => \N__19931\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_6\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_3_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19928\,
            in3 => \N__19919\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \bfn_3_10_0_\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_3_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011101111000"
        )
    port map (
            in0 => \N__20139\,
            in1 => \N__19916\,
            in2 => \N__19910\,
            in3 => \N__19898\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_3_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20494\,
            in1 => \N__20467\,
            in2 => \N__21025\,
            in3 => \N__19865\,
            lcout => \current_shift_inst.PI_CTRL.N_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIU1LD_7_LC_3_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20980\,
            in2 => \_gnd_net_\,
            in3 => \N__21061\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_3_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__20204\,
            in1 => \N__20186\,
            in2 => \N__20162\,
            in3 => \N__20138\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIQTKD_5_LC_3_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101110111"
        )
    port map (
            in0 => \N__21057\,
            in1 => \N__20493\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_3_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__20976\,
            in1 => \N__21024\,
            in2 => \N__20060\,
            in3 => \N__20463\,
            lcout => \current_shift_inst.PI_CTRL.N_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMJ62_12_LC_3_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21073\,
            in2 => \_gnd_net_\,
            in3 => \N__20920\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_9_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIU8H5_14_LC_3_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21359\,
            in1 => \N__21388\,
            in2 => \N__20027\,
            in3 => \N__20887\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIEAE4_15_LC_3_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20873\,
            in1 => \N__21107\,
            in2 => \N__21094\,
            in3 => \N__21074\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIFBE4_19_LC_3_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21121\,
            in1 => \N__21106\,
            in2 => \N__21095\,
            in3 => \N__21136\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_3_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20237\,
            in1 => \N__20015\,
            in2 => \N__20009\,
            in3 => \N__20243\,
            lcout => \current_shift_inst.PI_CTRL.N_118\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIPM62_13_LC_3_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21370\,
            in2 => \_gnd_net_\,
            in3 => \N__20905\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIRMD4_17_LC_3_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21389\,
            in1 => \N__21154\,
            in2 => \N__21358\,
            in3 => \N__21167\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIQJB4_15_LC_3_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21166\,
            in1 => \N__21178\,
            in2 => \N__21155\,
            in3 => \N__20872\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIKAQ8_27_LC_3_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21320\,
            in1 => \N__21335\,
            in2 => \N__20252\,
            in3 => \N__20249\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNID9E4_10_LC_3_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21304\,
            in1 => \N__20935\,
            in2 => \N__21290\,
            in3 => \N__20947\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIPL52_13_LC_3_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__20906\,
            in1 => \_gnd_net_\,
            in2 => \N__21182\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISHP8_10_LC_3_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20210\,
            in1 => \N__20936\,
            in2 => \N__20231\,
            in3 => \N__20948\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI9LI5_19_LC_3_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21371\,
            in1 => \N__20216\,
            in2 => \N__21140\,
            in3 => \N__21122\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI1082_27_LC_3_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21319\,
            in2 => \_gnd_net_\,
            in3 => \N__21334\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIIEE4_12_LC_3_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20924\,
            in1 => \N__21289\,
            in2 => \N__20894\,
            in3 => \N__21305\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_counter_cry_1_c_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21425\,
            in2 => \N__21467\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_7_0_\,
            carryout => un5_counter_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_2_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21443\,
            in2 => \_gnd_net_\,
            in3 => \N__20360\,
            lcout => \counterZ0Z_2\,
            ltout => OPEN,
            carryin => un5_counter_cry_1,
            carryout => un5_counter_cry_2,
            clk => \N__47347\,
            ce => 'H',
            sr => \N__46678\
        );

    \counter_3_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20357\,
            in2 => \_gnd_net_\,
            in3 => \N__20345\,
            lcout => \counterZ0Z_3\,
            ltout => OPEN,
            carryin => un5_counter_cry_2,
            carryout => un5_counter_cry_3,
            clk => \N__47347\,
            ce => 'H',
            sr => \N__46678\
        );

    \counter_4_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20342\,
            in2 => \_gnd_net_\,
            in3 => \N__20330\,
            lcout => \counterZ0Z_4\,
            ltout => OPEN,
            carryin => un5_counter_cry_3,
            carryout => un5_counter_cry_4,
            clk => \N__47347\,
            ce => 'H',
            sr => \N__46678\
        );

    \counter_5_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20327\,
            in2 => \_gnd_net_\,
            in3 => \N__20315\,
            lcout => \counterZ0Z_5\,
            ltout => OPEN,
            carryin => un5_counter_cry_4,
            carryout => un5_counter_cry_5,
            clk => \N__47347\,
            ce => 'H',
            sr => \N__46678\
        );

    \counter_6_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20311\,
            in2 => \_gnd_net_\,
            in3 => \N__20297\,
            lcout => \counterZ0Z_6\,
            ltout => OPEN,
            carryin => un5_counter_cry_5,
            carryout => un5_counter_cry_6,
            clk => \N__47347\,
            ce => 'H',
            sr => \N__46678\
        );

    \counter_RNO_0_7_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21479\,
            in2 => \_gnd_net_\,
            in3 => \N__20294\,
            lcout => \counter_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => un5_counter_cry_6,
            carryout => un5_counter_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_8_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20290\,
            in2 => \_gnd_net_\,
            in3 => \N__20276\,
            lcout => \counterZ0Z_8\,
            ltout => OPEN,
            carryin => un5_counter_cry_7,
            carryout => un5_counter_cry_8,
            clk => \N__47347\,
            ce => 'H',
            sr => \N__46678\
        );

    \counter_9_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20273\,
            in2 => \_gnd_net_\,
            in3 => \N__20261\,
            lcout => \counterZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_4_8_0_\,
            carryout => un5_counter_cry_9,
            clk => \N__47344\,
            ce => 'H',
            sr => \N__46685\
        );

    \counter_RNO_0_10_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21593\,
            in2 => \_gnd_net_\,
            in3 => \N__20435\,
            lcout => \counter_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => un5_counter_cry_9,
            carryout => un5_counter_cry_10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_11_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20432\,
            in2 => \_gnd_net_\,
            in3 => \N__20420\,
            lcout => \counterZ0Z_11\,
            ltout => OPEN,
            carryin => un5_counter_cry_10,
            carryout => un5_counter_cry_11,
            clk => \N__47344\,
            ce => 'H',
            sr => \N__46685\
        );

    \counter_RNO_0_12_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20417\,
            in2 => \_gnd_net_\,
            in3 => \N__20405\,
            lcout => \counter_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_0_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000001001100"
        )
    port map (
            in0 => \N__20772\,
            in1 => \N__20396\,
            in2 => \N__20861\,
            in3 => \N__20719\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47340\,
            ce => 'H',
            sr => \N__46695\
        );

    \pwm_generator_inst.threshold_ACC_4_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010011100000000"
        )
    port map (
            in0 => \N__20847\,
            in1 => \N__20775\,
            in2 => \N__20726\,
            in3 => \N__20390\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47340\,
            ce => 'H',
            sr => \N__46695\
        );

    \pwm_generator_inst.threshold_ACC_1_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111111011000"
        )
    port map (
            in0 => \N__20846\,
            in1 => \N__20774\,
            in2 => \N__20725\,
            in3 => \N__20384\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47340\,
            ce => 'H',
            sr => \N__46695\
        );

    \pwm_generator_inst.threshold_ACC_3_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101001100000000"
        )
    port map (
            in0 => \N__20773\,
            in1 => \N__20712\,
            in2 => \N__20860\,
            in3 => \N__20378\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47340\,
            ce => 'H',
            sr => \N__46695\
        );

    \pwm_generator_inst.threshold_ACC_6_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111111011000"
        )
    port map (
            in0 => \N__20855\,
            in1 => \N__20770\,
            in2 => \N__20722\,
            in3 => \N__20372\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47336\,
            ce => 'H',
            sr => \N__46704\
        );

    \pwm_generator_inst.threshold_ACC_5_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100011100000000"
        )
    port map (
            in0 => \N__20769\,
            in1 => \N__20857\,
            in2 => \N__20724\,
            in3 => \N__20366\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47336\,
            ce => 'H',
            sr => \N__46704\
        );

    \pwm_generator_inst.threshold_ACC_8_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111111011000"
        )
    port map (
            in0 => \N__20856\,
            in1 => \N__20771\,
            in2 => \N__20723\,
            in3 => \N__20657\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47336\,
            ce => 'H',
            sr => \N__46704\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_0_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23888\,
            in2 => \N__21530\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_4_13_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\,
            clk => \N__47315\,
            ce => \N__23649\,
            sr => \N__46720\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23834\,
            in2 => \N__21575\,
            in3 => \N__20618\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            clk => \N__47315\,
            ce => \N__23649\,
            sr => \N__46720\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_2_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23783\,
            in2 => \N__21785\,
            in3 => \N__20597\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            clk => \N__47315\,
            ce => \N__23649\,
            sr => \N__46720\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_3_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23711\,
            in2 => \N__21758\,
            in3 => \N__20555\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            clk => \N__47315\,
            ce => \N__23649\,
            sr => \N__46720\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_4_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23497\,
            in2 => \N__21521\,
            in3 => \N__20504\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            clk => \N__47315\,
            ce => \N__23649\,
            sr => \N__46720\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_5_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24476\,
            in2 => \N__21539\,
            in3 => \N__20474\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            clk => \N__47315\,
            ce => \N__23649\,
            sr => \N__46720\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_6_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24398\,
            in2 => \N__21767\,
            in3 => \N__20438\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            clk => \N__47315\,
            ce => \N__23649\,
            sr => \N__46720\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_7_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24302\,
            in2 => \N__22067\,
            in3 => \N__21032\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            clk => \N__47315\,
            ce => \N__23649\,
            sr => \N__46720\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_8_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24260\,
            in2 => \N__21776\,
            in3 => \N__20990\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_4_14_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            clk => \N__47303\,
            ce => \N__23637\,
            sr => \N__46724\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_9_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24197\,
            in2 => \N__21551\,
            in3 => \N__20951\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            clk => \N__47303\,
            ce => \N__23637\,
            sr => \N__46724\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_10_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24126\,
            in2 => \N__21734\,
            in3 => \N__20939\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            clk => \N__47303\,
            ce => \N__23637\,
            sr => \N__46724\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_11_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21560\,
            in2 => \N__24064\,
            in3 => \N__20927\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            clk => \N__47303\,
            ce => \N__23637\,
            sr => \N__46724\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_12_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23989\,
            in2 => \N__21497\,
            in3 => \N__20909\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            clk => \N__47303\,
            ce => \N__23637\,
            sr => \N__46724\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_13_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21725\,
            in2 => \N__24983\,
            in3 => \N__20897\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            clk => \N__47303\,
            ce => \N__23637\,
            sr => \N__46724\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_14_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21836\,
            in2 => \N__24887\,
            in3 => \N__20876\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            clk => \N__47303\,
            ce => \N__23637\,
            sr => \N__46724\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_15_LC_4_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21749\,
            in2 => \N__24836\,
            in3 => \N__21185\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            clk => \N__47303\,
            ce => \N__23637\,
            sr => \N__46724\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_16_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24754\,
            in2 => \N__21800\,
            in3 => \N__21170\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_4_15_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            clk => \N__47294\,
            ce => \N__23676\,
            sr => \N__46728\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_17_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24683\,
            in2 => \N__21512\,
            in3 => \N__21158\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            clk => \N__47294\,
            ce => \N__23676\,
            sr => \N__46728\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_18_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21938\,
            in2 => \N__24620\,
            in3 => \N__21143\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            clk => \N__47294\,
            ce => \N__23676\,
            sr => \N__46728\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_19_LC_4_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24539\,
            in2 => \N__21743\,
            in3 => \N__21125\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            clk => \N__47294\,
            ce => \N__23676\,
            sr => \N__46728\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_20_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21830\,
            in2 => \N__25469\,
            in3 => \N__21110\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            clk => \N__47294\,
            ce => \N__23676\,
            sr => \N__46728\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_21_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21791\,
            in2 => \N__25403\,
            in3 => \N__21098\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            clk => \N__47294\,
            ce => \N__23676\,
            sr => \N__46728\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_22_LC_4_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25322\,
            in2 => \N__21923\,
            in3 => \N__21077\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            clk => \N__47294\,
            ce => \N__23676\,
            sr => \N__46728\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_23_LC_4_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25259\,
            in2 => \N__21932\,
            in3 => \N__21065\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            clk => \N__47294\,
            ce => \N__23676\,
            sr => \N__46728\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_24_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21914\,
            in2 => \N__25184\,
            in3 => \N__21374\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_4_16_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            clk => \N__47286\,
            ce => \N__23673\,
            sr => \N__46731\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_25_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25106\,
            in2 => \N__21906\,
            in3 => \N__21362\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            clk => \N__47286\,
            ce => \N__23673\,
            sr => \N__46731\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_26_LC_4_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21896\,
            in2 => \N__25055\,
            in3 => \N__21338\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            clk => \N__47286\,
            ce => \N__23673\,
            sr => \N__46731\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_27_LC_4_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25955\,
            in2 => \N__21907\,
            in3 => \N__21323\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            clk => \N__47286\,
            ce => \N__23673\,
            sr => \N__46731\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_28_LC_4_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21900\,
            in2 => \N__25906\,
            in3 => \N__21308\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            clk => \N__47286\,
            ce => \N__23673\,
            sr => \N__46731\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_29_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25848\,
            in2 => \N__21908\,
            in3 => \N__21293\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            clk => \N__47286\,
            ce => \N__23673\,
            sr => \N__46731\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_30_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21904\,
            in2 => \N__25791\,
            in3 => \N__21275\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\,
            clk => \N__47286\,
            ce => \N__23673\,
            sr => \N__46731\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_31_LC_4_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__21905\,
            in1 => \N__25658\,
            in2 => \_gnd_net_\,
            in3 => \N__21272\,
            lcout => \current_shift_inst.PI_CTRL.un8_enablelto31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47286\,
            ce => \N__23673\,
            sr => \N__46731\
        );

    \current_shift_inst.PI_CTRL.prop_term_12_LC_4_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23956\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47279\,
            ce => \N__23678\,
            sr => \N__46736\
        );

    \CONSTANT_ONE_LUT4_LC_4_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_7_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__21485\,
            in1 => \N__21713\,
            in2 => \N__21629\,
            in3 => \N__21655\,
            lcout => \counterZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47345\,
            ce => 'H',
            sr => \N__46671\
        );

    \counter_RNI800G_7_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21592\,
            in2 => \_gnd_net_\,
            in3 => \N__21478\,
            lcout => OPEN,
            ltout => \un2_counter_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNI3BSP_1_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__21465\,
            in1 => \N__21442\,
            in2 => \N__21431\,
            in3 => \N__21428\,
            lcout => un2_counter_9,
            ltout => \un2_counter_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_10khz_RNIIENA2_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__21869\,
            in1 => \N__21712\,
            in2 => \N__21404\,
            in3 => \N__21620\,
            lcout => \clk_10khz_RNIIENAZ0Z2\,
            ltout => \clk_10khz_RNIIENAZ0Z2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_cnv_0_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__34537\,
            in1 => \_gnd_net_\,
            in2 => \N__21401\,
            in3 => \N__21870\,
            lcout => \N_702_g\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_10khz_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__21621\,
            in1 => \N__21871\,
            in2 => \N__21665\,
            in3 => \N__21715\,
            lcout => clk_10khz_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47345\,
            ce => 'H',
            sr => \N__46671\
        );

    \pwm_generator_inst.threshold_2_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21398\,
            lcout => \pwm_generator_inst.thresholdZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47341\,
            ce => 'H',
            sr => \N__46679\
        );

    \counter_10_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__21719\,
            in1 => \N__21680\,
            in2 => \N__21666\,
            in3 => \N__21628\,
            lcout => \counterZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47341\,
            ce => 'H',
            sr => \N__46679\
        );

    \pwm_generator_inst.threshold_8_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21581\,
            lcout => \pwm_generator_inst.thresholdZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47331\,
            ce => 'H',
            sr => \N__46696\
        );

    \current_shift_inst.PI_CTRL.prop_term_1_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23864\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47323\,
            ce => \N__23585\,
            sr => \N__46705\
        );

    \current_shift_inst.PI_CTRL.prop_term_11_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24032\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47316\,
            ce => \N__23635\,
            sr => \N__46709\
        );

    \current_shift_inst.PI_CTRL.prop_term_9_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24170\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47316\,
            ce => \N__23635\,
            sr => \N__46709\
        );

    \current_shift_inst.PI_CTRL.prop_term_5_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24443\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47316\,
            ce => \N__23635\,
            sr => \N__46709\
        );

    \current_shift_inst.PI_CTRL.prop_term_0_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23911\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47304\,
            ce => \N__23641\,
            sr => \N__46713\
        );

    \current_shift_inst.PI_CTRL.prop_term_4_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23461\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47304\,
            ce => \N__23641\,
            sr => \N__46713\
        );

    \current_shift_inst.PI_CTRL.prop_term_17_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24659\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47304\,
            ce => \N__23641\,
            sr => \N__46713\
        );

    \current_shift_inst.PI_CTRL.prop_term_2_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23806\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47304\,
            ce => \N__23641\,
            sr => \N__46713\
        );

    \current_shift_inst.PI_CTRL.prop_term_8_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24236\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47304\,
            ce => \N__23641\,
            sr => \N__46713\
        );

    \current_shift_inst.PI_CTRL.prop_term_6_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24364\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47304\,
            ce => \N__23641\,
            sr => \N__46713\
        );

    \current_shift_inst.PI_CTRL.prop_term_3_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23734\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47304\,
            ce => \N__23641\,
            sr => \N__46713\
        );

    \current_shift_inst.PI_CTRL.prop_term_15_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24797\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47295\,
            ce => \N__23636\,
            sr => \N__46721\
        );

    \current_shift_inst.PI_CTRL.prop_term_19_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24515\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47295\,
            ce => \N__23636\,
            sr => \N__46721\
        );

    \current_shift_inst.PI_CTRL.integrator_11_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000001100"
        )
    port map (
            in0 => \N__22726\,
            in1 => \N__25678\,
            in2 => \N__22625\,
            in3 => \N__24002\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47295\,
            ce => \N__23636\,
            sr => \N__46721\
        );

    \current_shift_inst.PI_CTRL.prop_term_10_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24100\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47295\,
            ce => \N__23636\,
            sr => \N__46721\
        );

    \current_shift_inst.PI_CTRL.prop_term_13_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24946\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47295\,
            ce => \N__23636\,
            sr => \N__46721\
        );

    \current_shift_inst.PI_CTRL.prop_term_14_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24911\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47295\,
            ce => \N__23636\,
            sr => \N__46721\
        );

    \current_shift_inst.PI_CTRL.prop_term_20_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25442\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47295\,
            ce => \N__23636\,
            sr => \N__46721\
        );

    \current_shift_inst.PI_CTRL.integrator_10_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100011111000"
        )
    port map (
            in0 => \N__24077\,
            in1 => \N__22725\,
            in2 => \N__25682\,
            in3 => \N__22619\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47295\,
            ce => \N__23636\,
            sr => \N__46721\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25907\,
            in1 => \N__25954\,
            in2 => \N__25787\,
            in3 => \N__23990\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_10_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIA53P2_10_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21818\,
            in1 => \N__21812\,
            in2 => \N__21821\,
            in3 => \N__21806\,
            lcout => \current_shift_inst.PI_CTRL.N_47_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25105\,
            in1 => \N__25180\,
            in2 => \N__25054\,
            in3 => \N__25396\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_11_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24875\,
            in1 => \N__24982\,
            in2 => \N__24755\,
            in3 => \N__24050\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_9_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIB98M_0_10_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25257\,
            in1 => \N__24825\,
            in2 => \N__25853\,
            in3 => \N__24119\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_8_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_16_LC_5_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24718\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47280\,
            ce => \N__23675\,
            sr => \N__46729\
        );

    \current_shift_inst.PI_CTRL.prop_term_21_LC_5_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25361\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47280\,
            ce => \N__23675\,
            sr => \N__46729\
        );

    \current_shift_inst.PI_CTRL.prop_term_18_LC_5_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24577\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47280\,
            ce => \N__23675\,
            sr => \N__46729\
        );

    \current_shift_inst.PI_CTRL.integrator_30_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010110000"
        )
    port map (
            in0 => \N__25745\,
            in1 => \N__22614\,
            in2 => \N__25677\,
            in3 => \N__22741\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47280\,
            ce => \N__23675\,
            sr => \N__46729\
        );

    \current_shift_inst.PI_CTRL.prop_term_23_LC_5_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25222\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47280\,
            ce => \N__23675\,
            sr => \N__46729\
        );

    \current_shift_inst.PI_CTRL.integrator_4_LC_5_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011101100"
        )
    port map (
            in0 => \N__22742\,
            in1 => \N__25654\,
            in2 => \N__23438\,
            in3 => \N__22615\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47280\,
            ce => \N__23675\,
            sr => \N__46729\
        );

    \current_shift_inst.PI_CTRL.prop_term_22_LC_5_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25288\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47280\,
            ce => \N__23675\,
            sr => \N__46729\
        );

    \current_shift_inst.PI_CTRL.prop_term_24_LC_5_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25144\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47267\,
            ce => \N__23677\,
            sr => \N__46732\
        );

    \current_shift_inst.PI_CTRL.prop_term_25_LC_5_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25730\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47267\,
            ce => \N__23677\,
            sr => \N__46732\
        );

    \current_shift_inst.phase_valid_RNISLOR2_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__32393\,
            in1 => \N__21875\,
            in2 => \N__34536\,
            in3 => \N__21854\,
            lcout => \current_shift_inst.phase_valid_RNISLORZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_7_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21845\,
            lcout => \pwm_generator_inst.thresholdZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47332\,
            ce => 'H',
            sr => \N__46660\
        );

    \pwm_generator_inst.threshold_1_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21977\,
            lcout => \pwm_generator_inst.thresholdZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47332\,
            ce => 'H',
            sr => \N__46660\
        );

    \pwm_generator_inst.threshold_4_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21965\,
            lcout => \pwm_generator_inst.thresholdZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47324\,
            ce => 'H',
            sr => \N__46672\
        );

    \pwm_generator_inst.threshold_9_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21956\,
            lcout => \pwm_generator_inst.thresholdZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47317\,
            ce => 'H',
            sr => \N__46680\
        );

    \phase_controller_inst1.stoper_hc.target_time_8_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__44157\,
            in1 => \N__41768\,
            in2 => \_gnd_net_\,
            in3 => \N__43851\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47305\,
            ce => \N__31226\,
            sr => \N__46686\
        );

    \current_shift_inst.PI_CTRL.integrator_5_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000101010001111"
        )
    port map (
            in0 => \N__24413\,
            in1 => \N__22604\,
            in2 => \N__25676\,
            in3 => \N__22739\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47296\,
            ce => \N__23679\,
            sr => \N__46697\
        );

    \current_shift_inst.PI_CTRL.integrator_6_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001100010001"
        )
    port map (
            in0 => \N__22740\,
            in1 => \N__25649\,
            in2 => \N__22624\,
            in3 => \N__24338\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47296\,
            ce => \N__23679\,
            sr => \N__46697\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001101"
        )
    port map (
            in0 => \N__23710\,
            in1 => \N__22406\,
            in2 => \N__23498\,
            in3 => \N__22049\,
            lcout => \current_shift_inst.PI_CTRL.N_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24190\,
            in1 => \N__24290\,
            in2 => \N__24465\,
            in3 => \N__24386\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__23709\,
            in1 => \N__23493\,
            in2 => \N__21941\,
            in3 => \N__24255\,
            lcout => \current_shift_inst.PI_CTRL.N_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIB4HQ_8_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24189\,
            in2 => \_gnd_net_\,
            in3 => \N__24254\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI4JA22_5_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__24459\,
            in1 => \N__24291\,
            in2 => \N__22052\,
            in3 => \N__24387\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIOU8U3_18_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24610\,
            in1 => \N__22447\,
            in2 => \N__25675\,
            in3 => \N__21988\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIE7HME_18_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__21998\,
            in1 => \N__22018\,
            in2 => \N__22043\,
            in3 => \N__22040\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNITMGQ3_18_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__24611\,
            in1 => \N__25632\,
            in2 => \N__22465\,
            in3 => \N__22033\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24880\,
            in1 => \N__24972\,
            in2 => \N__24753\,
            in3 => \N__24063\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIBHHP7_18_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__22034\,
            in1 => \N__24612\,
            in2 => \N__22466\,
            in3 => \N__22019\,
            lcout => \current_shift_inst.PI_CTRL.N_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25250\,
            in1 => \N__24821\,
            in2 => \N__25852\,
            in3 => \N__24127\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIA53P2_0_10_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22073\,
            in1 => \N__22082\,
            in2 => \N__22007\,
            in3 => \N__22004\,
            lcout => \current_shift_inst.PI_CTRL.N_46_21\,
            ltout => \current_shift_inst.PI_CTRL.N_46_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI1IOH6_18_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24613\,
            in1 => \N__22448\,
            in2 => \N__21992\,
            in3 => \N__21989\,
            lcout => \current_shift_inst.PI_CTRL.N_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25886\,
            in1 => \N__25946\,
            in2 => \N__25795\,
            in3 => \N__23981\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25091\,
            in1 => \N__25166\,
            in2 => \N__25040\,
            in3 => \N__25385\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_15_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110011010000"
        )
    port map (
            in0 => \N__22551\,
            in1 => \N__24770\,
            in2 => \N__25667\,
            in3 => \N__22689\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47268\,
            ce => \N__23683\,
            sr => \N__46714\
        );

    \current_shift_inst.PI_CTRL.integrator_23_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011101100"
        )
    port map (
            in0 => \N__22690\,
            in1 => \N__25614\,
            in2 => \N__25202\,
            in3 => \N__22552\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47268\,
            ce => \N__23683\,
            sr => \N__46714\
        );

    \current_shift_inst.PI_CTRL.integrator_27_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010110000"
        )
    port map (
            in0 => \N__25922\,
            in1 => \N__22591\,
            in2 => \N__25666\,
            in3 => \N__22735\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47259\,
            ce => \N__23671\,
            sr => \N__46722\
        );

    \current_shift_inst.PI_CTRL.integrator_28_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111110001000"
        )
    port map (
            in0 => \N__22736\,
            in1 => \N__25865\,
            in2 => \N__22621\,
            in3 => \N__25613\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47259\,
            ce => \N__23671\,
            sr => \N__46722\
        );

    \current_shift_inst.PI_CTRL.integrator_26_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010110000"
        )
    port map (
            in0 => \N__25007\,
            in1 => \N__22590\,
            in2 => \N__25665\,
            in3 => \N__22734\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47259\,
            ce => \N__23671\,
            sr => \N__46722\
        );

    \current_shift_inst.PI_CTRL.integrator_31_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000001100"
        )
    port map (
            in0 => \N__22738\,
            in1 => \N__25603\,
            in2 => \N__22623\,
            in3 => \N__25490\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47259\,
            ce => \N__23671\,
            sr => \N__46722\
        );

    \current_shift_inst.PI_CTRL.prop_term_7_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24316\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47259\,
            ce => \N__23671\,
            sr => \N__46722\
        );

    \current_shift_inst.PI_CTRL.integrator_29_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000001100"
        )
    port map (
            in0 => \N__22737\,
            in1 => \N__25602\,
            in2 => \N__22622\,
            in3 => \N__25808\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47259\,
            ce => \N__23671\,
            sr => \N__46722\
        );

    \current_shift_inst.PI_CTRL.integrator_24_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010110000"
        )
    port map (
            in0 => \N__25118\,
            in1 => \N__22589\,
            in2 => \N__25664\,
            in3 => \N__22732\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47259\,
            ce => \N__23671\,
            sr => \N__46722\
        );

    \current_shift_inst.PI_CTRL.integrator_25_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000001100"
        )
    port map (
            in0 => \N__22733\,
            in1 => \N__25601\,
            in2 => \N__22620\,
            in3 => \N__25070\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47259\,
            ce => \N__23671\,
            sr => \N__46722\
        );

    \current_shift_inst.control_input_0_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22751\,
            in2 => \N__31417\,
            in3 => \N__31418\,
            lcout => \current_shift_inst.control_inputZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_7_17_0_\,
            carryout => \current_shift_inst.control_input_1_cry_0\,
            clk => \N__47251\,
            ce => \N__23027\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_1_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22871\,
            in2 => \_gnd_net_\,
            in3 => \N__22100\,
            lcout => \current_shift_inst.control_inputZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_0\,
            carryout => \current_shift_inst.control_input_1_cry_1\,
            clk => \N__47251\,
            ce => \N__23027\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_2_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22862\,
            in2 => \_gnd_net_\,
            in3 => \N__22097\,
            lcout => \current_shift_inst.control_inputZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_1\,
            carryout => \current_shift_inst.control_input_1_cry_2\,
            clk => \N__47251\,
            ce => \N__23027\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_3_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22853\,
            in2 => \_gnd_net_\,
            in3 => \N__22094\,
            lcout => \current_shift_inst.control_inputZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_2\,
            carryout => \current_shift_inst.control_input_1_cry_3\,
            clk => \N__47251\,
            ce => \N__23027\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_4_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22844\,
            in2 => \_gnd_net_\,
            in3 => \N__22091\,
            lcout => \current_shift_inst.control_inputZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_3\,
            carryout => \current_shift_inst.control_input_1_cry_4\,
            clk => \N__47251\,
            ce => \N__23027\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_5_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22835\,
            in2 => \_gnd_net_\,
            in3 => \N__22088\,
            lcout => \current_shift_inst.control_inputZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_4\,
            carryout => \current_shift_inst.control_input_1_cry_5\,
            clk => \N__47251\,
            ce => \N__23027\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_6_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22826\,
            in2 => \_gnd_net_\,
            in3 => \N__22085\,
            lcout => \current_shift_inst.control_inputZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_5\,
            carryout => \current_shift_inst.control_input_1_cry_6\,
            clk => \N__47251\,
            ce => \N__23027\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_7_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22817\,
            in2 => \_gnd_net_\,
            in3 => \N__22127\,
            lcout => \current_shift_inst.control_inputZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_6\,
            carryout => \current_shift_inst.control_input_1_cry_7\,
            clk => \N__47251\,
            ce => \N__23027\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_8_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22796\,
            in2 => \_gnd_net_\,
            in3 => \N__22124\,
            lcout => \current_shift_inst.control_inputZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_7_18_0_\,
            carryout => \current_shift_inst.control_input_1_cry_8\,
            clk => \N__47243\,
            ce => \N__23026\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_9_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22988\,
            in2 => \_gnd_net_\,
            in3 => \N__22121\,
            lcout => \current_shift_inst.control_inputZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_8\,
            carryout => \current_shift_inst.control_input_1_cry_9\,
            clk => \N__47243\,
            ce => \N__23026\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_10_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22979\,
            in2 => \_gnd_net_\,
            in3 => \N__22118\,
            lcout => \current_shift_inst.control_inputZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_9\,
            carryout => \current_shift_inst.control_input_1_cry_10\,
            clk => \N__47243\,
            ce => \N__23026\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_11_LC_7_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22970\,
            in2 => \_gnd_net_\,
            in3 => \N__22115\,
            lcout => \current_shift_inst.control_inputZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_10\,
            carryout => \current_shift_inst.control_input_1_cry_11\,
            clk => \N__47243\,
            ce => \N__23026\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_12_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22949\,
            in2 => \_gnd_net_\,
            in3 => \N__22112\,
            lcout => \current_shift_inst.control_inputZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_11\,
            carryout => \current_shift_inst.control_input_1_cry_12\,
            clk => \N__47243\,
            ce => \N__23026\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_13_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22928\,
            in2 => \_gnd_net_\,
            in3 => \N__22109\,
            lcout => \current_shift_inst.control_inputZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_12\,
            carryout => \current_shift_inst.control_input_1_cry_13\,
            clk => \N__47243\,
            ce => \N__23026\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_14_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22907\,
            in2 => \_gnd_net_\,
            in3 => \N__22106\,
            lcout => \current_shift_inst.control_inputZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_13\,
            carryout => \current_shift_inst.control_input_1_cry_14\,
            clk => \N__47243\,
            ce => \N__23026\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_15_LC_7_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22898\,
            in2 => \_gnd_net_\,
            in3 => \N__22103\,
            lcout => \current_shift_inst.control_inputZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_14\,
            carryout => \current_shift_inst.control_input_1_cry_15\,
            clk => \N__47243\,
            ce => \N__23026\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_16_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22889\,
            in2 => \_gnd_net_\,
            in3 => \N__22154\,
            lcout => \current_shift_inst.control_inputZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_7_19_0_\,
            carryout => \current_shift_inst.control_input_1_cry_16\,
            clk => \N__47235\,
            ce => \N__23037\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_17_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22880\,
            in2 => \_gnd_net_\,
            in3 => \N__22151\,
            lcout => \current_shift_inst.control_inputZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_16\,
            carryout => \current_shift_inst.control_input_1_cry_17\,
            clk => \N__47235\,
            ce => \N__23037\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_18_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23117\,
            in2 => \_gnd_net_\,
            in3 => \N__22148\,
            lcout => \current_shift_inst.control_inputZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_17\,
            carryout => \current_shift_inst.control_input_1_cry_18\,
            clk => \N__47235\,
            ce => \N__23037\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_19_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23108\,
            in2 => \_gnd_net_\,
            in3 => \N__22145\,
            lcout => \current_shift_inst.control_inputZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_18\,
            carryout => \current_shift_inst.control_input_1_cry_19\,
            clk => \N__47235\,
            ce => \N__23037\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_20_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23099\,
            in2 => \_gnd_net_\,
            in3 => \N__22142\,
            lcout => \current_shift_inst.control_inputZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_19\,
            carryout => \current_shift_inst.control_input_1_cry_20\,
            clk => \N__47235\,
            ce => \N__23037\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_21_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23090\,
            in2 => \_gnd_net_\,
            in3 => \N__22139\,
            lcout => \current_shift_inst.control_inputZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_20\,
            carryout => \current_shift_inst.control_input_1_cry_21\,
            clk => \N__47235\,
            ce => \N__23037\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_22_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23081\,
            in2 => \_gnd_net_\,
            in3 => \N__22136\,
            lcout => \current_shift_inst.control_inputZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_21\,
            carryout => \current_shift_inst.control_input_1_cry_22\,
            clk => \N__47235\,
            ce => \N__23037\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_23_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23072\,
            in2 => \_gnd_net_\,
            in3 => \N__22133\,
            lcout => \current_shift_inst.control_inputZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_22\,
            carryout => \current_shift_inst.control_input_1_cry_23\,
            clk => \N__47235\,
            ce => \N__23037\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_24_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23063\,
            in2 => \_gnd_net_\,
            in3 => \N__22130\,
            lcout => \current_shift_inst.control_inputZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_7_20_0_\,
            carryout => \current_shift_inst.control_input_1_cry_24\,
            clk => \N__47228\,
            ce => \N__23038\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_1_cry_24_THRU_LUT4_0_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22226\,
            lcout => \current_shift_inst.control_input_1_cry_24_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MIN_D1_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22223\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_min_comp2_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MAX_D1_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22211\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_max_comp2_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47337\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_0_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22196\,
            lcout => \pwm_generator_inst.thresholdZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47325\,
            ce => 'H',
            sr => \N__46651\
        );

    \pwm_generator_inst.threshold_6_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22184\,
            lcout => \pwm_generator_inst.thresholdZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47318\,
            ce => 'H',
            sr => \N__46661\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__39678\,
            in1 => \N__39846\,
            in2 => \N__40006\,
            in3 => \N__28928\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47318\,
            ce => 'H',
            sr => \N__46661\
        );

    \pwm_generator_inst.threshold_3_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22172\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.thresholdZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47318\,
            ce => 'H',
            sr => \N__46661\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__39679\,
            in1 => \N__39847\,
            in2 => \N__40007\,
            in3 => \N__29237\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47318\,
            ce => 'H',
            sr => \N__46661\
        );

    \pwm_generator_inst.threshold_5_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22163\,
            lcout => \pwm_generator_inst.thresholdZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47306\,
            ce => 'H',
            sr => \N__46673\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010000010"
        )
    port map (
            in0 => \N__23921\,
            in1 => \N__39654\,
            in2 => \N__40018\,
            in3 => \N__39845\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47306\,
            ce => 'H',
            sr => \N__46673\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23381\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_11_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22322\,
            in2 => \N__22340\,
            in3 => \N__28377\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22298\,
            in2 => \N__22316\,
            in3 => \N__28354\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22274\,
            in2 => \N__22292\,
            in3 => \N__28312\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22268\,
            in2 => \N__23420\,
            in3 => \N__28279\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22262\,
            in2 => \N__23372\,
            in3 => \N__29074\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22238\,
            in2 => \N__22256\,
            in3 => \N__29041\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29008\,
            in1 => \N__22232\,
            in2 => \N__23930\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28978\,
            in1 => \N__22388\,
            in2 => \N__22400\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \bfn_8_12_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22382\,
            in2 => \N__27410\,
            in3 => \N__31142\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22376\,
            in2 => \N__23363\,
            in3 => \N__28945\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22370\,
            in2 => \N__27422\,
            in3 => \N__28916\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22364\,
            in2 => \N__23396\,
            in3 => \N__28886\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22358\,
            in2 => \N__23408\,
            in3 => \N__29282\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22352\,
            in2 => \N__27437\,
            in3 => \N__29254\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29225\,
            in1 => \N__22346\,
            in2 => \N__29354\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22433\,
            in2 => \N__31268\,
            in3 => \N__29198\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \bfn_8_13_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22427\,
            in2 => \N__31256\,
            in3 => \N__29171\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22421\,
            in2 => \N__29342\,
            in3 => \N__29144\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22415\,
            in2 => \N__31244\,
            in3 => \N__29117\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22409\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__23880\,
            in1 => \N__23778\,
            in2 => \_gnd_net_\,
            in3 => \N__23830\,
            lcout => \current_shift_inst.PI_CTRL.un1_enablelt3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__39769\,
            in1 => \N__39962\,
            in2 => \_gnd_net_\,
            in3 => \N__39610\,
            lcout => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_18_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000001100"
        )
    port map (
            in0 => \N__22684\,
            in1 => \N__25634\,
            in2 => \N__22609\,
            in3 => \N__24551\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47269\,
            ce => \N__23631\,
            sr => \N__46706\
        );

    \current_shift_inst.PI_CTRL.integrator_9_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000101010001111"
        )
    port map (
            in0 => \N__24140\,
            in1 => \N__22555\,
            in2 => \N__25674\,
            in3 => \N__22688\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47269\,
            ce => \N__23631\,
            sr => \N__46706\
        );

    \current_shift_inst.PI_CTRL.integrator_7_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100000011011101"
        )
    port map (
            in0 => \N__22686\,
            in1 => \N__24272\,
            in2 => \N__22611\,
            in3 => \N__25645\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47269\,
            ce => \N__23631\,
            sr => \N__46706\
        );

    \current_shift_inst.PI_CTRL.integrator_8_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000101010001111"
        )
    port map (
            in0 => \N__24206\,
            in1 => \N__22554\,
            in2 => \N__25673\,
            in3 => \N__22687\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47269\,
            ce => \N__23631\,
            sr => \N__46706\
        );

    \current_shift_inst.PI_CTRL.integrator_21_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000001100"
        )
    port map (
            in0 => \N__22685\,
            in1 => \N__25635\,
            in2 => \N__22610\,
            in3 => \N__25331\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47269\,
            ce => \N__23631\,
            sr => \N__46706\
        );

    \current_shift_inst.PI_CTRL.integrator_12_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010110000"
        )
    port map (
            in0 => \N__24992\,
            in1 => \N__22553\,
            in2 => \N__25672\,
            in3 => \N__22682\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47269\,
            ce => \N__23631\,
            sr => \N__46706\
        );

    \current_shift_inst.PI_CTRL.integrator_13_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000001100"
        )
    port map (
            in0 => \N__22683\,
            in1 => \N__25633\,
            in2 => \N__22608\,
            in3 => \N__24923\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47269\,
            ce => \N__23631\,
            sr => \N__46706\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25460\,
            in1 => \N__24533\,
            in2 => \N__25320\,
            in3 => \N__24677\,
            lcout => \current_shift_inst.PI_CTRL.N_47_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_17_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100011111000"
        )
    port map (
            in0 => \N__22721\,
            in1 => \N__24629\,
            in2 => \N__25669\,
            in3 => \N__22575\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47260\,
            ce => \N__23684\,
            sr => \N__46710\
        );

    \current_shift_inst.PI_CTRL.integrator_19_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111010001100"
        )
    port map (
            in0 => \N__24485\,
            in1 => \N__25619\,
            in2 => \N__22613\,
            in3 => \N__22722\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47260\,
            ce => \N__23684\,
            sr => \N__46710\
        );

    \current_shift_inst.PI_CTRL.integrator_20_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100011111000"
        )
    port map (
            in0 => \N__22723\,
            in1 => \N__25412\,
            in2 => \N__25670\,
            in3 => \N__22576\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47260\,
            ce => \N__23684\,
            sr => \N__46710\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25461\,
            in1 => \N__24534\,
            in2 => \N__25321\,
            in3 => \N__24678\,
            lcout => \current_shift_inst.PI_CTRL.N_46_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_22_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100011111000"
        )
    port map (
            in0 => \N__22724\,
            in1 => \N__25268\,
            in2 => \N__25671\,
            in3 => \N__22577\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47260\,
            ce => \N__23684\,
            sr => \N__46710\
        );

    \current_shift_inst.PI_CTRL.integrator_14_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111010001100"
        )
    port map (
            in0 => \N__24845\,
            in1 => \N__25618\,
            in2 => \N__22612\,
            in3 => \N__22719\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47260\,
            ce => \N__23684\,
            sr => \N__46710\
        );

    \current_shift_inst.PI_CTRL.integrator_16_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100011111000"
        )
    port map (
            in0 => \N__22720\,
            in1 => \N__24692\,
            in2 => \N__25668\,
            in3 => \N__22574\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47260\,
            ce => \N__23684\,
            sr => \N__46710\
        );

    \current_shift_inst.un38_control_input_0_cry_5_c_RNO_0_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27487\,
            in2 => \_gnd_net_\,
            in3 => \N__29530\,
            lcout => \current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4H5J_19_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__30417\,
            in1 => \N__30463\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI4H5J_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIH6661_17_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__28001\,
            in1 => \N__29640\,
            in2 => \N__29684\,
            in3 => \N__27949\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIH6661_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR0UI_13_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29968\,
            in2 => \_gnd_net_\,
            in3 => \N__29929\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIR0UI_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQKU1_5_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__29488\,
            in1 => \N__27803\,
            in2 => \N__27857\,
            in3 => \N__29453\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIVQKU1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_5_c_RNO_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__27852\,
            in1 => \N__27488\,
            in2 => \N__29534\,
            in3 => \N__29487\,
            lcout => \current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAL3J_18_LC_8_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27948\,
            in2 => \_gnd_net_\,
            in3 => \N__29641\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIAL3J_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CRY_0_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30599\,
            in2 => \N__30605\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_17_0_\,
            carryout => \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_0_c_inv_LC_8_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22787\,
            in2 => \N__29306\,
            in3 => \N__31435\,
            lcout => \current_shift_inst.z_i_0_31\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CO\,
            carryout => \current_shift_inst.un38_control_input_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_1_c_LC_8_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25481\,
            in2 => \N__29615\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_0\,
            carryout => \current_shift_inst.un38_control_input_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_2_c_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29581\,
            in2 => \N__26033\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_1\,
            carryout => \current_shift_inst.un38_control_input_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_3_c_inv_LC_8_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25475\,
            in1 => \N__29555\,
            in2 => \N__22781\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un38_control_input_0_cry_3_c_invZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_2\,
            carryout => \current_shift_inst.un38_control_input_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_4_c_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26012\,
            in2 => \N__26024\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_3\,
            carryout => \current_shift_inst.un38_control_input_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_5_c_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22772\,
            in2 => \N__22766\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_4\,
            carryout => \current_shift_inst.un38_control_input_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_5_c_RNI7HN13_LC_8_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22757\,
            in2 => \N__25991\,
            in3 => \N__22745\,
            lcout => \current_shift_inst.control_input_1_axb_0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_5\,
            carryout => \current_shift_inst.un38_control_input_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_6_c_RNIHVR13_LC_8_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26090\,
            in2 => \N__25967\,
            in3 => \N__22865\,
            lcout => \current_shift_inst.control_input_1_axb_1\,
            ltout => OPEN,
            carryin => \bfn_8_18_0_\,
            carryout => \current_shift_inst.un38_control_input_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_7_c_RNIRD023_LC_8_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26051\,
            in2 => \N__26006\,
            in3 => \N__22856\,
            lcout => \current_shift_inst.control_input_1_axb_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_7\,
            carryout => \current_shift_inst.un38_control_input_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_8_c_RNIC9753_LC_8_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30002\,
            in2 => \N__29807\,
            in3 => \N__22847\,
            lcout => \current_shift_inst.control_input_1_axb_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_8\,
            carryout => \current_shift_inst.un38_control_input_0_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_9_c_RNII9PR2_LC_8_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26045\,
            in2 => \N__25982\,
            in3 => \N__22838\,
            lcout => \current_shift_inst.control_input_1_axb_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_9\,
            carryout => \current_shift_inst.un38_control_input_0_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_10_c_RNIV96V1_LC_8_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26096\,
            in2 => \N__26078\,
            in3 => \N__22829\,
            lcout => \current_shift_inst.control_input_1_axb_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_10\,
            carryout => \current_shift_inst.un38_control_input_0_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_11_c_RNI9OAV1_LC_8_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30647\,
            in2 => \N__29993\,
            in3 => \N__22820\,
            lcout => \current_shift_inst.control_input_1_axb_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_11\,
            carryout => \current_shift_inst.un38_control_input_0_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_12_c_RNIJ6FV1_LC_8_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29891\,
            in2 => \N__29981\,
            in3 => \N__22811\,
            lcout => \current_shift_inst.control_input_1_axb_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_12\,
            carryout => \current_shift_inst.un38_control_input_0_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_13_c_RNITKJV1_LC_8_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25997\,
            in2 => \N__22808\,
            in3 => \N__22790\,
            lcout => \current_shift_inst.control_input_1_axb_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_13\,
            carryout => \current_shift_inst.un38_control_input_0_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_14_c_RNI73OV1_LC_8_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30137\,
            in2 => \N__26066\,
            in3 => \N__22982\,
            lcout => \current_shift_inst.control_input_1_axb_9\,
            ltout => OPEN,
            carryin => \bfn_8_19_0_\,
            carryout => \current_shift_inst.un38_control_input_0_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_15_c_RNIHHSV1_LC_8_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30287\,
            in2 => \N__30374\,
            in3 => \N__22973\,
            lcout => \current_shift_inst.control_input_1_axb_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_15\,
            carryout => \current_shift_inst.un38_control_input_0_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_16_c_RNIRV002_LC_8_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26057\,
            in2 => \N__26117\,
            in3 => \N__22964\,
            lcout => \current_shift_inst.control_input_1_axb_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_16\,
            carryout => \current_shift_inst.un38_control_input_0_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_17_c_RNI5E502_LC_8_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26084\,
            in2 => \N__22961\,
            in3 => \N__22943\,
            lcout => \current_shift_inst.control_input_1_axb_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_17\,
            carryout => \current_shift_inst.un38_control_input_0_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_18_c_RNI6KA02_LC_8_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25973\,
            in2 => \N__22940\,
            in3 => \N__22922\,
            lcout => \current_shift_inst.control_input_1_axb_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_18\,
            carryout => \current_shift_inst.un38_control_input_0_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_19_c_RNICO912_LC_8_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30383\,
            in2 => \N__22919\,
            in3 => \N__22901\,
            lcout => \current_shift_inst.control_input_1_axb_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_19\,
            carryout => \current_shift_inst.un38_control_input_0_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_20_c_RNI92P32_LC_8_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31085\,
            in2 => \N__31019\,
            in3 => \N__22892\,
            lcout => \current_shift_inst.control_input_1_axb_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_20\,
            carryout => \current_shift_inst.un38_control_input_0_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_21_c_RNIJGT32_LC_8_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26141\,
            in2 => \N__30938\,
            in3 => \N__22883\,
            lcout => \current_shift_inst.control_input_1_axb_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_21\,
            carryout => \current_shift_inst.un38_control_input_0_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_22_c_RNITU142_LC_8_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26147\,
            in2 => \N__26156\,
            in3 => \N__22874\,
            lcout => \current_shift_inst.control_input_1_axb_17\,
            ltout => OPEN,
            carryin => \bfn_8_20_0_\,
            carryout => \current_shift_inst.un38_control_input_0_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_23_c_RNI7D642_LC_8_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31481\,
            in2 => \N__30923\,
            in3 => \N__23111\,
            lcout => \current_shift_inst.control_input_1_axb_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_23\,
            carryout => \current_shift_inst.un38_control_input_0_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_24_c_RNIHRA42_LC_8_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30785\,
            in2 => \N__31886\,
            in3 => \N__23102\,
            lcout => \current_shift_inst.control_input_1_axb_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_24\,
            carryout => \current_shift_inst.un38_control_input_0_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_25_c_RNIR9F42_LC_8_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31796\,
            in2 => \N__31730\,
            in3 => \N__23093\,
            lcout => \current_shift_inst.control_input_1_axb_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_25\,
            carryout => \current_shift_inst.un38_control_input_0_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_26_c_RNI5OJ42_LC_8_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26102\,
            in2 => \N__30911\,
            in3 => \N__23084\,
            lcout => \current_shift_inst.control_input_1_axb_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_26\,
            carryout => \current_shift_inst.un38_control_input_0_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_27_c_RNIF6O42_LC_8_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26039\,
            in2 => \N__26126\,
            in3 => \N__23075\,
            lcout => \current_shift_inst.control_input_1_axb_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_27\,
            carryout => \current_shift_inst.un38_control_input_0_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_28_c_RNIGCT42_LC_8_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26108\,
            in2 => \N__30800\,
            in3 => \N__23066\,
            lcout => \current_shift_inst.control_input_1_axb_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_28\,
            carryout => \current_shift_inst.un38_control_input_0_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_29_c_RNIMGS52_LC_8_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26132\,
            in2 => \N__31654\,
            in3 => \N__23057\,
            lcout => \current_shift_inst.control_input_1_axb_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_29\,
            carryout => \current_shift_inst.un38_control_input_0_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_25_LC_8_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30476\,
            in2 => \N__23054\,
            in3 => \N__23045\,
            lcout => \current_shift_inst.control_inputZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47221\,
            ce => \N__23042\,
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MIN_D2_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23246\,
            lcout => \il_min_comp2_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47338\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MAX_D1_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23240\,
            lcout => \il_max_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47333\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23216\,
            in2 => \N__23225\,
            in3 => \N__27196\,
            lcout => \pwm_generator_inst.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_9_8_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27174\,
            in1 => \N__23210\,
            in2 => \N__23201\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_0\,
            carryout => \pwm_generator_inst.un14_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23180\,
            in2 => \N__23192\,
            in3 => \N__27154\,
            lcout => \pwm_generator_inst.counter_i_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_1\,
            carryout => \pwm_generator_inst.un14_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23174\,
            in2 => \N__23168\,
            in3 => \N__27132\,
            lcout => \pwm_generator_inst.counter_i_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_2\,
            carryout => \pwm_generator_inst.un14_counter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23159\,
            in2 => \N__23147\,
            in3 => \N__27111\,
            lcout => \pwm_generator_inst.counter_i_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_3\,
            carryout => \pwm_generator_inst.un14_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23123\,
            in2 => \N__23135\,
            in3 => \N__27090\,
            lcout => \pwm_generator_inst.counter_i_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_4\,
            carryout => \pwm_generator_inst.un14_counter_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23339\,
            in2 => \N__23351\,
            in3 => \N__27345\,
            lcout => \pwm_generator_inst.counter_i_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_5\,
            carryout => \pwm_generator_inst.un14_counter_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23333\,
            in2 => \N__23324\,
            in3 => \N__27324\,
            lcout => \pwm_generator_inst.counter_i_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_6\,
            carryout => \pwm_generator_inst.un14_counter_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23300\,
            in2 => \N__23315\,
            in3 => \N__27303\,
            lcout => \pwm_generator_inst.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_9_9_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23279\,
            in2 => \N__23294\,
            in3 => \N__27228\,
            lcout => \pwm_generator_inst.counter_i_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_8\,
            carryout => \pwm_generator_inst.un14_counter_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.pwm_out_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23273\,
            lcout => pwm_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47307\,
            ce => 'H',
            sr => \N__46652\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__39823\,
            in1 => \N__39661\,
            in2 => \N__40017\,
            in3 => \N__29030\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47297\,
            ce => 'H',
            sr => \N__46662\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__39658\,
            in1 => \N__40002\,
            in2 => \N__39854\,
            in3 => \N__28964\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47297\,
            ce => 'H',
            sr => \N__46662\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__39822\,
            in1 => \N__39660\,
            in2 => \N__40016\,
            in3 => \N__29063\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47297\,
            ce => 'H',
            sr => \N__46662\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__39656\,
            in1 => \N__39994\,
            in2 => \N__39852\,
            in3 => \N__28268\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47297\,
            ce => 'H',
            sr => \N__46662\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__39657\,
            in1 => \N__40001\,
            in2 => \N__39853\,
            in3 => \N__28997\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47297\,
            ce => 'H',
            sr => \N__46662\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__39821\,
            in1 => \N__39659\,
            in2 => \N__40015\,
            in3 => \N__28301\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47297\,
            ce => 'H',
            sr => \N__46662\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__39655\,
            in1 => \N__39990\,
            in2 => \N__39851\,
            in3 => \N__28343\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47297\,
            ce => 'H',
            sr => \N__46662\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__43848\,
            in1 => \N__35432\,
            in2 => \N__44186\,
            in3 => \N__40346\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47287\,
            ce => \N__31227\,
            sr => \N__46674\
        );

    \phase_controller_inst1.stoper_hc.target_time_13_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__44281\,
            in1 => \N__44144\,
            in2 => \_gnd_net_\,
            in3 => \N__43847\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47287\,
            ce => \N__31227\,
            sr => \N__46674\
        );

    \phase_controller_inst1.stoper_hc.target_time_12_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__43846\,
            in1 => \_gnd_net_\,
            in2 => \N__44185\,
            in3 => \N__39407\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47287\,
            ce => \N__31227\,
            sr => \N__46674\
        );

    \phase_controller_inst1.stoper_hc.target_time_0_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__40345\,
            in1 => \N__43844\,
            in2 => \N__42260\,
            in3 => \N__44139\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47287\,
            ce => \N__31227\,
            sr => \N__46674\
        );

    \phase_controller_inst1.stoper_hc.target_time_5_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100000001000"
        )
    port map (
            in0 => \N__43849\,
            in1 => \N__43956\,
            in2 => \N__44187\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47287\,
            ce => \N__31227\,
            sr => \N__46674\
        );

    \phase_controller_inst1.stoper_hc.target_time_10_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__35678\,
            in1 => \N__44140\,
            in2 => \_gnd_net_\,
            in3 => \N__43845\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47287\,
            ce => \N__31227\,
            sr => \N__46674\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__43850\,
            in1 => \_gnd_net_\,
            in2 => \N__44188\,
            in3 => \N__41670\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47287\,
            ce => \N__31227\,
            sr => \N__46674\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__40040\,
            in1 => \N__27393\,
            in2 => \_gnd_net_\,
            in3 => \N__28387\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27389\,
            in2 => \_gnd_net_\,
            in3 => \N__40039\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_0_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23881\,
            in2 => \N__23912\,
            in3 => \N__23755\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_9_13_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_0\,
            clk => \N__47270\,
            ce => \N__23674\,
            sr => \N__46687\
        );

    \current_shift_inst.PI_CTRL.integrator_1_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__23753\,
            in1 => \N__23829\,
            in2 => \N__23863\,
            in3 => \N__23810\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\,
            clk => \N__47270\,
            ce => \N__23674\,
            sr => \N__46687\
        );

    \current_shift_inst.PI_CTRL.integrator_2_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__23756\,
            in1 => \N__23779\,
            in2 => \N__23807\,
            in3 => \N__23759\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\,
            clk => \N__47270\,
            ce => \N__23674\,
            sr => \N__46687\
        );

    \current_shift_inst.PI_CTRL.integrator_3_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1101011101111101"
        )
    port map (
            in0 => \N__23754\,
            in1 => \N__23708\,
            in2 => \N__23735\,
            in3 => \N__23687\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\,
            clk => \N__47270\,
            ce => \N__23674\,
            sr => \N__46687\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23489\,
            in2 => \N__23462\,
            in3 => \N__23423\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24472\,
            in2 => \N__24442\,
            in3 => \N__24401\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24394\,
            in2 => \N__24365\,
            in3 => \N__24326\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24323\,
            in2 => \N__24298\,
            in3 => \N__24263\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24256\,
            in2 => \N__24235\,
            in3 => \N__24200\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \bfn_9_14_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24188\,
            in2 => \N__24169\,
            in3 => \N__24134\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24131\,
            in2 => \N__24101\,
            in3 => \N__24068\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24065\,
            in2 => \N__24031\,
            in3 => \N__23993\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23988\,
            in2 => \N__23957\,
            in3 => \N__24986\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24971\,
            in2 => \N__24947\,
            in3 => \N__24914\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24910\,
            in2 => \N__24879\,
            in3 => \N__24839\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24832\,
            in2 => \N__24796\,
            in3 => \N__24758\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24746\,
            in2 => \N__24719\,
            in3 => \N__24686\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \bfn_9_15_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24679\,
            in2 => \N__24658\,
            in3 => \N__24623\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24599\,
            in2 => \N__24578\,
            in3 => \N__24542\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24535\,
            in2 => \N__24514\,
            in3 => \N__24479\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25462\,
            in2 => \N__25441\,
            in3 => \N__25406\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25386\,
            in2 => \N__25360\,
            in3 => \N__25325\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25316\,
            in2 => \N__25292\,
            in3 => \N__25262\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25258\,
            in2 => \N__25226\,
            in3 => \N__25187\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25176\,
            in2 => \N__25145\,
            in3 => \N__25109\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \bfn_9_16_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25101\,
            in2 => \N__25731\,
            in3 => \N__25058\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25720\,
            in2 => \N__25050\,
            in3 => \N__24995\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25950\,
            in2 => \N__25732\,
            in3 => \N__25910\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25724\,
            in2 => \N__25905\,
            in3 => \N__25856\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25847\,
            in2 => \N__25733\,
            in3 => \N__25799\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25728\,
            in2 => \N__25796\,
            in3 => \N__25736\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__25729\,
            in1 => \N__25653\,
            in2 => \_gnd_net_\,
            in3 => \N__25493\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_1_c_RNO_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__30594\,
            in1 => \N__29614\,
            in2 => \_gnd_net_\,
            in3 => \N__27596\,
            lcout => \current_shift_inst.un38_control_input_0_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_2_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26423\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47236\,
            ce => \N__26477\,
            sr => \N__46715\
        );

    \current_shift_inst.un38_control_input_0_cry_3_c_inv_RNO_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101100101"
        )
    port map (
            in0 => \N__27526\,
            in1 => \N__27564\,
            in2 => \N__30603\,
            in3 => \N__27595\,
            lcout => \current_shift_inst.N_1717_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_1_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26456\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47236\,
            ce => \N__26477\,
            sr => \N__46715\
        );

    \current_shift_inst.un38_control_input_0_cry_2_c_RNO_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001101010011010"
        )
    port map (
            in0 => \N__27568\,
            in1 => \N__27597\,
            in2 => \N__30604\,
            in3 => \N__29582\,
            lcout => \current_shift_inst.un38_control_input_0_cry_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5LGN1_3_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__27598\,
            in1 => \N__27527\,
            in2 => \N__27569\,
            in3 => \N__30598\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3\,
            ltout => \current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_4_c_RNO_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27486\,
            in2 => \N__26015\,
            in3 => \N__29529\,
            lcout => \current_shift_inst.un38_control_input_0_cry_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIK3CV_7_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27758\,
            in3 => \N__29403\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIK3CV_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIP5T51_13_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__30271\,
            in1 => \N__29969\,
            in2 => \N__29933\,
            in3 => \N__30207\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIP5T51_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIER9V_5_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27853\,
            in2 => \_gnd_net_\,
            in3 => \N__29489\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIER9V_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJDBL1_10_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__27676\,
            in1 => \N__30074\,
            in2 => \N__30041\,
            in3 => \N__29736\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJDBL1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIE6961_18_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100110011001"
        )
    port map (
            in0 => \N__30462\,
            in1 => \N__30424\,
            in2 => \N__27953\,
            in3 => \N__29645\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIE6961_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHVAV_6_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__27798\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29451\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIHVAV_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7DM51_10_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \N__29737\,
            in1 => \N__27677\,
            in2 => \N__30773\,
            in3 => \N__30715\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI7DM51_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI53NU1_6_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001111000011"
        )
    port map (
            in0 => \N__27799\,
            in1 => \N__27752\,
            in2 => \N__29407\,
            in3 => \N__29452\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI53NU1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7H2J_17_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__29679\,
            in1 => \_gnd_net_\,
            in2 => \N__28000\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI7H2J_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIIKQI_10_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__27675\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29738\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIIKQI_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU4VI_14_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30270\,
            in2 => \_gnd_net_\,
            in3 => \N__30211\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIU4VI_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBU361_16_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__30320\,
            in1 => \N__27993\,
            in2 => \N__30358\,
            in3 => \N__29680\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIBU361_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBBPU1_7_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__27756\,
            in1 => \N__29846\,
            in2 => \N__29414\,
            in3 => \N__29880\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIBBPU1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1PG21_9_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30069\,
            in2 => \_gnd_net_\,
            in3 => \N__30037\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI1PG21_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNINKG81_27_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__28144\,
            in1 => \N__30879\,
            in2 => \N__30128\,
            in3 => \N__30838\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNINKG81_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR32K_22_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28249\,
            in2 => \_gnd_net_\,
            in3 => \N__29779\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIR32K_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPB581_22_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__28250\,
            in1 => \N__31544\,
            in2 => \N__29783\,
            in3 => \N__31588\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPB581_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJ3381_21_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__30968\,
            in1 => \N__28248\,
            in2 => \N__31007\,
            in3 => \N__29778\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJ3381_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQF91_30_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__31655\,
            in1 => \N__30631\,
            in2 => \_gnd_net_\,
            in3 => \N__30500\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIVQF91_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAO7K_27_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__30120\,
            in1 => \_gnd_net_\,
            in2 => \N__28145\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIAO7K_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4D1J_16_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30350\,
            in2 => \_gnd_net_\,
            in3 => \N__30319\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI4D1J_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIKKJ81_29_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__30883\,
            in1 => \N__31679\,
            in2 => \N__30842\,
            in3 => \N__31705\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIKKJ81_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHCE81_26_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__31866\,
            in1 => \N__28140\,
            in2 => \N__31832\,
            in3 => \N__30121\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIHCE81_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_3_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26455\,
            in2 => \N__26398\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_3\,
            ltout => OPEN,
            carryin => \bfn_9_21_0_\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_2\,
            clk => \N__47215\,
            ce => \N__26476\,
            sr => \N__46733\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_4_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26422\,
            in2 => \N__26371\,
            in3 => \N__26183\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_2\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_3\,
            clk => \N__47215\,
            ce => \N__26476\,
            sr => \N__46733\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_5_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26341\,
            in2 => \N__26399\,
            in3 => \N__26180\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_3\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_4\,
            clk => \N__47215\,
            ce => \N__26476\,
            sr => \N__46733\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_6_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26320\,
            in2 => \N__26372\,
            in3 => \N__26177\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_4\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_5\,
            clk => \N__47215\,
            ce => \N__26476\,
            sr => \N__46733\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_7_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26342\,
            in2 => \N__26297\,
            in3 => \N__26174\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_5\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_6\,
            clk => \N__47215\,
            ce => \N__26476\,
            sr => \N__46733\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_8_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26321\,
            in2 => \N__26263\,
            in3 => \N__26171\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_6\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_7\,
            clk => \N__47215\,
            ce => \N__26476\,
            sr => \N__46733\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_9_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26296\,
            in2 => \N__26696\,
            in3 => \N__26168\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_7\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_8\,
            clk => \N__47215\,
            ce => \N__26476\,
            sr => \N__46733\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_10_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26665\,
            in2 => \N__26264\,
            in3 => \N__26165\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_8\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_9\,
            clk => \N__47215\,
            ce => \N__26476\,
            sr => \N__46733\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_11_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26695\,
            in2 => \N__26638\,
            in3 => \N__26162\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_11\,
            ltout => OPEN,
            carryin => \bfn_9_22_0_\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_10\,
            clk => \N__47211\,
            ce => \N__26475\,
            sr => \N__46737\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_12_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26666\,
            in2 => \N__26608\,
            in3 => \N__26159\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_10\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_11\,
            clk => \N__47211\,
            ce => \N__26475\,
            sr => \N__46737\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_13_LC_9_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26581\,
            in2 => \N__26639\,
            in3 => \N__26210\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_11\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_12\,
            clk => \N__47211\,
            ce => \N__26475\,
            sr => \N__46737\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_14_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26560\,
            in2 => \N__26609\,
            in3 => \N__26207\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_12\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_13\,
            clk => \N__47211\,
            ce => \N__26475\,
            sr => \N__46737\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_15_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26582\,
            in2 => \N__26536\,
            in3 => \N__26204\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_13\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_14\,
            clk => \N__47211\,
            ce => \N__26475\,
            sr => \N__46737\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_16_LC_9_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26561\,
            in2 => \N__26509\,
            in3 => \N__26201\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_14\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_15\,
            clk => \N__47211\,
            ce => \N__26475\,
            sr => \N__46737\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_17_LC_9_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26914\,
            in2 => \N__26537\,
            in3 => \N__26198\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_15\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_16\,
            clk => \N__47211\,
            ce => \N__26475\,
            sr => \N__46737\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_18_LC_9_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26887\,
            in2 => \N__26510\,
            in3 => \N__26195\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_16\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_17\,
            clk => \N__47211\,
            ce => \N__26475\,
            sr => \N__46737\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_19_LC_9_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26915\,
            in2 => \N__26860\,
            in3 => \N__26192\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_19\,
            ltout => OPEN,
            carryin => \bfn_9_23_0_\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_18\,
            clk => \N__47208\,
            ce => \N__26474\,
            sr => \N__46738\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_20_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26888\,
            in2 => \N__26830\,
            in3 => \N__26189\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_18\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_19\,
            clk => \N__47208\,
            ce => \N__26474\,
            sr => \N__46738\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_21_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26800\,
            in2 => \N__26861\,
            in3 => \N__26186\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_19\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_20\,
            clk => \N__47208\,
            ce => \N__26474\,
            sr => \N__46738\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_22_LC_9_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26776\,
            in2 => \N__26831\,
            in3 => \N__26237\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_20\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_21\,
            clk => \N__47208\,
            ce => \N__26474\,
            sr => \N__46738\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_23_LC_9_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26801\,
            in2 => \N__26752\,
            in3 => \N__26234\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_21\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_22\,
            clk => \N__47208\,
            ce => \N__26474\,
            sr => \N__46738\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_24_LC_9_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26777\,
            in2 => \N__26722\,
            in3 => \N__26231\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_22\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_23\,
            clk => \N__47208\,
            ce => \N__26474\,
            sr => \N__46738\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_25_LC_9_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27070\,
            in2 => \N__26753\,
            in3 => \N__26228\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_23\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_24\,
            clk => \N__47208\,
            ce => \N__26474\,
            sr => \N__46738\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_26_LC_9_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27043\,
            in2 => \N__26723\,
            in3 => \N__26225\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_24\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_25\,
            clk => \N__47208\,
            ce => \N__26474\,
            sr => \N__46738\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_27_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27071\,
            in2 => \N__27016\,
            in3 => \N__26222\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_27\,
            ltout => OPEN,
            carryin => \bfn_9_24_0_\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_26\,
            clk => \N__47204\,
            ce => \N__26473\,
            sr => \N__46740\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_28_LC_9_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27044\,
            in2 => \N__26986\,
            in3 => \N__26219\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_26\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_27\,
            clk => \N__47204\,
            ce => \N__26473\,
            sr => \N__46740\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_29_LC_9_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26960\,
            in2 => \N__27017\,
            in3 => \N__26216\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_27\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_28\,
            clk => \N__47204\,
            ce => \N__26473\,
            sr => \N__46740\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_30_LC_9_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26936\,
            in2 => \N__26987\,
            in3 => \N__26213\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_28\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_29\,
            clk => \N__47204\,
            ce => \N__26473\,
            sr => \N__46740\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_31_LC_9_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26480\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47204\,
            ce => \N__26473\,
            sr => \N__46740\
        );

    \current_shift_inst.timer_phase.counter_0_LC_9_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32081\,
            in1 => \N__26442\,
            in2 => \_gnd_net_\,
            in3 => \N__26426\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_9_25_0_\,
            carryout => \current_shift_inst.timer_phase.counter_cry_0\,
            clk => \N__47199\,
            ce => \N__32134\,
            sr => \N__46741\
        );

    \current_shift_inst.timer_phase.counter_1_LC_9_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32077\,
            in1 => \N__26415\,
            in2 => \_gnd_net_\,
            in3 => \N__26402\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_0\,
            carryout => \current_shift_inst.timer_phase.counter_cry_1\,
            clk => \N__47199\,
            ce => \N__32134\,
            sr => \N__46741\
        );

    \current_shift_inst.timer_phase.counter_2_LC_9_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32082\,
            in1 => \N__26391\,
            in2 => \_gnd_net_\,
            in3 => \N__26375\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_1\,
            carryout => \current_shift_inst.timer_phase.counter_cry_2\,
            clk => \N__47199\,
            ce => \N__32134\,
            sr => \N__46741\
        );

    \current_shift_inst.timer_phase.counter_3_LC_9_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32078\,
            in1 => \N__26359\,
            in2 => \_gnd_net_\,
            in3 => \N__26345\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_2\,
            carryout => \current_shift_inst.timer_phase.counter_cry_3\,
            clk => \N__47199\,
            ce => \N__32134\,
            sr => \N__46741\
        );

    \current_shift_inst.timer_phase.counter_4_LC_9_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32083\,
            in1 => \N__26340\,
            in2 => \_gnd_net_\,
            in3 => \N__26324\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_3\,
            carryout => \current_shift_inst.timer_phase.counter_cry_4\,
            clk => \N__47199\,
            ce => \N__32134\,
            sr => \N__46741\
        );

    \current_shift_inst.timer_phase.counter_5_LC_9_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32079\,
            in1 => \N__26314\,
            in2 => \_gnd_net_\,
            in3 => \N__26300\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_4\,
            carryout => \current_shift_inst.timer_phase.counter_cry_5\,
            clk => \N__47199\,
            ce => \N__32134\,
            sr => \N__46741\
        );

    \current_shift_inst.timer_phase.counter_6_LC_9_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32084\,
            in1 => \N__26286\,
            in2 => \_gnd_net_\,
            in3 => \N__26267\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_5\,
            carryout => \current_shift_inst.timer_phase.counter_cry_6\,
            clk => \N__47199\,
            ce => \N__32134\,
            sr => \N__46741\
        );

    \current_shift_inst.timer_phase.counter_7_LC_9_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32080\,
            in1 => \N__26256\,
            in2 => \_gnd_net_\,
            in3 => \N__26240\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_6\,
            carryout => \current_shift_inst.timer_phase.counter_cry_7\,
            clk => \N__47199\,
            ce => \N__32134\,
            sr => \N__46741\
        );

    \current_shift_inst.timer_phase.counter_8_LC_9_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32064\,
            in1 => \N__26685\,
            in2 => \_gnd_net_\,
            in3 => \N__26669\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_9_26_0_\,
            carryout => \current_shift_inst.timer_phase.counter_cry_8\,
            clk => \N__47197\,
            ce => \N__32126\,
            sr => \N__46742\
        );

    \current_shift_inst.timer_phase.counter_9_LC_9_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32068\,
            in1 => \N__26658\,
            in2 => \_gnd_net_\,
            in3 => \N__26642\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_8\,
            carryout => \current_shift_inst.timer_phase.counter_cry_9\,
            clk => \N__47197\,
            ce => \N__32126\,
            sr => \N__46742\
        );

    \current_shift_inst.timer_phase.counter_10_LC_9_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32061\,
            in1 => \N__26626\,
            in2 => \_gnd_net_\,
            in3 => \N__26612\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_9\,
            carryout => \current_shift_inst.timer_phase.counter_cry_10\,
            clk => \N__47197\,
            ce => \N__32126\,
            sr => \N__46742\
        );

    \current_shift_inst.timer_phase.counter_11_LC_9_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32065\,
            in1 => \N__26601\,
            in2 => \_gnd_net_\,
            in3 => \N__26585\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_10\,
            carryout => \current_shift_inst.timer_phase.counter_cry_11\,
            clk => \N__47197\,
            ce => \N__32126\,
            sr => \N__46742\
        );

    \current_shift_inst.timer_phase.counter_12_LC_9_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32062\,
            in1 => \N__26580\,
            in2 => \_gnd_net_\,
            in3 => \N__26564\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_11\,
            carryout => \current_shift_inst.timer_phase.counter_cry_12\,
            clk => \N__47197\,
            ce => \N__32126\,
            sr => \N__46742\
        );

    \current_shift_inst.timer_phase.counter_13_LC_9_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32066\,
            in1 => \N__26554\,
            in2 => \_gnd_net_\,
            in3 => \N__26540\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_12\,
            carryout => \current_shift_inst.timer_phase.counter_cry_13\,
            clk => \N__47197\,
            ce => \N__32126\,
            sr => \N__46742\
        );

    \current_shift_inst.timer_phase.counter_14_LC_9_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32063\,
            in1 => \N__26529\,
            in2 => \_gnd_net_\,
            in3 => \N__26513\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_13\,
            carryout => \current_shift_inst.timer_phase.counter_cry_14\,
            clk => \N__47197\,
            ce => \N__32126\,
            sr => \N__46742\
        );

    \current_shift_inst.timer_phase.counter_15_LC_9_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32067\,
            in1 => \N__26497\,
            in2 => \_gnd_net_\,
            in3 => \N__26483\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_14\,
            carryout => \current_shift_inst.timer_phase.counter_cry_15\,
            clk => \N__47197\,
            ce => \N__32126\,
            sr => \N__46742\
        );

    \current_shift_inst.timer_phase.counter_16_LC_9_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32069\,
            in1 => \N__26907\,
            in2 => \_gnd_net_\,
            in3 => \N__26891\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_9_27_0_\,
            carryout => \current_shift_inst.timer_phase.counter_cry_16\,
            clk => \N__47195\,
            ce => \N__32135\,
            sr => \N__46744\
        );

    \current_shift_inst.timer_phase.counter_17_LC_9_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32073\,
            in1 => \N__26880\,
            in2 => \_gnd_net_\,
            in3 => \N__26864\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_16\,
            carryout => \current_shift_inst.timer_phase.counter_cry_17\,
            clk => \N__47195\,
            ce => \N__32135\,
            sr => \N__46744\
        );

    \current_shift_inst.timer_phase.counter_18_LC_9_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32070\,
            in1 => \N__26848\,
            in2 => \_gnd_net_\,
            in3 => \N__26834\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_17\,
            carryout => \current_shift_inst.timer_phase.counter_cry_18\,
            clk => \N__47195\,
            ce => \N__32135\,
            sr => \N__46744\
        );

    \current_shift_inst.timer_phase.counter_19_LC_9_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32074\,
            in1 => \N__26818\,
            in2 => \_gnd_net_\,
            in3 => \N__26804\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_18\,
            carryout => \current_shift_inst.timer_phase.counter_cry_19\,
            clk => \N__47195\,
            ce => \N__32135\,
            sr => \N__46744\
        );

    \current_shift_inst.timer_phase.counter_20_LC_9_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32071\,
            in1 => \N__26794\,
            in2 => \_gnd_net_\,
            in3 => \N__26780\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_19\,
            carryout => \current_shift_inst.timer_phase.counter_cry_20\,
            clk => \N__47195\,
            ce => \N__32135\,
            sr => \N__46744\
        );

    \current_shift_inst.timer_phase.counter_21_LC_9_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32075\,
            in1 => \N__26770\,
            in2 => \_gnd_net_\,
            in3 => \N__26756\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_20\,
            carryout => \current_shift_inst.timer_phase.counter_cry_21\,
            clk => \N__47195\,
            ce => \N__32135\,
            sr => \N__46744\
        );

    \current_shift_inst.timer_phase.counter_22_LC_9_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32072\,
            in1 => \N__26740\,
            in2 => \_gnd_net_\,
            in3 => \N__26726\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_21\,
            carryout => \current_shift_inst.timer_phase.counter_cry_22\,
            clk => \N__47195\,
            ce => \N__32135\,
            sr => \N__46744\
        );

    \current_shift_inst.timer_phase.counter_23_LC_9_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32076\,
            in1 => \N__26715\,
            in2 => \_gnd_net_\,
            in3 => \N__26699\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_22\,
            carryout => \current_shift_inst.timer_phase.counter_cry_23\,
            clk => \N__47195\,
            ce => \N__32135\,
            sr => \N__46744\
        );

    \current_shift_inst.timer_phase.counter_24_LC_9_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32085\,
            in1 => \N__27063\,
            in2 => \_gnd_net_\,
            in3 => \N__27047\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_9_28_0_\,
            carryout => \current_shift_inst.timer_phase.counter_cry_24\,
            clk => \N__47193\,
            ce => \N__32133\,
            sr => \N__46745\
        );

    \current_shift_inst.timer_phase.counter_25_LC_9_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32089\,
            in1 => \N__27036\,
            in2 => \_gnd_net_\,
            in3 => \N__27020\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_24\,
            carryout => \current_shift_inst.timer_phase.counter_cry_25\,
            clk => \N__47193\,
            ce => \N__32133\,
            sr => \N__46745\
        );

    \current_shift_inst.timer_phase.counter_26_LC_9_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32086\,
            in1 => \N__27004\,
            in2 => \_gnd_net_\,
            in3 => \N__26990\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_25\,
            carryout => \current_shift_inst.timer_phase.counter_cry_26\,
            clk => \N__47193\,
            ce => \N__32133\,
            sr => \N__46745\
        );

    \current_shift_inst.timer_phase.counter_27_LC_9_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32090\,
            in1 => \N__26979\,
            in2 => \_gnd_net_\,
            in3 => \N__26963\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_26\,
            carryout => \current_shift_inst.timer_phase.counter_cry_27\,
            clk => \N__47193\,
            ce => \N__32133\,
            sr => \N__46745\
        );

    \current_shift_inst.timer_phase.counter_28_LC_9_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32087\,
            in1 => \N__26956\,
            in2 => \_gnd_net_\,
            in3 => \N__26942\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_27\,
            carryout => \current_shift_inst.timer_phase.counter_cry_28\,
            clk => \N__47193\,
            ce => \N__32133\,
            sr => \N__46745\
        );

    \current_shift_inst.timer_phase.counter_29_LC_9_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__26935\,
            in1 => \N__32088\,
            in2 => \_gnd_net_\,
            in3 => \N__26939\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47193\,
            ce => \N__32133\,
            sr => \N__46745\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27397\,
            in2 => \_gnd_net_\,
            in3 => \N__40067\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MAX_D2_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26921\,
            lcout => \il_max_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47308\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNISQD2_0_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27153\,
            in2 => \_gnd_net_\,
            in3 => \N__27195\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlto2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIBO26_1_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__27112\,
            in1 => \N__27133\,
            in2 => \N__27209\,
            in3 => \N__27175\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlt9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIFA6C_5_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__27203\,
            in1 => \N__27347\,
            in2 => \N__27206\,
            in3 => \N__27092\,
            lcout => \pwm_generator_inst.un1_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIVDL3_9_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__27230\,
            in1 => \N__27305\,
            in2 => \_gnd_net_\,
            in3 => \N__27325\,
            lcout => \pwm_generator_inst.un1_counterlto9_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_0_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27276\,
            in1 => \N__27197\,
            in2 => \_gnd_net_\,
            in3 => \N__27179\,
            lcout => \pwm_generator_inst.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_10_9_0_\,
            carryout => \pwm_generator_inst.counter_cry_0\,
            clk => \N__47288\,
            ce => 'H',
            sr => \N__46638\
        );

    \pwm_generator_inst.counter_1_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27272\,
            in1 => \N__27176\,
            in2 => \_gnd_net_\,
            in3 => \N__27158\,
            lcout => \pwm_generator_inst.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_0\,
            carryout => \pwm_generator_inst.counter_cry_1\,
            clk => \N__47288\,
            ce => 'H',
            sr => \N__46638\
        );

    \pwm_generator_inst.counter_2_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27277\,
            in1 => \N__27155\,
            in2 => \_gnd_net_\,
            in3 => \N__27137\,
            lcout => \pwm_generator_inst.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_1\,
            carryout => \pwm_generator_inst.counter_cry_2\,
            clk => \N__47288\,
            ce => 'H',
            sr => \N__46638\
        );

    \pwm_generator_inst.counter_3_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27273\,
            in1 => \N__27134\,
            in2 => \_gnd_net_\,
            in3 => \N__27116\,
            lcout => \pwm_generator_inst.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_2\,
            carryout => \pwm_generator_inst.counter_cry_3\,
            clk => \N__47288\,
            ce => 'H',
            sr => \N__46638\
        );

    \pwm_generator_inst.counter_4_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27278\,
            in1 => \N__27113\,
            in2 => \_gnd_net_\,
            in3 => \N__27095\,
            lcout => \pwm_generator_inst.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_3\,
            carryout => \pwm_generator_inst.counter_cry_4\,
            clk => \N__47288\,
            ce => 'H',
            sr => \N__46638\
        );

    \pwm_generator_inst.counter_5_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27274\,
            in1 => \N__27091\,
            in2 => \_gnd_net_\,
            in3 => \N__27074\,
            lcout => \pwm_generator_inst.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_4\,
            carryout => \pwm_generator_inst.counter_cry_5\,
            clk => \N__47288\,
            ce => 'H',
            sr => \N__46638\
        );

    \pwm_generator_inst.counter_6_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27279\,
            in1 => \N__27346\,
            in2 => \_gnd_net_\,
            in3 => \N__27329\,
            lcout => \pwm_generator_inst.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_5\,
            carryout => \pwm_generator_inst.counter_cry_6\,
            clk => \N__47288\,
            ce => 'H',
            sr => \N__46638\
        );

    \pwm_generator_inst.counter_7_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27275\,
            in1 => \N__27326\,
            in2 => \_gnd_net_\,
            in3 => \N__27308\,
            lcout => \pwm_generator_inst.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_6\,
            carryout => \pwm_generator_inst.counter_cry_7\,
            clk => \N__47288\,
            ce => 'H',
            sr => \N__46638\
        );

    \pwm_generator_inst.counter_8_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27281\,
            in1 => \N__27304\,
            in2 => \_gnd_net_\,
            in3 => \N__27284\,
            lcout => \pwm_generator_inst.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_10_10_0_\,
            carryout => \pwm_generator_inst.counter_cry_8\,
            clk => \N__47281\,
            ce => 'H',
            sr => \N__46645\
        );

    \pwm_generator_inst.counter_9_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27280\,
            in1 => \N__27229\,
            in2 => \_gnd_net_\,
            in3 => \N__27233\,
            lcout => \pwm_generator_inst.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47281\,
            ce => 'H',
            sr => \N__46645\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__39662\,
            in1 => \N__39978\,
            in2 => \N__39848\,
            in3 => \N__28895\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47281\,
            ce => 'H',
            sr => \N__46645\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__39820\,
            in1 => \N__39667\,
            in2 => \N__40014\,
            in3 => \N__29207\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47281\,
            ce => 'H',
            sr => \N__46645\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__39663\,
            in1 => \N__39988\,
            in2 => \N__39849\,
            in3 => \N__29180\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47281\,
            ce => 'H',
            sr => \N__46645\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__39819\,
            in1 => \N__39666\,
            in2 => \N__40013\,
            in3 => \N__29264\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47281\,
            ce => 'H',
            sr => \N__46645\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__39664\,
            in1 => \N__39989\,
            in2 => \N__39850\,
            in3 => \N__29096\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47281\,
            ce => 'H',
            sr => \N__46645\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__39818\,
            in1 => \N__39665\,
            in2 => \N__40012\,
            in3 => \N__28865\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47281\,
            ce => 'H',
            sr => \N__46645\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100010001100"
        )
    port map (
            in0 => \N__39811\,
            in1 => \N__29126\,
            in2 => \N__39680\,
            in3 => \N__39932\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47272\,
            ce => 'H',
            sr => \N__46653\
        );

    \phase_controller_inst1.stoper_hc.time_passed_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__31106\,
            in1 => \N__27398\,
            in2 => \N__27368\,
            in3 => \N__40064\,
            lcout => \phase_controller_inst1.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47272\,
            ce => 'H',
            sr => \N__46653\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010000100"
        )
    port map (
            in0 => \N__39669\,
            in1 => \N__29153\,
            in2 => \N__39977\,
            in3 => \N__39812\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47272\,
            ce => 'H',
            sr => \N__46653\
        );

    \phase_controller_inst1.stoper_hc.target_time_14_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__43899\,
            in1 => \N__44087\,
            in2 => \_gnd_net_\,
            in3 => \N__33878\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47262\,
            ce => \N__31225\,
            sr => \N__46663\
        );

    \phase_controller_inst1.stoper_hc.target_time_11_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__44086\,
            in1 => \N__39352\,
            in2 => \_gnd_net_\,
            in3 => \N__43898\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47262\,
            ce => \N__31225\,
            sr => \N__46663\
        );

    \phase_controller_inst1.stoper_hc.target_time_9_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010000000101"
        )
    port map (
            in0 => \N__40344\,
            in1 => \N__34048\,
            in2 => \N__44155\,
            in3 => \N__43900\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47262\,
            ce => \N__31225\,
            sr => \N__46663\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39608\,
            in2 => \_gnd_net_\,
            in3 => \N__39766\,
            lcout => \phase_controller_inst1.stoper_hc.time_passed11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__39961\,
            in1 => \N__39609\,
            in2 => \_gnd_net_\,
            in3 => \N__39767\,
            lcout => \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_0_c_inv_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29293\,
            in2 => \N__27356\,
            in3 => \N__29325\,
            lcout => \G_407\,
            ltout => OPEN,
            carryin => \bfn_10_14_0_\,
            carryout => \current_shift_inst.z_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_1_c_inv_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27443\,
            in2 => \N__29604\,
            in3 => \N__27599\,
            lcout => \G_406\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_0\,
            carryout => \current_shift_inst.z_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_2_c_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29569\,
            in2 => \N__27545\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_1\,
            carryout => \current_shift_inst.z_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_3_c_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29548\,
            in2 => \N__27506\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_2\,
            carryout => \current_shift_inst.z_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_4_c_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27458\,
            in2 => \N__29519\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_3\,
            carryout => \current_shift_inst.z_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_5_c_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29472\,
            in2 => \N__27821\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_4\,
            carryout => \current_shift_inst.z_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_6_c_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27773\,
            in2 => \N__29442\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_5\,
            carryout => \current_shift_inst.z_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_7_c_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27722\,
            in2 => \N__29391\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_6\,
            carryout => \current_shift_inst.z_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_8_c_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27707\,
            in2 => \N__29837\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_15_0_\,
            carryout => \current_shift_inst.z_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_9_c_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27692\,
            in2 => \N__30029\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_8\,
            carryout => \current_shift_inst.z_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_10_c_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29721\,
            in2 => \N__27650\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_9\,
            carryout => \current_shift_inst.z_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_11_c_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27632\,
            in2 => \N__30707\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_10\,
            carryout => \current_shift_inst.z_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_12_c_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27617\,
            in2 => \N__30737\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_11\,
            carryout => \current_shift_inst.z_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_13_c_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28064\,
            in2 => \N__29921\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_12\,
            carryout => \current_shift_inst.z_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_14_c_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28049\,
            in2 => \N__30197\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_13\,
            carryout => \current_shift_inst.z_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_15_c_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28034\,
            in2 => \N__30233\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_14\,
            carryout => \current_shift_inst.z_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_16_c_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30303\,
            in2 => \N__28019\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_16_0_\,
            carryout => \current_shift_inst.z_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_17_c_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27968\,
            in2 => \N__29670\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_16\,
            carryout => \current_shift_inst.z_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_18_c_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29631\,
            in2 => \N__27920\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_17\,
            carryout => \current_shift_inst.z_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_19_c_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27902\,
            in2 => \N__30416\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_18\,
            carryout => \current_shift_inst.z_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_20_c_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27887\,
            in2 => \N__31070\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_19\,
            carryout => \current_shift_inst.z_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_21_c_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30954\,
            in2 => \N__27872\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_20\,
            carryout => \current_shift_inst.z_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_22_c_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28226\,
            in2 => \N__29770\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_21\,
            carryout => \current_shift_inst.z_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_23_c_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31572\,
            in2 => \N__28211\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_22\,
            carryout => \current_shift_inst.z_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_24_c_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28193\,
            in2 => \N__31507\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_17_0_\,
            carryout => \current_shift_inst.z_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_25_c_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31748\,
            in2 => \N__28178\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_24\,
            carryout => \current_shift_inst.z_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_26_c_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28160\,
            in2 => \N__31824\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_25\,
            carryout => \current_shift_inst.z_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_27_c_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28112\,
            in2 => \N__30111\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_26\,
            carryout => \current_shift_inst.z_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_28_c_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28097\,
            in2 => \N__30831\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_27\,
            carryout => \current_shift_inst.z_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_29_c_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31671\,
            in2 => \N__28082\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_28\,
            carryout => \current_shift_inst.z_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_30_c_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30489\,
            in2 => \N__28469\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_29\,
            carryout => \current_shift_inst.z_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_s_31_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__30574\,
            in1 => \N__28448\,
            in2 => \N__30529\,
            in3 => \N__27602\,
            lcout => \current_shift_inst.z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_1_c_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27591\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_18_0_\,
            carryout => \current_shift_inst.z_5_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_2_s_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27563\,
            in2 => \N__28693\,
            in3 => \N__27530\,
            lcout => \current_shift_inst.z_5_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_1\,
            carryout => \current_shift_inst.z_5_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_3_s_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27520\,
            in2 => \N__28697\,
            in3 => \N__27491\,
            lcout => \current_shift_inst.z_5_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_2\,
            carryout => \current_shift_inst.z_5_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_4_s_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27485\,
            in2 => \N__28694\,
            in3 => \N__27446\,
            lcout => \current_shift_inst.z_5_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_3\,
            carryout => \current_shift_inst.z_5_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_5_s_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27842\,
            in2 => \N__28698\,
            in3 => \N__27806\,
            lcout => \current_shift_inst.z_5_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_4\,
            carryout => \current_shift_inst.z_5_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_6_s_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27797\,
            in2 => \N__28695\,
            in3 => \N__27761\,
            lcout => \current_shift_inst.z_5_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_5\,
            carryout => \current_shift_inst.z_5_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_7_s_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27757\,
            in2 => \N__28699\,
            in3 => \N__27710\,
            lcout => \current_shift_inst.z_5_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_6\,
            carryout => \current_shift_inst.z_5_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_8_s_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29873\,
            in2 => \N__28696\,
            in3 => \N__27695\,
            lcout => \current_shift_inst.z_5_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_7\,
            carryout => \current_shift_inst.z_5_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_9_s_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30065\,
            in2 => \N__28847\,
            in3 => \N__27680\,
            lcout => \current_shift_inst.z_5_9\,
            ltout => OPEN,
            carryin => \bfn_10_19_0_\,
            carryout => \current_shift_inst.z_5_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_10_s_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27674\,
            in2 => \N__28841\,
            in3 => \N__27635\,
            lcout => \current_shift_inst.z_5_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_9\,
            carryout => \current_shift_inst.z_5_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_11_s_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30762\,
            in2 => \N__28844\,
            in3 => \N__27620\,
            lcout => \current_shift_inst.z_5_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_10\,
            carryout => \current_shift_inst.z_5_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_12_s_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30663\,
            in2 => \N__28842\,
            in3 => \N__27605\,
            lcout => \current_shift_inst.z_5_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_11\,
            carryout => \current_shift_inst.z_5_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_13_s_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29957\,
            in2 => \N__28845\,
            in3 => \N__28052\,
            lcout => \current_shift_inst.z_5_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_12\,
            carryout => \current_shift_inst.z_5_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_14_s_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30269\,
            in2 => \N__28843\,
            in3 => \N__28037\,
            lcout => \current_shift_inst.z_5_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_13\,
            carryout => \current_shift_inst.z_5_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_15_s_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30164\,
            in2 => \N__28846\,
            in3 => \N__28022\,
            lcout => \current_shift_inst.z_5_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_14\,
            carryout => \current_shift_inst.z_5_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_16_s_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28792\,
            in2 => \N__30357\,
            in3 => \N__28004\,
            lcout => \current_shift_inst.z_5_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_15\,
            carryout => \current_shift_inst.z_5_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_17_s_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27992\,
            in2 => \N__28833\,
            in3 => \N__27956\,
            lcout => \current_shift_inst.z_5_17\,
            ltout => OPEN,
            carryin => \bfn_10_20_0_\,
            carryout => \current_shift_inst.z_5_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_18_s_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27939\,
            in2 => \N__28837\,
            in3 => \N__27905\,
            lcout => \current_shift_inst.z_5_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_17\,
            carryout => \current_shift_inst.z_5_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_19_s_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30452\,
            in2 => \N__28834\,
            in3 => \N__27890\,
            lcout => \current_shift_inst.z_5_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_18\,
            carryout => \current_shift_inst.z_5_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_20_s_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31033\,
            in2 => \N__28838\,
            in3 => \N__27875\,
            lcout => \current_shift_inst.z_5_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_19\,
            carryout => \current_shift_inst.z_5_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_21_s_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30992\,
            in2 => \N__28835\,
            in3 => \N__28253\,
            lcout => \current_shift_inst.z_5_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_20\,
            carryout => \current_shift_inst.z_5_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_22_s_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28247\,
            in2 => \N__28839\,
            in3 => \N__28214\,
            lcout => \current_shift_inst.z_5_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_21\,
            carryout => \current_shift_inst.z_5_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_23_s_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31548\,
            in2 => \N__28836\,
            in3 => \N__28196\,
            lcout => \current_shift_inst.z_5_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_22\,
            carryout => \current_shift_inst.z_5_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_24_s_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31622\,
            in2 => \N__28840\,
            in3 => \N__28181\,
            lcout => \current_shift_inst.z_5_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_23\,
            carryout => \current_shift_inst.z_5_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_25_s_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31768\,
            in2 => \N__28827\,
            in3 => \N__28163\,
            lcout => \current_shift_inst.z_5_25\,
            ltout => OPEN,
            carryin => \bfn_10_21_0_\,
            carryout => \current_shift_inst.z_5_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_26_s_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31859\,
            in2 => \N__28830\,
            in3 => \N__28148\,
            lcout => \current_shift_inst.z_5_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_25\,
            carryout => \current_shift_inst.z_5_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_27_s_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28139\,
            in2 => \N__28828\,
            in3 => \N__28100\,
            lcout => \current_shift_inst.z_5_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_26\,
            carryout => \current_shift_inst.z_5_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_28_s_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30869\,
            in2 => \N__28831\,
            in3 => \N__28085\,
            lcout => \current_shift_inst.z_5_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_27\,
            carryout => \current_shift_inst.z_5_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_29_s_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31704\,
            in2 => \N__28829\,
            in3 => \N__28067\,
            lcout => \current_shift_inst.z_5_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_28\,
            carryout => \current_shift_inst.z_5_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_30_s_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30630\,
            in2 => \N__28832\,
            in3 => \N__28454\,
            lcout => \current_shift_inst.z_5_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_29\,
            carryout => \current_shift_inst.z_5_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.z_5_cry_30_THRU_LUT4_0_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28451\,
            lcout => \current_shift_inst.z_5_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.S2_LC_10_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32255\,
            lcout => s4_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47190\,
            ce => 'H',
            sr => \N__46743\
        );

    \SB_DFF_inst_PH1_MIN_D1_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28421\,
            lcout => \il_min_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47309\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28406\,
            in2 => \N__28391\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_8_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28361\,
            in2 => \_gnd_net_\,
            in3 => \N__28331\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28328\,
            in2 => \N__28322\,
            in3 => \N__28289\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28286\,
            in2 => \_gnd_net_\,
            in3 => \N__28256\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29081\,
            in2 => \_gnd_net_\,
            in3 => \N__29051\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29048\,
            in2 => \_gnd_net_\,
            in3 => \N__29018\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29015\,
            in2 => \_gnd_net_\,
            in3 => \N__28985\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28982\,
            in2 => \_gnd_net_\,
            in3 => \N__28952\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31138\,
            in2 => \_gnd_net_\,
            in3 => \N__28949\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_11_9_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28946\,
            in2 => \_gnd_net_\,
            in3 => \N__28919\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28915\,
            in3 => \N__28889\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28885\,
            in3 => \N__28859\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29278\,
            in2 => \_gnd_net_\,
            in3 => \N__29258\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29255\,
            in2 => \_gnd_net_\,
            in3 => \N__29228\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29221\,
            in2 => \_gnd_net_\,
            in3 => \N__29201\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29194\,
            in2 => \_gnd_net_\,
            in3 => \N__29174\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29167\,
            in2 => \_gnd_net_\,
            in3 => \N__29147\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \bfn_11_10_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29140\,
            in2 => \_gnd_net_\,
            in3 => \N__29120\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29113\,
            in2 => \_gnd_net_\,
            in3 => \N__29099\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MIN_D2_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29090\,
            lcout => \il_min_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47273\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_6_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__34150\,
            in1 => \N__34047\,
            in2 => \_gnd_net_\,
            in3 => \N__35431\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_10_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001110000"
        )
    port map (
            in0 => \N__35513\,
            in1 => \N__34107\,
            in2 => \N__29357\,
            in3 => \N__41253\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_15_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__44084\,
            in1 => \N__33916\,
            in2 => \_gnd_net_\,
            in3 => \N__43878\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47253\,
            ce => \N__31229\,
            sr => \N__46654\
        );

    \phase_controller_inst1.stoper_hc.target_time_18_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__43879\,
            in1 => \N__44085\,
            in2 => \_gnd_net_\,
            in3 => \N__42191\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47253\,
            ce => \N__31229\,
            sr => \N__46654\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35854\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47245\,
            ce => \N__32738\,
            sr => \N__46664\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35827\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47245\,
            ce => \N__32738\,
            sr => \N__46664\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32716\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47245\,
            ce => \N__32738\,
            sr => \N__46664\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32717\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_1_fast_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47245\,
            ce => \N__32738\,
            sr => \N__46664\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_RNI48NB_31_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31328\,
            in2 => \N__29327\,
            in3 => \N__29326\,
            lcout => \current_shift_inst.un38_control_input_0\,
            ltout => OPEN,
            carryin => \bfn_11_14_0_\,
            carryout => \current_shift_inst.un4_control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_1_c_RNIJF2G_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31316\,
            in2 => \_gnd_net_\,
            in3 => \N__29585\,
            lcout => \current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_1\,
            carryout => \current_shift_inst.un4_control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_2_c_RNILI3G_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31163\,
            in3 => \N__29558\,
            lcout => \current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_2\,
            carryout => \current_shift_inst.un4_control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_3_c_RNINL4G_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31154\,
            in2 => \_gnd_net_\,
            in3 => \N__29537\,
            lcout => \current_shift_inst.un4_control_input_cry_3_c_RNINL4GZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_3\,
            carryout => \current_shift_inst.un4_control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_4_c_RNIPO5G_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31298\,
            in2 => \_gnd_net_\,
            in3 => \N__29492\,
            lcout => \current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_4\,
            carryout => \current_shift_inst.un4_control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_5_c_RNIRR6G_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31289\,
            in3 => \N__29456\,
            lcout => \current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_5\,
            carryout => \current_shift_inst.un4_control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_6_c_RNITU7G_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31277\,
            in2 => \_gnd_net_\,
            in3 => \N__29417\,
            lcout => \current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_6\,
            carryout => \current_shift_inst.un4_control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_7_c_RNIV19G_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33749\,
            in2 => \_gnd_net_\,
            in3 => \N__29366\,
            lcout => \current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_7\,
            carryout => \current_shift_inst.un4_control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_8_c_RNI15AG_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33980\,
            in2 => \_gnd_net_\,
            in3 => \N__29363\,
            lcout => \current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0\,
            ltout => OPEN,
            carryin => \bfn_11_15_0_\,
            carryout => \current_shift_inst.un4_control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_9_c_RNIALDJ_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31376\,
            in2 => \_gnd_net_\,
            in3 => \N__29360\,
            lcout => \current_shift_inst.un4_control_input_cry_9_c_RNIALDJZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_9\,
            carryout => \current_shift_inst.un4_control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_10_c_RNIJLTG_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31391\,
            in2 => \_gnd_net_\,
            in3 => \N__29705\,
            lcout => \current_shift_inst.un4_control_input_cry_10_c_RNIJLTGZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_10\,
            carryout => \current_shift_inst.un4_control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_11_c_RNILOUG_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31370\,
            in2 => \_gnd_net_\,
            in3 => \N__29702\,
            lcout => \current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_11\,
            carryout => \current_shift_inst.un4_control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_12_c_RNINRVG_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33926\,
            in2 => \_gnd_net_\,
            in3 => \N__29699\,
            lcout => \current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_12\,
            carryout => \current_shift_inst.un4_control_input_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_13_c_RNIPU0H_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31364\,
            in2 => \_gnd_net_\,
            in3 => \N__29696\,
            lcout => \current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_13\,
            carryout => \current_shift_inst.un4_control_input_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_14_c_RNIR12H_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31304\,
            in2 => \_gnd_net_\,
            in3 => \N__29693\,
            lcout => \current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_14\,
            carryout => \current_shift_inst.un4_control_input_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_15_c_RNIT43H_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33962\,
            in2 => \_gnd_net_\,
            in3 => \N__29690\,
            lcout => \current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_15\,
            carryout => \current_shift_inst.un4_control_input_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_16_c_RNIV74H_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33944\,
            in2 => \_gnd_net_\,
            in3 => \N__29687\,
            lcout => \current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0\,
            ltout => OPEN,
            carryin => \bfn_11_16_0_\,
            carryout => \current_shift_inst.un4_control_input_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_17_c_RNI1B5H_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31358\,
            in2 => \_gnd_net_\,
            in3 => \N__29648\,
            lcout => \current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_17\,
            carryout => \current_shift_inst.un4_control_input_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_18_c_RNI3E6H_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31385\,
            in3 => \N__29795\,
            lcout => \current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_18\,
            carryout => \current_shift_inst.un4_control_input_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_19_c_RNIS88H_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31442\,
            in2 => \_gnd_net_\,
            in3 => \N__29792\,
            lcout => \current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_19\,
            carryout => \current_shift_inst.un4_control_input_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_20_c_RNILQ1I_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31454\,
            in2 => \_gnd_net_\,
            in3 => \N__29789\,
            lcout => \current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_20\,
            carryout => \current_shift_inst.un4_control_input_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_21_c_RNINT2I_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31346\,
            in2 => \_gnd_net_\,
            in3 => \N__29786\,
            lcout => \current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_21\,
            carryout => \current_shift_inst.un4_control_input_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_22_c_RNIP04I_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33734\,
            in2 => \_gnd_net_\,
            in3 => \N__29753\,
            lcout => \current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_22\,
            carryout => \current_shift_inst.un4_control_input_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_23_c_RNIR35I_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31310\,
            in2 => \_gnd_net_\,
            in3 => \N__29750\,
            lcout => \current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_23\,
            carryout => \current_shift_inst.un4_control_input_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_24_c_RNIT66I_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31448\,
            in2 => \_gnd_net_\,
            in3 => \N__29747\,
            lcout => \current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0\,
            ltout => OPEN,
            carryin => \bfn_11_17_0_\,
            carryout => \current_shift_inst.un4_control_input_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_25_c_RNIV97I_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31340\,
            in2 => \_gnd_net_\,
            in3 => \N__29744\,
            lcout => \current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_25\,
            carryout => \current_shift_inst.un4_control_input_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_26_c_RNI1D8I_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31466\,
            in2 => \_gnd_net_\,
            in3 => \N__29741\,
            lcout => \current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_26\,
            carryout => \current_shift_inst.un4_control_input_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_27_c_RNI3G9I_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31397\,
            in2 => \_gnd_net_\,
            in3 => \N__30086\,
            lcout => \current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_27\,
            carryout => \current_shift_inst.un4_control_input_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_28_c_RNI5JAI_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31352\,
            in2 => \_gnd_net_\,
            in3 => \N__30083\,
            lcout => \current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_28\,
            carryout => \current_shift_inst.un4_control_input_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_29_c_RNIUDCI_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31460\,
            in2 => \_gnd_net_\,
            in3 => \N__30080\,
            lcout => \current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_29\,
            carryout => \current_shift_inst.un4_control_input_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_30_c_RNINV5J_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30560\,
            in2 => \_gnd_net_\,
            in3 => \N__30077\,
            lcout => \current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIO0U12_8_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__29882\,
            in1 => \N__30073\,
            in2 => \N__29845\,
            in3 => \N__30030\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIO0U12_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILORI_11_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__30771\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30708\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNILORI_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOSSI_12_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__30739\,
            in1 => \_gnd_net_\,
            in2 => \N__30679\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIOSSI_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJTQ51_12_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__29967\,
            in1 => \N__30740\,
            in2 => \N__30680\,
            in3 => \N__29925\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJTQ51_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIN7DV_8_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29881\,
            in2 => \_gnd_net_\,
            in3 => \N__29838\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIN7DV_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDS8K_28_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30884\,
            in2 => \_gnd_net_\,
            in3 => \N__30827\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIDS8K_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5S981_24_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__31628\,
            in1 => \N__31749\,
            in2 => \N__31508\,
            in3 => \N__31784\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5S981_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDLO51_11_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__30772\,
            in1 => \N__30738\,
            in2 => \N__30716\,
            in3 => \N__30672\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIDLO51_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_RNO_0_25_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110010110"
        )
    port map (
            in0 => \N__30638\,
            in1 => \N__30590\,
            in2 => \N__30533\,
            in3 => \N__30499\,
            lcout => \current_shift_inst.un38_control_input_0_axb_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPC571_19_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__30464\,
            in1 => \N__31041\,
            in2 => \N__30425\,
            in3 => \N__31071\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPC571_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI190J_15_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30166\,
            in2 => \_gnd_net_\,
            in3 => \N__30234\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI190J_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5M161_15_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__30167\,
            in1 => \N__30359\,
            in2 => \N__30239\,
            in3 => \N__30312\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5M161_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVDV51_14_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__30278\,
            in1 => \N__30235\,
            in2 => \N__30212\,
            in3 => \N__30165\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIVDV51_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDR081_20_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__31003\,
            in1 => \N__31045\,
            in2 => \N__31076\,
            in3 => \N__30963\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIDR081_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILRVJ_20_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__31072\,
            in1 => \_gnd_net_\,
            in2 => \N__31046\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNILRVJ_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOV0K_21_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31002\,
            in2 => \_gnd_net_\,
            in3 => \N__30964\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIOV0K_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU73K_23_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31549\,
            in2 => \_gnd_net_\,
            in3 => \N__31592\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIU73K_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.start_timer_tr_RNO_1_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32250\,
            in2 => \_gnd_net_\,
            in3 => \N__32217\,
            lcout => \phase_controller_slave.start_timer_tr_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7K6K_26_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31867\,
            in2 => \_gnd_net_\,
            in3 => \N__31825\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI7K6K_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MAX_D2_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30899\,
            lcout => \il_max_comp2_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47205\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.state_1_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__32218\,
            in1 => \N__47637\,
            in2 => \N__32251\,
            in3 => \N__47665\,
            lcout => \phase_controller_slave.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47201\,
            ce => 'H',
            sr => \N__46725\
        );

    \delay_measurement_inst.delay_hc_reg_6_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011111111"
        )
    port map (
            in0 => \N__35129\,
            in1 => \N__42648\,
            in2 => \N__34158\,
            in3 => \N__42102\,
            lcout => measured_delay_hc_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47271\,
            ce => 'H',
            sr => \N__46627\
        );

    \phase_controller_inst1.state_1_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__43076\,
            in1 => \N__31115\,
            in2 => \N__33787\,
            in3 => \N__43023\,
            lcout => \phase_controller_inst1.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47261\,
            ce => 'H',
            sr => \N__46633\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__39668\,
            in1 => \N__39768\,
            in2 => \N__39928\,
            in3 => \N__31148\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47261\,
            ce => 'H',
            sr => \N__46633\
        );

    \phase_controller_inst1.start_timer_hc_RNO_1_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32504\,
            in2 => \_gnd_net_\,
            in3 => \N__32538\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.start_timer_hc_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__43153\,
            in1 => \N__39910\,
            in2 => \N__31124\,
            in3 => \N__31121\,
            lcout => \phase_controller_inst1.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47252\,
            ce => 'H',
            sr => \N__46639\
        );

    \phase_controller_inst1.start_timer_hc_RNO_0_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33773\,
            in2 => \_gnd_net_\,
            in3 => \N__31110\,
            lcout => \phase_controller_inst1.N_88\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_2_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__31111\,
            in1 => \N__32505\,
            in2 => \N__33783\,
            in3 => \N__32539\,
            lcout => \phase_controller_inst1.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47252\,
            ce => 'H',
            sr => \N__46639\
        );

    \phase_controller_slave.stoper_tr.target_time_10_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__47598\,
            in1 => \N__39473\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47244\,
            ce => \N__44417\,
            sr => \N__46646\
        );

    \phase_controller_slave.stoper_tr.target_time_11_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47595\,
            in2 => \_gnd_net_\,
            in3 => \N__41531\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47244\,
            ce => \N__44417\,
            sr => \N__46646\
        );

    \phase_controller_slave.stoper_tr.target_time_12_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47596\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39500\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47244\,
            ce => \N__44417\,
            sr => \N__46646\
        );

    \phase_controller_slave.stoper_tr.target_time_13_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__41999\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47597\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47244\,
            ce => \N__44417\,
            sr => \N__46646\
        );

    \phase_controller_slave.stoper_tr.target_time_15_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41489\,
            in2 => \_gnd_net_\,
            in3 => \N__47520\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47244\,
            ce => \N__44417\,
            sr => \N__46646\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32471\,
            lcout => \current_shift_inst.un4_control_input_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32462\,
            lcout => \current_shift_inst.un4_control_input_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32453\,
            lcout => \current_shift_inst.un4_control_input_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_16_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__44061\,
            in1 => \N__40453\,
            in2 => \_gnd_net_\,
            in3 => \N__43887\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47237\,
            ce => \N__31228\,
            sr => \N__46655\
        );

    \phase_controller_inst1.stoper_hc.target_time_17_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__43888\,
            in1 => \N__44062\,
            in2 => \_gnd_net_\,
            in3 => \N__42346\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47237\,
            ce => \N__31228\,
            sr => \N__46655\
        );

    \phase_controller_inst1.stoper_hc.target_time_19_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100110011"
        )
    port map (
            in0 => \N__41887\,
            in1 => \N__44060\,
            in2 => \_gnd_net_\,
            in3 => \N__40389\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47237\,
            ce => \N__31228\,
            sr => \N__46655\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32486\,
            lcout => \current_shift_inst.un4_control_input_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32480\,
            lcout => \current_shift_inst.un4_control_input_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.stoper_state_1_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000001100100"
        )
    port map (
            in0 => \N__40981\,
            in1 => \N__40655\,
            in2 => \N__40916\,
            in3 => \N__40739\,
            lcout => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47229\,
            ce => \N__40514\,
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.stoper_state_0_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__37793\,
            in1 => \N__38103\,
            in2 => \N__38051\,
            in3 => \N__34417\,
            lcout => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47229\,
            ce => \N__40514\,
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.stoper_state_1_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001010000"
        )
    port map (
            in0 => \N__34418\,
            in1 => \N__38039\,
            in2 => \N__38144\,
            in3 => \N__37794\,
            lcout => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47229\,
            ce => \N__40514\,
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.tr_state_0_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001100110"
        )
    port map (
            in0 => \N__34910\,
            in1 => \N__33826\,
            in2 => \_gnd_net_\,
            in3 => \N__33812\,
            lcout => \delay_measurement_inst.tr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47229\,
            ce => \N__40514\,
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.hc_state_0_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__35881\,
            in1 => \N__35916\,
            in2 => \_gnd_net_\,
            in3 => \N__41939\,
            lcout => \delay_measurement_inst.hc_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47229\,
            ce => \N__40514\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31334\,
            lcout => \current_shift_inst.un4_control_input_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31322\,
            lcout => \current_shift_inst.un4_control_input_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32621\,
            lcout => \current_shift_inst.un4_control_input_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32555\,
            lcout => \current_shift_inst.un4_control_input_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32585\,
            lcout => \current_shift_inst.un4_control_input_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32660\,
            lcout => \current_shift_inst.un4_control_input_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32597\,
            lcout => \current_shift_inst.un4_control_input_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32576\,
            lcout => \current_shift_inst.un4_control_input_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32564\,
            lcout => \current_shift_inst.un4_control_input_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32669\,
            lcout => \current_shift_inst.un4_control_input_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32759\,
            lcout => \current_shift_inst.un4_control_input_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32633\,
            lcout => \current_shift_inst.un4_control_input_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32786\,
            lcout => \current_shift_inst.un4_control_input_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32777\,
            lcout => \current_shift_inst.un4_control_input_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32750\,
            lcout => \current_shift_inst.un4_control_input_axb_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32642\,
            lcout => \current_shift_inst.un4_control_input_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32612\,
            lcout => \current_shift_inst.un4_control_input_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32651\,
            lcout => \current_shift_inst.un4_control_input_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__32426\,
            in1 => \N__40393\,
            in2 => \_gnd_net_\,
            in3 => \N__41886\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlt31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_i_31_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31436\,
            lcout => \current_shift_inst.z_i_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32768\,
            lcout => \current_shift_inst.un4_control_input_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_ibuf_gb_io_RNI79U7_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46777\,
            lcout => red_c_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1C4K_24_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__31502\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31627\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI1C4K_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIB4C81_25_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \N__31751\,
            in1 => \N__31783\,
            in2 => \N__31871\,
            in3 => \N__31823\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIB4C81_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4G5K_25_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__31782\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31750\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI4G5K_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7OAK_29_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31712\,
            in2 => \_gnd_net_\,
            in3 => \N__31675\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI7OAK_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVJ781_23_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__31626\,
            in1 => \N__31587\,
            in2 => \N__31556\,
            in3 => \N__31503\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIVJ781_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.S3_sync0_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31903\,
            lcout => \current_shift_inst.S3_syncZ0Z0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47212\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__47443\,
            in1 => \N__34223\,
            in2 => \N__31931\,
            in3 => \N__47401\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.target_time_2_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000110000000000"
        )
    port map (
            in0 => \N__40217\,
            in1 => \N__40094\,
            in2 => \N__31469\,
            in3 => \N__37465\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47209\,
            ce => \N__44449\,
            sr => \N__46707\
        );

    \phase_controller_slave.stoper_tr.target_time_3_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__37466\,
            in1 => \N__40216\,
            in2 => \_gnd_net_\,
            in3 => \N__37422\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47209\,
            ce => \N__44449\,
            sr => \N__46707\
        );

    \phase_controller_slave.stoper_tr.target_time_1_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__37423\,
            in1 => \N__37046\,
            in2 => \N__40121\,
            in3 => \N__37464\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47209\,
            ce => \N__44449\,
            sr => \N__46707\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1_6_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__37224\,
            in1 => \N__37326\,
            in2 => \_gnd_net_\,
            in3 => \N__40248\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1Z0Z_6\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0_6_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47537\,
            in2 => \N__31922\,
            in3 => \N__47400\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.target_time_5_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__40178\,
            in1 => \N__41490\,
            in2 => \N__31919\,
            in3 => \N__37260\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47209\,
            ce => \N__44449\,
            sr => \N__46707\
        );

    \phase_controller_slave.start_timer_hc_RNO_1_LC_12_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32150\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32166\,
            lcout => OPEN,
            ltout => \phase_controller_slave.start_timer_hc_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.start_timer_hc_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__33288\,
            in1 => \N__40802\,
            in2 => \N__31916\,
            in3 => \N__47615\,
            lcout => \phase_controller_slave.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47200\,
            ce => 'H',
            sr => \N__46716\
        );

    \phase_controller_slave.state_2_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101000110000"
        )
    port map (
            in0 => \N__32167\,
            in1 => \N__47664\,
            in2 => \N__47641\,
            in3 => \N__32151\,
            lcout => \phase_controller_slave.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47200\,
            ce => 'H',
            sr => \N__46716\
        );

    \phase_controller_slave.stoper_hc.time_passed_LC_12_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__47663\,
            in1 => \N__37076\,
            in2 => \N__34187\,
            in3 => \N__40738\,
            lcout => \phase_controller_slave.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47200\,
            ce => 'H',
            sr => \N__46716\
        );

    \phase_controller_slave.S1_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32153\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => s3_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47198\,
            ce => 'H',
            sr => \N__46723\
        );

    \phase_controller_slave.state_0_LC_12_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111000001010"
        )
    port map (
            in0 => \N__33304\,
            in1 => \N__32246\,
            in2 => \N__33248\,
            in3 => \N__32219\,
            lcout => \phase_controller_slave.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47198\,
            ce => 'H',
            sr => \N__46723\
        );

    \phase_controller_slave.state_4_LC_12_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__33305\,
            in1 => \N__33247\,
            in2 => \N__33290\,
            in3 => \N__34453\,
            lcout => \phase_controller_slave.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47198\,
            ce => 'H',
            sr => \N__46723\
        );

    \phase_controller_slave.state_3_LC_12_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000001100"
        )
    port map (
            in0 => \N__34454\,
            in1 => \N__32152\,
            in2 => \N__32171\,
            in3 => \N__33287\,
            lcout => \phase_controller_slave.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47198\,
            ce => 'H',
            sr => \N__46723\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_16_LC_12_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__41027\,
            in1 => \N__40853\,
            in2 => \N__40691\,
            in3 => \N__33374\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47194\,
            ce => 'H',
            sr => \N__46730\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_14_LC_12_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__40683\,
            in1 => \N__41028\,
            in2 => \N__40899\,
            in3 => \N__33386\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47194\,
            ce => 'H',
            sr => \N__46730\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_12_LC_12_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__41026\,
            in1 => \N__40852\,
            in2 => \N__40690\,
            in3 => \N__33398\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47194\,
            ce => 'H',
            sr => \N__46730\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_19_LC_12_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__41058\,
            in1 => \N__40682\,
            in2 => \N__40918\,
            in3 => \N__33356\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47191\,
            ce => 'H',
            sr => \N__46734\
        );

    \current_shift_inst.timer_phase.running_RNIL91O_LC_12_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__33491\,
            in1 => \N__33541\,
            in2 => \_gnd_net_\,
            in3 => \N__33514\,
            lcout => \current_shift_inst.timer_phase.N_192_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.running_RNIB31B_LC_12_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33513\,
            lcout => \current_shift_inst.timer_phase.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_12_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31955\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_clk_12mhz_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33426\,
            in2 => \_gnd_net_\,
            in3 => \N__33585\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_321_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_13_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__34960\,
            in1 => \N__42551\,
            in2 => \N__44260\,
            in3 => \N__42461\,
            lcout => measured_delay_hc_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47310\,
            ce => 'H',
            sr => \N__46604\
        );

    \current_shift_inst.meas_state_0_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111110101010"
        )
    port map (
            in0 => \N__32701\,
            in1 => \N__32385\,
            in2 => \N__32357\,
            in3 => \N__32305\,
            lcout => \current_shift_inst.meas_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47298\,
            ce => 'H',
            sr => \N__46609\
        );

    \current_shift_inst.phase_valid_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100011111000"
        )
    port map (
            in0 => \N__32304\,
            in1 => \N__32843\,
            in2 => \N__32392\,
            in3 => \N__32702\,
            lcout => \current_shift_inst.phase_validZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47298\,
            ce => 'H',
            sr => \N__46609\
        );

    \current_shift_inst.timer_s1.running_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__32352\,
            in1 => \N__32330\,
            in2 => \_gnd_net_\,
            in3 => \N__35569\,
            lcout => \current_shift_inst.timer_s1.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47298\,
            ce => 'H',
            sr => \N__46609\
        );

    \delay_measurement_inst.delay_hc_reg_1_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__42526\,
            in1 => \N__34865\,
            in2 => \N__41252\,
            in3 => \N__42099\,
            lcout => measured_delay_hc_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47298\,
            ce => 'H',
            sr => \N__46609\
        );

    \delay_measurement_inst.delay_hc_reg_31_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__42101\,
            in1 => \N__44017\,
            in2 => \_gnd_net_\,
            in3 => \N__42525\,
            lcout => measured_delay_hc_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47298\,
            ce => 'H',
            sr => \N__46609\
        );

    \delay_measurement_inst.delay_hc_reg_2_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__42527\,
            in1 => \N__34847\,
            in2 => \N__34106\,
            in3 => \N__42100\,
            lcout => measured_delay_hc_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47298\,
            ce => 'H',
            sr => \N__46609\
        );

    \current_shift_inst.stop_timer_s1_RNO_0_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32380\,
            in1 => \N__32300\,
            in2 => \N__32356\,
            in3 => \N__32696\,
            lcout => OPEN,
            ltout => \current_shift_inst.N_199_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.stop_timer_s1_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111110000"
        )
    port map (
            in0 => \N__32700\,
            in1 => \N__32308\,
            in2 => \N__32258\,
            in3 => \N__32329\,
            lcout => \current_shift_inst.stop_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47289\,
            ce => \N__40522\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNII51H_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35558\,
            in2 => \_gnd_net_\,
            in3 => \N__32327\,
            lcout => \current_shift_inst.timer_s1.N_187_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.start_timer_s1_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100001010"
        )
    port map (
            in0 => \N__32698\,
            in1 => \N__32381\,
            in2 => \N__32309\,
            in3 => \N__32351\,
            lcout => \current_shift_inst.start_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47289\,
            ce => \N__40522\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__32350\,
            in1 => \N__35559\,
            in2 => \_gnd_net_\,
            in3 => \N__32328\,
            lcout => \current_shift_inst.timer_s1.N_191_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.start_timer_phase_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011111100100010"
        )
    port map (
            in0 => \N__32697\,
            in1 => \N__32307\,
            in2 => \N__32842\,
            in3 => \N__33529\,
            lcout => \current_shift_inst.start_timer_phaseZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47289\,
            ce => \N__40522\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.stop_timer_phase_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101010110000"
        )
    port map (
            in0 => \N__32306\,
            in1 => \N__32699\,
            in2 => \N__33482\,
            in3 => \N__32838\,
            lcout => \current_shift_inst.stop_timer_phaseZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47289\,
            ce => \N__40522\,
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.stop_timer_hc_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__41930\,
            in1 => \N__35882\,
            in2 => \N__46781\,
            in3 => \N__35930\,
            lcout => \delay_measurement_inst.stop_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47282\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_13_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35080\,
            in1 => \N__35128\,
            in2 => \N__34961\,
            in3 => \N__35206\,
            lcout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto5_3_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__34099\,
            in1 => \N__41248\,
            in2 => \N__35517\,
            in3 => \N__42243\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un1_startlto5Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto6_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001100"
        )
    port map (
            in0 => \N__43954\,
            in1 => \N__34151\,
            in2 => \N__32276\,
            in3 => \N__35426\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlt8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto9_0_0_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000000110000"
        )
    port map (
            in0 => \N__34030\,
            in1 => \N__33719\,
            in2 => \N__33876\,
            in3 => \N__32444\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlt15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_9_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011111111"
        )
    port map (
            in0 => \N__35081\,
            in1 => \N__42624\,
            in2 => \N__34046\,
            in3 => \N__42092\,
            lcout => measured_delay_hc_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47274\,
            ce => 'H',
            sr => \N__46628\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_8_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__44274\,
            in1 => \N__33901\,
            in2 => \N__40439\,
            in3 => \N__33853\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_13_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35633\,
            in1 => \N__39302\,
            in2 => \N__32438\,
            in3 => \N__32435\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_5_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__42628\,
            in1 => \N__34814\,
            in2 => \N__43958\,
            in3 => \N__42421\,
            lcout => measured_delay_hc_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47263\,
            ce => 'H',
            sr => \N__46634\
        );

    \delay_measurement_inst.delay_hc_reg_14_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011111010"
        )
    port map (
            in0 => \N__42418\,
            in1 => \N__35303\,
            in2 => \N__33866\,
            in3 => \N__42625\,
            lcout => measured_delay_hc_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47263\,
            ce => 'H',
            sr => \N__46634\
        );

    \delay_measurement_inst.delay_hc_reg_15_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__42626\,
            in1 => \N__33902\,
            in2 => \N__35267\,
            in3 => \N__42419\,
            lcout => measured_delay_hc_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47263\,
            ce => 'H',
            sr => \N__46634\
        );

    \delay_measurement_inst.delay_hc_reg_16_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111101010"
        )
    port map (
            in0 => \N__42420\,
            in1 => \N__42627\,
            in2 => \N__35210\,
            in3 => \N__40429\,
            lcout => measured_delay_hc_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47263\,
            ce => 'H',
            sr => \N__46634\
        );

    \phase_controller_inst1.state_RNIR0JF_1_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43077\,
            in2 => \_gnd_net_\,
            in3 => \N__43033\,
            lcout => \phase_controller_inst1.T01_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_RNO_0_3_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__34545\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43150\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.N_86_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_3_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__32507\,
            in1 => \N__32543\,
            in2 => \N__32510\,
            in3 => \N__43175\,
            lcout => \phase_controller_inst1.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47254\,
            ce => 'H',
            sr => \N__46640\
        );

    \phase_controller_inst1.state_4_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__43151\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34544\,
            lcout => \phase_controller_inst1.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47254\,
            ce => 'H',
            sr => \N__46640\
        );

    \phase_controller_inst1.S1_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32506\,
            lcout => s1_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47254\,
            ce => 'H',
            sr => \N__46640\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35797\,
            in2 => \N__35855\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_3\,
            ltout => OPEN,
            carryin => \bfn_13_13_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            clk => \N__47246\,
            ce => \N__32741\,
            sr => \N__46647\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35776\,
            in2 => \N__35828\,
            in3 => \N__32474\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            clk => \N__47246\,
            ce => \N__32741\,
            sr => \N__46647\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35798\,
            in2 => \N__35755\,
            in3 => \N__32465\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            clk => \N__47246\,
            ce => \N__32741\,
            sr => \N__46647\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35777\,
            in2 => \N__35725\,
            in3 => \N__32456\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            clk => \N__47246\,
            ce => \N__32741\,
            sr => \N__46647\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36130\,
            in2 => \N__35756\,
            in3 => \N__32447\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            clk => \N__47246\,
            ce => \N__32741\,
            sr => \N__46647\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36109\,
            in2 => \N__35726\,
            in3 => \N__32603\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            clk => \N__47246\,
            ce => \N__32741\,
            sr => \N__46647\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36131\,
            in2 => \N__36089\,
            in3 => \N__32600\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            clk => \N__47246\,
            ce => \N__32741\,
            sr => \N__46647\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36110\,
            in2 => \N__36056\,
            in3 => \N__32588\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            clk => \N__47246\,
            ce => \N__32741\,
            sr => \N__46647\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36082\,
            in2 => \N__36025\,
            in3 => \N__32579\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_11\,
            ltout => OPEN,
            carryin => \bfn_13_14_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            clk => \N__47238\,
            ce => \N__32740\,
            sr => \N__46656\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36055\,
            in2 => \N__35998\,
            in3 => \N__32570\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            clk => \N__47238\,
            ce => \N__32740\,
            sr => \N__46656\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35971\,
            in2 => \N__36026\,
            in3 => \N__32567\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            clk => \N__47238\,
            ce => \N__32740\,
            sr => \N__46656\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35950\,
            in2 => \N__35999\,
            in3 => \N__32558\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            clk => \N__47238\,
            ce => \N__32740\,
            sr => \N__46656\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35972\,
            in2 => \N__36364\,
            in3 => \N__32549\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            clk => \N__47238\,
            ce => \N__32740\,
            sr => \N__46656\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35951\,
            in2 => \N__36337\,
            in3 => \N__32546\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            clk => \N__47238\,
            ce => \N__32740\,
            sr => \N__46656\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36310\,
            in2 => \N__36365\,
            in3 => \N__32672\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            clk => \N__47238\,
            ce => \N__32740\,
            sr => \N__46656\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36281\,
            in2 => \N__36338\,
            in3 => \N__32663\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            clk => \N__47238\,
            ce => \N__32740\,
            sr => \N__46656\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36311\,
            in2 => \N__36253\,
            in3 => \N__32654\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_19\,
            ltout => OPEN,
            carryin => \bfn_13_15_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            clk => \N__47230\,
            ce => \N__32739\,
            sr => \N__46665\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36280\,
            in2 => \N__36226\,
            in3 => \N__32645\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            clk => \N__47230\,
            ce => \N__32739\,
            sr => \N__46665\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36199\,
            in2 => \N__36254\,
            in3 => \N__32636\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            clk => \N__47230\,
            ce => \N__32739\,
            sr => \N__46665\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36178\,
            in2 => \N__36227\,
            in3 => \N__32627\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            clk => \N__47230\,
            ce => \N__32739\,
            sr => \N__46665\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36200\,
            in2 => \N__36157\,
            in3 => \N__32624\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            clk => \N__47230\,
            ce => \N__32739\,
            sr => \N__46665\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36179\,
            in2 => \N__36700\,
            in3 => \N__32615\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            clk => \N__47230\,
            ce => \N__32739\,
            sr => \N__46665\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36674\,
            in2 => \N__36158\,
            in3 => \N__32606\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            clk => \N__47230\,
            ce => \N__32739\,
            sr => \N__46665\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36647\,
            in2 => \N__36701\,
            in3 => \N__32780\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            clk => \N__47230\,
            ce => \N__32739\,
            sr => \N__46665\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36673\,
            in2 => \N__36619\,
            in3 => \N__32771\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_27\,
            ltout => OPEN,
            carryin => \bfn_13_16_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            clk => \N__47225\,
            ce => \N__32737\,
            sr => \N__46675\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36646\,
            in2 => \N__36592\,
            in3 => \N__32762\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            clk => \N__47225\,
            ce => \N__32737\,
            sr => \N__46675\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36566\,
            in2 => \N__36620\,
            in3 => \N__32753\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            clk => \N__47225\,
            ce => \N__32737\,
            sr => \N__46675\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36425\,
            in2 => \N__36593\,
            in3 => \N__32744\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\,
            clk => \N__47225\,
            ce => \N__32737\,
            sr => \N__46675\
        );

    \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32720\,
            lcout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.S1_rise_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32807\,
            in2 => \_gnd_net_\,
            in3 => \N__32815\,
            lcout => \current_shift_inst.S1_riseZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47222\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.S3_sync_prev_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32795\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.S3_sync_prevZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47222\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.S1_sync0_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32875\,
            lcout => \current_shift_inst.S1_syncZ0Z0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47222\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.S1_sync1_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32855\,
            lcout => \current_shift_inst.S1_syncZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47222\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.S3_rise_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32849\,
            in2 => \_gnd_net_\,
            in3 => \N__32794\,
            lcout => \current_shift_inst.S3_riseZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47222\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.S1_sync_prev_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32816\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.S1_sync_prevZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47222\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.S3_sync1_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32801\,
            lcout => \current_shift_inst.S3_syncZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47222\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.target_time_6_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001000101"
        )
    port map (
            in0 => \N__37350\,
            in1 => \N__40249\,
            in2 => \N__41492\,
            in3 => \N__37256\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47216\,
            ce => \N__44444\,
            sr => \N__46688\
        );

    \phase_controller_slave.stoper_tr.target_time_4_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__37255\,
            in1 => \N__41485\,
            in2 => \N__43501\,
            in3 => \N__37349\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47216\,
            ce => \N__44444\,
            sr => \N__46688\
        );

    \phase_controller_slave.stoper_tr.target_time_7_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__41482\,
            in1 => \N__37328\,
            in2 => \_gnd_net_\,
            in3 => \N__37254\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47216\,
            ce => \N__44444\,
            sr => \N__46688\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_6_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100010001"
        )
    port map (
            in0 => \N__47534\,
            in1 => \N__47707\,
            in2 => \N__47442\,
            in3 => \N__47390\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.target_time_8_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__41483\,
            in1 => \_gnd_net_\,
            in2 => \N__32978\,
            in3 => \N__37226\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47216\,
            ce => \N__44444\,
            sr => \N__46688\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_13_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41481\,
            in2 => \_gnd_net_\,
            in3 => \N__47831\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.target_time_9_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111111001101"
        )
    port map (
            in0 => \N__47391\,
            in1 => \N__47435\,
            in2 => \N__32975\,
            in3 => \N__47536\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47216\,
            ce => \N__44444\,
            sr => \N__46688\
        );

    \phase_controller_slave.stoper_tr.target_time_14_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__47535\,
            in1 => \N__41484\,
            in2 => \_gnd_net_\,
            in3 => \N__47708\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47216\,
            ce => \N__44444\,
            sr => \N__46688\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32960\,
            in2 => \N__32972\,
            in3 => \N__34365\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_13_19_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32945\,
            in2 => \N__32954\,
            in3 => \N__34345\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32930\,
            in2 => \N__32939\,
            in3 => \N__34309\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32912\,
            in2 => \N__32924\,
            in3 => \N__34279\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32894\,
            in2 => \N__32906\,
            in3 => \N__34249\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33128\,
            in2 => \N__33137\,
            in3 => \N__34726\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33110\,
            in2 => \N__33122\,
            in3 => \N__34699\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33095\,
            in2 => \N__33104\,
            in3 => \N__34666\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33077\,
            in2 => \N__33089\,
            in3 => \N__37517\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_13_20_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34636\,
            in1 => \N__33056\,
            in2 => \N__33071\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33032\,
            in2 => \N__33050\,
            in3 => \N__34607\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33008\,
            in2 => \N__33026\,
            in3 => \N__37655\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32984\,
            in2 => \N__33002\,
            in3 => \N__37541\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33203\,
            in2 => \N__33218\,
            in3 => \N__38324\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33179\,
            in2 => \N__33197\,
            in3 => \N__37679\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33173\,
            in2 => \N__44471\,
            in3 => \N__37631\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33167\,
            in2 => \N__33146\,
            in3 => \N__38222\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_13_21_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_13_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33161\,
            in2 => \N__33323\,
            in3 => \N__38198\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_13_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33155\,
            in2 => \N__33314\,
            in3 => \N__37760\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33149\,
            lcout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.target_time_17_LC_13_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__43297\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47206\,
            ce => \N__44445\,
            sr => \N__46711\
        );

    \phase_controller_slave.stoper_tr.target_time_18_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43211\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47206\,
            ce => \N__44445\,
            sr => \N__46711\
        );

    \phase_controller_slave.stoper_tr.target_time_19_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__41576\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47206\,
            ce => \N__44445\,
            sr => \N__46711\
        );

    \phase_controller_slave.start_timer_tr_RNO_0_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33242\,
            in2 => \_gnd_net_\,
            in3 => \N__33303\,
            lcout => OPEN,
            ltout => \phase_controller_slave.N_210_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.start_timer_tr_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110111001100"
        )
    port map (
            in0 => \N__33289\,
            in1 => \N__33266\,
            in2 => \N__33254\,
            in3 => \N__37951\,
            lcout => \phase_controller_slave.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47202\,
            ce => 'H',
            sr => \N__46717\
        );

    \phase_controller_slave.stoper_tr.stoper_state_RNI38A6_0_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37859\,
            in2 => \_gnd_net_\,
            in3 => \N__38145\,
            lcout => \phase_controller_slave.stoper_tr.time_passed11\,
            ltout => \phase_controller_slave.stoper_tr.time_passed11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.time_passed_LC_13_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010111000"
        )
    port map (
            in0 => \N__33243\,
            in1 => \N__33224\,
            in2 => \N__33251\,
            in3 => \N__34410\,
            lcout => \phase_controller_slave.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47202\,
            ce => 'H',
            sr => \N__46717\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_11_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__37861\,
            in1 => \N__38147\,
            in2 => \N__37998\,
            in3 => \N__34592\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47202\,
            ce => 'H',
            sr => \N__46717\
        );

    \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__37947\,
            in1 => \N__37860\,
            in2 => \_gnd_net_\,
            in3 => \N__38146\,
            lcout => \phase_controller_slave.stoper_tr.time_passed_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_13_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34208\,
            in2 => \N__38291\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_23_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_13_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38252\,
            in2 => \_gnd_net_\,
            in3 => \N__33350\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34577\,
            in2 => \N__36833\,
            in3 => \N__33347\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_13_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37601\,
            in2 => \_gnd_net_\,
            in3 => \N__33344\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37568\,
            in2 => \_gnd_net_\,
            in3 => \N__33341\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_13_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37487\,
            in2 => \_gnd_net_\,
            in3 => \N__33338\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_13_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36749\,
            in2 => \_gnd_net_\,
            in3 => \N__33335\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_13_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36725\,
            in2 => \_gnd_net_\,
            in3 => \N__33332\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38509\,
            in2 => \_gnd_net_\,
            in3 => \N__33329\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9\,
            ltout => OPEN,
            carryin => \bfn_13_24_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37733\,
            in2 => \_gnd_net_\,
            in3 => \N__33326\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_13_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37705\,
            in2 => \_gnd_net_\,
            in3 => \N__33401\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_13_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36961\,
            in2 => \_gnd_net_\,
            in3 => \N__33392\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_13_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36934\,
            in2 => \_gnd_net_\,
            in3 => \N__33389\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_13_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36895\,
            in2 => \_gnd_net_\,
            in3 => \N__33380\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_13_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38476\,
            in2 => \_gnd_net_\,
            in3 => \N__33377\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_13_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37174\,
            in2 => \_gnd_net_\,
            in3 => \N__33368\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_13_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37150\,
            in2 => \_gnd_net_\,
            in3 => \N__33365\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17\,
            ltout => OPEN,
            carryin => \bfn_13_25_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_13_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37126\,
            in2 => \_gnd_net_\,
            in3 => \N__33362\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_13_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37099\,
            in2 => \_gnd_net_\,
            in3 => \N__33359\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.running_LC_13_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__33542\,
            in1 => \N__33515\,
            in2 => \_gnd_net_\,
            in3 => \N__33489\,
            lcout => \current_shift_inst.timer_phase.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47192\,
            ce => 'H',
            sr => \N__46735\
        );

    \current_shift_inst.timer_phase.running_RNIC90O_LC_13_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33512\,
            in2 => \_gnd_net_\,
            in3 => \N__33490\,
            lcout => \current_shift_inst.timer_phase.N_188_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.S2_LC_13_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43100\,
            lcout => s2_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47189\,
            ce => 'H',
            sr => \N__46739\
        );

    \delay_measurement_inst.delay_hc_timer.running_LC_14_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__35903\,
            in1 => \N__33431\,
            in2 => \_gnd_net_\,
            in3 => \N__33591\,
            lcout => \delay_measurement_inst.delay_hc_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47326\,
            ce => 'H',
            sr => \N__46596\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJG9N1_1_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35538\,
            in1 => \N__34839\,
            in2 => \N__34813\,
            in3 => \N__34858\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINGQU3_9_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100101010"
        )
    port map (
            in0 => \N__35075\,
            in1 => \N__34871\,
            in2 => \N__33434\,
            in3 => \N__35259\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_2_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__33593\,
            in1 => \N__35899\,
            in2 => \_gnd_net_\,
            in3 => \N__33427\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_322_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOHNN2_6_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101000001010"
        )
    port map (
            in0 => \N__33691\,
            in1 => \N__35117\,
            in2 => \N__35076\,
            in3 => \N__33611\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1LC84_14_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111000000000"
        )
    port map (
            in0 => \N__35302\,
            in1 => \N__35257\,
            in2 => \N__33404\,
            in3 => \N__33554\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt30_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41792\,
            in2 => \_gnd_net_\,
            in3 => \N__41697\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0\,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_10_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__33620\,
            in1 => \N__34823\,
            in2 => \N__33605\,
            in3 => \N__33560\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOVQ9D_14_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__35597\,
            in1 => \N__33656\,
            in2 => \N__33602\,
            in3 => \N__33599\,
            lcout => \delay_measurement_inst.un1_elapsed_time_hc\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__33592\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI93LG1_14_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__35249\,
            in1 => \N__35288\,
            in2 => \_gnd_net_\,
            in3 => \N__33553\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI537G_17_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__42205\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42481\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4UNN2_4_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__33569\,
            in1 => \N__35449\,
            in2 => \N__33563\,
            in3 => \N__34803\,
            lcout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35002\,
            in1 => \N__34947\,
            in2 => \N__34983\,
            in3 => \N__35031\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__42204\,
            in1 => \N__42480\,
            in2 => \N__42129\,
            in3 => \N__35194\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ0JH1_6_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41793\,
            in1 => \N__41698\,
            in2 => \N__35124\,
            in3 => \N__35256\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52G18_14_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100000000"
        )
    port map (
            in0 => \N__33692\,
            in1 => \N__33680\,
            in2 => \N__33671\,
            in3 => \N__33668\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP8VO1_20_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__35144\,
            in1 => \N__35156\,
            in2 => \N__35171\,
            in3 => \N__33646\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_1\,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5483B_31_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__35593\,
            in1 => \N__35315\,
            in2 => \N__33662\,
            in3 => \N__33629\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto31_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35143\,
            in2 => \_gnd_net_\,
            in3 => \N__35155\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINN412_20_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__33647\,
            in1 => \N__35313\,
            in2 => \N__33659\,
            in3 => \N__35170\,
            lcout => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35351\,
            in1 => \N__35360\,
            in2 => \N__35342\,
            in3 => \N__35369\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5483B_0_31_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010011"
        )
    port map (
            in0 => \N__35592\,
            in1 => \N__35314\,
            in2 => \N__33638\,
            in3 => \N__33628\,
            lcout => \delay_measurement_inst.delay_hc_reg3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOJD01_11_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35260\,
            in1 => \N__34984\,
            in2 => \N__35012\,
            in3 => \N__35298\,
            lcout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_10_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__42621\,
            in1 => \N__35039\,
            in2 => \N__35677\,
            in3 => \N__42378\,
            lcout => measured_delay_hc_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47283\,
            ce => 'H',
            sr => \N__46618\
        );

    \delay_measurement_inst.delay_hc_reg_11_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__42622\,
            in1 => \N__35011\,
            in2 => \N__39350\,
            in3 => \N__42379\,
            lcout => measured_delay_hc_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47283\,
            ce => 'H',
            sr => \N__46618\
        );

    \delay_measurement_inst.delay_hc_reg_12_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__42380\,
            in1 => \N__34985\,
            in2 => \N__39405\,
            in3 => \N__42623\,
            lcout => measured_delay_hc_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47283\,
            ce => 'H',
            sr => \N__46618\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto13_3_1_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__39379\,
            in1 => \N__39331\,
            in2 => \N__44273\,
            in3 => \N__35657\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un1_startlto13_3Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto13_3_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001110000"
        )
    port map (
            in0 => \N__34029\,
            in1 => \N__41756\,
            in2 => \N__33722\,
            in3 => \N__41671\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_26_1_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__42019\,
            in1 => \N__33711\,
            in2 => \N__42682\,
            in3 => \N__42049\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_20_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__33713\,
            in1 => \N__42620\,
            in2 => \_gnd_net_\,
            in3 => \N__42417\,
            lcout => measured_delay_hc_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47275\,
            ce => 'H',
            sr => \N__46629\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto30_2_0_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__42020\,
            in1 => \N__33712\,
            in2 => \N__42683\,
            in3 => \N__41876\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un1_startlto30_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto30_3_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001110000"
        )
    port map (
            in0 => \N__33903\,
            in1 => \N__35576\,
            in2 => \N__33701\,
            in3 => \N__33698\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlt31_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.stoper_state_RNII60D_0_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__38045\,
            in1 => \N__37826\,
            in2 => \_gnd_net_\,
            in3 => \N__38117\,
            lcout => \phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.start_timer_tr_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__34905\,
            in1 => \N__33833\,
            in2 => \_gnd_net_\,
            in3 => \N__33805\,
            lcout => \delay_measurement_inst.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47255\,
            ce => 'H',
            sr => \N__46641\
        );

    \delay_measurement_inst.prev_tr_sig_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34906\,
            lcout => \delay_measurement_inst.prev_tr_sigZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47255\,
            ce => 'H',
            sr => \N__46641\
        );

    \delay_measurement_inst.tr_state_RNIMR6L_0_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__34904\,
            in1 => \N__33832\,
            in2 => \_gnd_net_\,
            in3 => \N__33804\,
            lcout => \delay_measurement_inst.tr_state_RNIMR6LZ0Z_0\,
            ltout => \delay_measurement_inst.tr_state_RNIMR6LZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.stop_timer_tr_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33791\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.stop_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47255\,
            ce => 'H',
            sr => \N__46641\
        );

    \delay_measurement_inst.delay_tr_timer.running_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101111100001010"
        )
    port map (
            in0 => \N__39255\,
            in1 => \_gnd_net_\,
            in2 => \N__37405\,
            in3 => \N__37378\,
            lcout => \delay_measurement_inst.delay_tr_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47255\,
            ce => 'H',
            sr => \N__46641\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37398\,
            in2 => \_gnd_net_\,
            in3 => \N__39254\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_323_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.T01_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010111010"
        )
    port map (
            in0 => \N__33788\,
            in1 => \N__43117\,
            in2 => \N__34474\,
            in3 => \N__43152\,
            lcout => shift_flag_start,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47255\,
            ce => 'H',
            sr => \N__46641\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33755\,
            lcout => \current_shift_inst.un4_control_input_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33740\,
            lcout => \current_shift_inst.un4_control_input_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33986\,
            lcout => \current_shift_inst.un4_control_input_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33968\,
            lcout => \current_shift_inst.un4_control_input_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33950\,
            lcout => \current_shift_inst.un4_control_input_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_10_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47605\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39469\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47239\,
            ce => \N__46858\,
            sr => \N__46657\
        );

    \phase_controller_inst1.stoper_tr.target_time_12_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47606\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39496\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47239\,
            ce => \N__46858\,
            sr => \N__46657\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33932\,
            lcout => \current_shift_inst.un4_control_input_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.target_time_0_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__44164\,
            in1 => \N__43853\,
            in2 => \N__42259\,
            in3 => \N__40336\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47231\,
            ce => \N__43700\,
            sr => \N__46666\
        );

    \phase_controller_slave.stoper_hc.target_time_15_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__43855\,
            in1 => \N__44166\,
            in2 => \_gnd_net_\,
            in3 => \N__33917\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47231\,
            ce => \N__43700\,
            sr => \N__46666\
        );

    \phase_controller_slave.stoper_hc.target_time_14_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__43854\,
            in1 => \N__44165\,
            in2 => \_gnd_net_\,
            in3 => \N__33877\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47231\,
            ce => \N__43700\,
            sr => \N__46666\
        );

    \phase_controller_slave.stoper_hc.target_timeZ0Z_6_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001000000011"
        )
    port map (
            in0 => \N__34165\,
            in1 => \N__40335\,
            in2 => \N__44198\,
            in3 => \N__43852\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ1Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47231\,
            ce => \N__43700\,
            sr => \N__46666\
        );

    \phase_controller_slave.stoper_hc.target_time_10_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__44167\,
            in1 => \N__35670\,
            in2 => \_gnd_net_\,
            in3 => \N__43856\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47226\,
            ce => \N__43687\,
            sr => \N__46676\
        );

    \phase_controller_slave.stoper_hc.target_time_3_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110101000"
        )
    port map (
            in0 => \N__43860\,
            in1 => \N__40318\,
            in2 => \N__35518\,
            in3 => \N__44173\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47226\,
            ce => \N__43687\,
            sr => \N__46676\
        );

    \phase_controller_slave.stoper_hc.target_time_12_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__44169\,
            in1 => \N__39406\,
            in2 => \_gnd_net_\,
            in3 => \N__43858\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47226\,
            ce => \N__43687\,
            sr => \N__46676\
        );

    \phase_controller_slave.stoper_hc.target_time_11_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__43857\,
            in1 => \N__44168\,
            in2 => \_gnd_net_\,
            in3 => \N__39353\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47226\,
            ce => \N__43687\,
            sr => \N__46676\
        );

    \phase_controller_slave.stoper_hc.target_time_2_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__40316\,
            in1 => \N__34115\,
            in2 => \N__44199\,
            in3 => \N__43859\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47226\,
            ce => \N__43687\,
            sr => \N__46676\
        );

    \phase_controller_slave.stoper_hc.target_time_9_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000110001"
        )
    port map (
            in0 => \N__43863\,
            in1 => \N__44178\,
            in2 => \N__34055\,
            in3 => \N__40319\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47226\,
            ce => \N__43687\,
            sr => \N__46676\
        );

    \phase_controller_slave.stoper_hc.target_time_4_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__40317\,
            in1 => \N__35427\,
            in2 => \N__44200\,
            in3 => \N__43861\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47226\,
            ce => \N__43687\,
            sr => \N__46676\
        );

    \phase_controller_slave.stoper_hc.target_time_7_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__43862\,
            in1 => \N__44177\,
            in2 => \_gnd_net_\,
            in3 => \N__41675\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47226\,
            ce => \N__43687\,
            sr => \N__46676\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_7_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__40663\,
            in1 => \N__40860\,
            in2 => \N__41029\,
            in3 => \N__33998\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47223\,
            ce => 'H',
            sr => \N__46681\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_8_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__40859\,
            in1 => \N__41000\,
            in2 => \N__40667\,
            in3 => \N__34199\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47223\,
            ce => 'H',
            sr => \N__46681\
        );

    \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__40858\,
            in1 => \_gnd_net_\,
            in2 => \N__40666\,
            in3 => \N__40999\,
            lcout => \phase_controller_slave.stoper_hc.time_passed_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34439\,
            in1 => \N__34369\,
            in2 => \_gnd_net_\,
            in3 => \N__34411\,
            lcout => OPEN,
            ltout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_1_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__38024\,
            in1 => \N__37892\,
            in2 => \N__34172\,
            in3 => \N__38143\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47223\,
            ce => 'H',
            sr => \N__46681\
        );

    \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_0_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__40998\,
            in1 => \N__40640\,
            in2 => \_gnd_net_\,
            in3 => \N__40857\,
            lcout => \phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_10_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__37858\,
            in1 => \N__38142\,
            in2 => \N__38047\,
            in3 => \N__34619\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47223\,
            ce => 'H',
            sr => \N__46681\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_2_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010000010"
        )
    port map (
            in0 => \N__34334\,
            in1 => \N__37875\,
            in2 => \N__38046\,
            in3 => \N__38173\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47217\,
            ce => 'H',
            sr => \N__46689\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_3_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100011000100"
        )
    port map (
            in0 => \N__37873\,
            in1 => \N__34298\,
            in2 => \N__38179\,
            in3 => \N__38022\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47217\,
            ce => 'H',
            sr => \N__46689\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_4_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__38015\,
            in1 => \N__37876\,
            in2 => \N__34268\,
            in3 => \N__38165\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47217\,
            ce => 'H',
            sr => \N__46689\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_5_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100011000100"
        )
    port map (
            in0 => \N__37874\,
            in1 => \N__34745\,
            in2 => \N__38180\,
            in3 => \N__38023\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47217\,
            ce => 'H',
            sr => \N__46689\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_3_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__41053\,
            in1 => \N__40664\,
            in2 => \N__40914\,
            in3 => \N__34238\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47217\,
            ce => 'H',
            sr => \N__46689\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_7_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__38164\,
            in1 => \N__38018\,
            in2 => \N__37899\,
            in3 => \N__34688\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47217\,
            ce => 'H',
            sr => \N__46689\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_8_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__38016\,
            in1 => \N__37877\,
            in2 => \N__34655\,
            in3 => \N__38166\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47217\,
            ce => 'H',
            sr => \N__46689\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_6_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__38163\,
            in1 => \N__38017\,
            in2 => \N__37898\,
            in3 => \N__34715\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47217\,
            ce => 'H',
            sr => \N__46689\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_3_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__43205\,
            in1 => \N__41568\,
            in2 => \N__43296\,
            in3 => \N__44386\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_5_3_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__40164\,
            in1 => \N__43497\,
            in2 => \N__34226\,
            in3 => \N__47824\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_5Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_15_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__44387\,
            in1 => \N__43206\,
            in2 => \N__41575\,
            in3 => \N__43289\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.stoper_state_RNIDEUE_0_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41022\,
            in2 => \_gnd_net_\,
            in3 => \N__40628\,
            lcout => \phase_controller_slave.stoper_hc.time_passed11\,
            ltout => \phase_controller_slave.stoper_hc.time_passed11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34211\,
            in3 => \N__40716\,
            lcout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSR_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__40717\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37062\,
            lcout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1B6_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34432\,
            in2 => \_gnd_net_\,
            in3 => \N__34403\,
            lcout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.un1_start_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__34557\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34475\,
            lcout => \phase_controller_slave.un1_startZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34431\,
            in2 => \_gnd_net_\,
            in3 => \N__34402\,
            lcout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34379\,
            in2 => \N__34373\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_22_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_14_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34349\,
            in2 => \_gnd_net_\,
            in3 => \N__34325\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_14_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34322\,
            in2 => \N__34316\,
            in3 => \N__34286\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34283\,
            in2 => \_gnd_net_\,
            in3 => \N__34256\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_14_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34253\,
            in2 => \_gnd_net_\,
            in3 => \N__34733\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_14_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34730\,
            in2 => \_gnd_net_\,
            in3 => \N__34706\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_14_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34703\,
            in2 => \_gnd_net_\,
            in3 => \N__34673\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_14_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34670\,
            in2 => \_gnd_net_\,
            in3 => \N__34643\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37513\,
            in2 => \_gnd_net_\,
            in3 => \N__34640\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9\,
            ltout => OPEN,
            carryin => \bfn_14_23_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_14_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34637\,
            in2 => \_gnd_net_\,
            in3 => \N__34610\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_14_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34606\,
            in2 => \_gnd_net_\,
            in3 => \N__34586\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_14_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37651\,
            in2 => \_gnd_net_\,
            in3 => \N__34583\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_14_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37537\,
            in2 => \_gnd_net_\,
            in3 => \N__34580\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_14_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38320\,
            in2 => \_gnd_net_\,
            in3 => \N__34781\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_14_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37675\,
            in2 => \_gnd_net_\,
            in3 => \N__34778\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_14_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37627\,
            in2 => \_gnd_net_\,
            in3 => \N__34775\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_14_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38218\,
            in2 => \_gnd_net_\,
            in3 => \N__34772\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17\,
            ltout => OPEN,
            carryin => \bfn_14_24_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_14_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38194\,
            in2 => \_gnd_net_\,
            in3 => \N__34769\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_14_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37756\,
            in2 => \_gnd_net_\,
            in3 => \N__34766\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_13_LC_14_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__41066\,
            in1 => \N__40680\,
            in2 => \N__40909\,
            in3 => \N__34763\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47196\,
            ce => 'H',
            sr => \N__46726\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_17_LC_14_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__41067\,
            in1 => \N__40681\,
            in2 => \N__40910\,
            in3 => \N__34757\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47196\,
            ce => 'H',
            sr => \N__46726\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_18_LC_14_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__40679\,
            in1 => \N__41068\,
            in2 => \N__40917\,
            in3 => \N__34751\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47196\,
            ce => 'H',
            sr => \N__46726\
        );

    \SB_DFF_inst_DELAY_TR1_LC_15_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__34925\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => delay_tr_d1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47334\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_DELAY_TR2_LC_15_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34916\,
            lcout => delay_tr_d2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47334\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHUIH1_4_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41696\,
            in1 => \N__35448\,
            in2 => \N__41797\,
            in3 => \N__35258\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38456\,
            lcout => \delay_measurement_inst.elapsed_time_hc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47327\,
            ce => \N__35695\,
            sr => \N__46597\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38435\,
            lcout => \delay_measurement_inst.elapsed_time_hc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47327\,
            ce => \N__35695\,
            sr => \N__46597\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOKRB1_10_LC_15_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__35539\,
            in1 => \N__42130\,
            in2 => \N__35038\,
            in3 => \N__34840\,
            lcout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38455\,
            in2 => \N__38413\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.elapsed_time_hc_3\,
            ltout => OPEN,
            carryin => \bfn_15_7_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__47319\,
            ce => \N__35696\,
            sr => \N__46600\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38434\,
            in2 => \N__38389\,
            in3 => \N__34817\,
            lcout => \delay_measurement_inst.elapsed_time_hc_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__47319\,
            ce => \N__35696\,
            sr => \N__46600\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38364\,
            in2 => \N__38414\,
            in3 => \N__34784\,
            lcout => \delay_measurement_inst.elapsed_time_hc_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__47319\,
            ce => \N__35696\,
            sr => \N__46600\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38346\,
            in2 => \N__38390\,
            in3 => \N__35090\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__47319\,
            ce => \N__35696\,
            sr => \N__46600\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38365\,
            in2 => \N__38698\,
            in3 => \N__35087\,
            lcout => \delay_measurement_inst.elapsed_time_hc_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__47319\,
            ce => \N__35696\,
            sr => \N__46600\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38347\,
            in2 => \N__38674\,
            in3 => \N__35084\,
            lcout => \delay_measurement_inst.elapsed_time_hc_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__47319\,
            ce => \N__35696\,
            sr => \N__46600\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38651\,
            in2 => \N__38699\,
            in3 => \N__35042\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__47319\,
            ce => \N__35696\,
            sr => \N__46600\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38627\,
            in2 => \N__38675\,
            in3 => \N__35015\,
            lcout => \delay_measurement_inst.elapsed_time_hc_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__47319\,
            ce => \N__35696\,
            sr => \N__46600\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38650\,
            in2 => \N__38602\,
            in3 => \N__34988\,
            lcout => \delay_measurement_inst.elapsed_time_hc_11\,
            ltout => OPEN,
            carryin => \bfn_15_8_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__47311\,
            ce => \N__35697\,
            sr => \N__46605\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38626\,
            in2 => \N__38578\,
            in3 => \N__34964\,
            lcout => \delay_measurement_inst.elapsed_time_hc_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__47311\,
            ce => \N__35697\,
            sr => \N__46605\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38553\,
            in2 => \N__38603\,
            in3 => \N__34928\,
            lcout => \delay_measurement_inst.elapsed_time_hc_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__47311\,
            ce => \N__35697\,
            sr => \N__46605\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38535\,
            in2 => \N__38579\,
            in3 => \N__35270\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__47311\,
            ce => \N__35697\,
            sr => \N__46605\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38554\,
            in2 => \N__38878\,
            in3 => \N__35213\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__47311\,
            ce => \N__35697\,
            sr => \N__46605\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38536\,
            in2 => \N__38854\,
            in3 => \N__35183\,
            lcout => \delay_measurement_inst.elapsed_time_hc_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__47311\,
            ce => \N__35697\,
            sr => \N__46605\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38831\,
            in2 => \N__38879\,
            in3 => \N__35180\,
            lcout => \delay_measurement_inst.elapsed_time_hc_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__47311\,
            ce => \N__35697\,
            sr => \N__46605\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38807\,
            in2 => \N__38855\,
            in3 => \N__35177\,
            lcout => \delay_measurement_inst.elapsed_time_hc_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__47311\,
            ce => \N__35697\,
            sr => \N__46605\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38830\,
            in2 => \N__38782\,
            in3 => \N__35174\,
            lcout => \delay_measurement_inst.elapsed_time_hc_19\,
            ltout => OPEN,
            carryin => \bfn_15_9_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__47299\,
            ce => \N__35698\,
            sr => \N__46610\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38806\,
            in2 => \N__38758\,
            in3 => \N__35159\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__47299\,
            ce => \N__35698\,
            sr => \N__46610\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38733\,
            in2 => \N__38783\,
            in3 => \N__35147\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__47299\,
            ce => \N__35698\,
            sr => \N__46610\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38715\,
            in2 => \N__38759\,
            in3 => \N__35132\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__47299\,
            ce => \N__35698\,
            sr => \N__46610\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38734\,
            in2 => \N__39232\,
            in3 => \N__35363\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__47299\,
            ce => \N__35698\,
            sr => \N__46610\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38716\,
            in2 => \N__39208\,
            in3 => \N__35354\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__47299\,
            ce => \N__35698\,
            sr => \N__46610\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39185\,
            in2 => \N__39233\,
            in3 => \N__35345\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__47299\,
            ce => \N__35698\,
            sr => \N__46610\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39161\,
            in2 => \N__39209\,
            in3 => \N__35333\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__47299\,
            ce => \N__35698\,
            sr => \N__46610\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39184\,
            in2 => \N__39136\,
            in3 => \N__35330\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\,
            ltout => OPEN,
            carryin => \bfn_15_10_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__47290\,
            ce => \N__35699\,
            sr => \N__46614\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39160\,
            in2 => \N__39112\,
            in3 => \N__35327\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__47290\,
            ce => \N__35699\,
            sr => \N__46614\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39088\,
            in2 => \N__39137\,
            in3 => \N__35324\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__47290\,
            ce => \N__35699\,
            sr => \N__46614\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38935\,
            in2 => \N__39113\,
            in3 => \N__35321\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__47290\,
            ce => \N__35699\,
            sr => \N__46614\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35318\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47290\,
            ce => \N__35699\,
            sr => \N__46614\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41660\,
            in1 => \N__43955\,
            in2 => \N__41763\,
            in3 => \N__35656\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35624\,
            in1 => \N__35618\,
            in2 => \N__35612\,
            in3 => \N__35603\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__40440\,
            in1 => \N__42183\,
            in2 => \N__42053\,
            in3 => \N__42339\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIUKI8_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35570\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.timer_s1.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_3_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__42649\,
            in1 => \N__35543\,
            in2 => \N__35500\,
            in3 => \N__42442\,
            lcout => measured_delay_hc_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47276\,
            ce => 'H',
            sr => \N__46630\
        );

    \delay_measurement_inst.delay_hc_reg_4_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__42443\,
            in1 => \N__42650\,
            in2 => \N__35422\,
            in3 => \N__35453\,
            lcout => measured_delay_hc_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47276\,
            ce => 'H',
            sr => \N__46630\
        );

    \delay_measurement_inst.delay_tr_reg_15_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__45159\,
            in1 => \N__47487\,
            in2 => \N__47806\,
            in3 => \N__47723\,
            lcout => measured_delay_tr_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47276\,
            ce => 'H',
            sr => \N__46630\
        );

    \delay_measurement_inst.delay_tr_reg_7_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__47724\,
            in1 => \N__43594\,
            in2 => \N__37313\,
            in3 => \N__44717\,
            lcout => measured_delay_tr_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47276\,
            ce => 'H',
            sr => \N__46630\
        );

    \delay_measurement_inst.delay_tr_reg_8_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__44663\,
            in1 => \N__37202\,
            in2 => \N__43603\,
            in3 => \N__47725\,
            lcout => measured_delay_tr_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47276\,
            ce => 'H',
            sr => \N__46630\
        );

    \delay_measurement_inst.start_timer_hc_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100110101010"
        )
    port map (
            in0 => \N__35929\,
            in1 => \N__35868\,
            in2 => \_gnd_net_\,
            in3 => \N__41931\,
            lcout => \delay_measurement_inst.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47276\,
            ce => 'H',
            sr => \N__46630\
        );

    \delay_measurement_inst.prev_hc_sig_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__41932\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.prev_hc_sigZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47276\,
            ce => 'H',
            sr => \N__46630\
        );

    \current_shift_inst.timer_s1.counter_0_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36533\,
            in1 => \N__35850\,
            in2 => \_gnd_net_\,
            in3 => \N__35831\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_15_13_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_0\,
            clk => \N__47264\,
            ce => \N__36409\,
            sr => \N__46635\
        );

    \current_shift_inst.timer_s1.counter_1_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36541\,
            in1 => \N__35820\,
            in2 => \_gnd_net_\,
            in3 => \N__35801\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_0\,
            carryout => \current_shift_inst.timer_s1.counter_cry_1\,
            clk => \N__47264\,
            ce => \N__36409\,
            sr => \N__46635\
        );

    \current_shift_inst.timer_s1.counter_2_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36534\,
            in1 => \N__35796\,
            in2 => \_gnd_net_\,
            in3 => \N__35780\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_1\,
            carryout => \current_shift_inst.timer_s1.counter_cry_2\,
            clk => \N__47264\,
            ce => \N__36409\,
            sr => \N__46635\
        );

    \current_shift_inst.timer_s1.counter_3_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36542\,
            in1 => \N__35775\,
            in2 => \_gnd_net_\,
            in3 => \N__35759\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_2\,
            carryout => \current_shift_inst.timer_s1.counter_cry_3\,
            clk => \N__47264\,
            ce => \N__36409\,
            sr => \N__46635\
        );

    \current_shift_inst.timer_s1.counter_4_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36535\,
            in1 => \N__35743\,
            in2 => \_gnd_net_\,
            in3 => \N__35729\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_3\,
            carryout => \current_shift_inst.timer_s1.counter_cry_4\,
            clk => \N__47264\,
            ce => \N__36409\,
            sr => \N__46635\
        );

    \current_shift_inst.timer_s1.counter_5_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36543\,
            in1 => \N__35718\,
            in2 => \_gnd_net_\,
            in3 => \N__35702\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_4\,
            carryout => \current_shift_inst.timer_s1.counter_cry_5\,
            clk => \N__47264\,
            ce => \N__36409\,
            sr => \N__46635\
        );

    \current_shift_inst.timer_s1.counter_6_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36536\,
            in1 => \N__36129\,
            in2 => \_gnd_net_\,
            in3 => \N__36113\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_5\,
            carryout => \current_shift_inst.timer_s1.counter_cry_6\,
            clk => \N__47264\,
            ce => \N__36409\,
            sr => \N__46635\
        );

    \current_shift_inst.timer_s1.counter_7_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36544\,
            in1 => \N__36108\,
            in2 => \_gnd_net_\,
            in3 => \N__36092\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_6\,
            carryout => \current_shift_inst.timer_s1.counter_cry_7\,
            clk => \N__47264\,
            ce => \N__36409\,
            sr => \N__46635\
        );

    \current_shift_inst.timer_s1.counter_8_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36548\,
            in1 => \N__36078\,
            in2 => \_gnd_net_\,
            in3 => \N__36059\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_15_14_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_8\,
            clk => \N__47256\,
            ce => \N__36407\,
            sr => \N__46642\
        );

    \current_shift_inst.timer_s1.counter_9_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36540\,
            in1 => \N__36045\,
            in2 => \_gnd_net_\,
            in3 => \N__36029\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_8\,
            carryout => \current_shift_inst.timer_s1.counter_cry_9\,
            clk => \N__47256\,
            ce => \N__36407\,
            sr => \N__46642\
        );

    \current_shift_inst.timer_s1.counter_10_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36545\,
            in1 => \N__36018\,
            in2 => \_gnd_net_\,
            in3 => \N__36002\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_9\,
            carryout => \current_shift_inst.timer_s1.counter_cry_10\,
            clk => \N__47256\,
            ce => \N__36407\,
            sr => \N__46642\
        );

    \current_shift_inst.timer_s1.counter_11_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36537\,
            in1 => \N__35991\,
            in2 => \_gnd_net_\,
            in3 => \N__35975\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_10\,
            carryout => \current_shift_inst.timer_s1.counter_cry_11\,
            clk => \N__47256\,
            ce => \N__36407\,
            sr => \N__46642\
        );

    \current_shift_inst.timer_s1.counter_12_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36546\,
            in1 => \N__35970\,
            in2 => \_gnd_net_\,
            in3 => \N__35954\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_11\,
            carryout => \current_shift_inst.timer_s1.counter_cry_12\,
            clk => \N__47256\,
            ce => \N__36407\,
            sr => \N__46642\
        );

    \current_shift_inst.timer_s1.counter_13_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36538\,
            in1 => \N__35949\,
            in2 => \_gnd_net_\,
            in3 => \N__35933\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_12\,
            carryout => \current_shift_inst.timer_s1.counter_cry_13\,
            clk => \N__47256\,
            ce => \N__36407\,
            sr => \N__46642\
        );

    \current_shift_inst.timer_s1.counter_14_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36547\,
            in1 => \N__36357\,
            in2 => \_gnd_net_\,
            in3 => \N__36341\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_13\,
            carryout => \current_shift_inst.timer_s1.counter_cry_14\,
            clk => \N__47256\,
            ce => \N__36407\,
            sr => \N__46642\
        );

    \current_shift_inst.timer_s1.counter_15_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36539\,
            in1 => \N__36330\,
            in2 => \_gnd_net_\,
            in3 => \N__36314\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_14\,
            carryout => \current_shift_inst.timer_s1.counter_cry_15\,
            clk => \N__47256\,
            ce => \N__36407\,
            sr => \N__46642\
        );

    \current_shift_inst.timer_s1.counter_16_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36519\,
            in1 => \N__36303\,
            in2 => \_gnd_net_\,
            in3 => \N__36284\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_15_15_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_16\,
            clk => \N__47247\,
            ce => \N__36410\,
            sr => \N__46648\
        );

    \current_shift_inst.timer_s1.counter_17_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36523\,
            in1 => \N__36276\,
            in2 => \_gnd_net_\,
            in3 => \N__36257\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_16\,
            carryout => \current_shift_inst.timer_s1.counter_cry_17\,
            clk => \N__47247\,
            ce => \N__36410\,
            sr => \N__46648\
        );

    \current_shift_inst.timer_s1.counter_18_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36520\,
            in1 => \N__36246\,
            in2 => \_gnd_net_\,
            in3 => \N__36230\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_17\,
            carryout => \current_shift_inst.timer_s1.counter_cry_18\,
            clk => \N__47247\,
            ce => \N__36410\,
            sr => \N__46648\
        );

    \current_shift_inst.timer_s1.counter_19_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36524\,
            in1 => \N__36219\,
            in2 => \_gnd_net_\,
            in3 => \N__36203\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_18\,
            carryout => \current_shift_inst.timer_s1.counter_cry_19\,
            clk => \N__47247\,
            ce => \N__36410\,
            sr => \N__46648\
        );

    \current_shift_inst.timer_s1.counter_20_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36521\,
            in1 => \N__36198\,
            in2 => \_gnd_net_\,
            in3 => \N__36182\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_19\,
            carryout => \current_shift_inst.timer_s1.counter_cry_20\,
            clk => \N__47247\,
            ce => \N__36410\,
            sr => \N__46648\
        );

    \current_shift_inst.timer_s1.counter_21_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36525\,
            in1 => \N__36177\,
            in2 => \_gnd_net_\,
            in3 => \N__36161\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_20\,
            carryout => \current_shift_inst.timer_s1.counter_cry_21\,
            clk => \N__47247\,
            ce => \N__36410\,
            sr => \N__46648\
        );

    \current_shift_inst.timer_s1.counter_22_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36522\,
            in1 => \N__36150\,
            in2 => \_gnd_net_\,
            in3 => \N__36134\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_21\,
            carryout => \current_shift_inst.timer_s1.counter_cry_22\,
            clk => \N__47247\,
            ce => \N__36410\,
            sr => \N__46648\
        );

    \current_shift_inst.timer_s1.counter_23_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36526\,
            in1 => \N__36693\,
            in2 => \_gnd_net_\,
            in3 => \N__36677\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_22\,
            carryout => \current_shift_inst.timer_s1.counter_cry_23\,
            clk => \N__47247\,
            ce => \N__36410\,
            sr => \N__46648\
        );

    \current_shift_inst.timer_s1.counter_24_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36527\,
            in1 => \N__36669\,
            in2 => \_gnd_net_\,
            in3 => \N__36650\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_15_16_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_24\,
            clk => \N__47240\,
            ce => \N__36408\,
            sr => \N__46658\
        );

    \current_shift_inst.timer_s1.counter_25_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36531\,
            in1 => \N__36642\,
            in2 => \_gnd_net_\,
            in3 => \N__36623\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_24\,
            carryout => \current_shift_inst.timer_s1.counter_cry_25\,
            clk => \N__47240\,
            ce => \N__36408\,
            sr => \N__46658\
        );

    \current_shift_inst.timer_s1.counter_26_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36528\,
            in1 => \N__36612\,
            in2 => \_gnd_net_\,
            in3 => \N__36596\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_25\,
            carryout => \current_shift_inst.timer_s1.counter_cry_26\,
            clk => \N__47240\,
            ce => \N__36408\,
            sr => \N__46658\
        );

    \current_shift_inst.timer_s1.counter_27_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36532\,
            in1 => \N__36585\,
            in2 => \_gnd_net_\,
            in3 => \N__36569\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_26\,
            carryout => \current_shift_inst.timer_s1.counter_cry_27\,
            clk => \N__47240\,
            ce => \N__36408\,
            sr => \N__46658\
        );

    \current_shift_inst.timer_s1.counter_28_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36529\,
            in1 => \N__36565\,
            in2 => \_gnd_net_\,
            in3 => \N__36551\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_27\,
            carryout => \current_shift_inst.timer_s1.counter_cry_28\,
            clk => \N__47240\,
            ce => \N__36408\,
            sr => \N__46658\
        );

    \current_shift_inst.timer_s1.counter_29_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__36424\,
            in1 => \N__36530\,
            in2 => \_gnd_net_\,
            in3 => \N__36428\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47240\,
            ce => \N__36408\,
            sr => \N__46658\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0_c_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36371\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_17_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36854\,
            in2 => \N__41210\,
            in3 => \N__38286\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36839\,
            in2 => \N__36848\,
            in3 => \N__38251\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__36826\,
            in1 => \N__36800\,
            in2 => \N__36809\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36785\,
            in2 => \N__36794\,
            in3 => \N__37597\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36779\,
            in2 => \N__43730\,
            in3 => \N__37564\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36764\,
            in2 => \N__36773\,
            in3 => \N__37486\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36731\,
            in2 => \N__36758\,
            in3 => \N__36742\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__36718\,
            in1 => \N__36707\,
            in2 => \N__40466\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \bfn_15_18_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37034\,
            in2 => \N__37028\,
            in3 => \N__38510\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37732\,
            in1 => \N__37004\,
            in2 => \N__37019\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36986\,
            in2 => \N__36998\,
            in3 => \N__37706\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36947\,
            in2 => \N__36980\,
            in3 => \N__36968\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36920\,
            in2 => \N__44225\,
            in3 => \N__36941\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36881\,
            in2 => \N__36914\,
            in3 => \N__36899\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36860\,
            in2 => \N__36875\,
            in3 => \N__38477\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37160\,
            in2 => \N__40409\,
            in3 => \N__37181\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \bfn_15_19_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37136\,
            in2 => \N__40475\,
            in3 => \N__37154\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40400\,
            in2 => \N__37112\,
            in3 => \N__37130\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37103\,
            in1 => \N__37085\,
            in2 => \N__40355\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37079\,
            lcout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_2_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__41437\,
            in1 => \N__37275\,
            in2 => \_gnd_net_\,
            in3 => \N__37361\,
            lcout => \phase_controller_inst1.stoper_tr.N_20_li\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__37075\,
            in1 => \N__38287\,
            in2 => \_gnd_net_\,
            in3 => \N__40718\,
            lcout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_2_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010001000000000"
        )
    port map (
            in0 => \N__40093\,
            in1 => \N__37437\,
            in2 => \N__40215\,
            in3 => \N__37455\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47218\,
            ce => \N__46827\,
            sr => \N__46690\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2_1_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40205\,
            in2 => \_gnd_net_\,
            in3 => \N__40092\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_1_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__40117\,
            in1 => \N__37438\,
            in2 => \N__37469\,
            in3 => \N__37454\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47218\,
            ce => \N__46827\,
            sr => \N__46690\
        );

    \phase_controller_inst1.stoper_tr.target_time_3_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__37456\,
            in1 => \N__40206\,
            in2 => \_gnd_net_\,
            in3 => \N__37439\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47218\,
            ce => \N__46827\,
            sr => \N__46690\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__37409\,
            in1 => \N__37385\,
            in2 => \_gnd_net_\,
            in3 => \N__39266\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_324_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_5_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__37279\,
            in1 => \N__41452\,
            in2 => \N__40177\,
            in3 => \N__37363\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47213\,
            ce => \N__46857\,
            sr => \N__46701\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001000101"
        )
    port map (
            in0 => \N__37364\,
            in1 => \N__40250\,
            in2 => \N__41480\,
            in3 => \N__37280\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47213\,
            ce => \N__46857\,
            sr => \N__46701\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__37278\,
            in1 => \N__43502\,
            in2 => \N__41479\,
            in3 => \N__37362\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47213\,
            ce => \N__46857\,
            sr => \N__46701\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__41451\,
            in1 => \N__37327\,
            in2 => \_gnd_net_\,
            in3 => \N__37276\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47213\,
            ce => \N__46857\,
            sr => \N__46701\
        );

    \phase_controller_inst1.stoper_tr.target_time_8_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__37277\,
            in1 => \N__41453\,
            in2 => \_gnd_net_\,
            in3 => \N__37225\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47213\,
            ce => \N__46857\,
            sr => \N__46701\
        );

    \phase_controller_inst1.stoper_tr.target_time_14_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__41447\,
            in1 => \N__47539\,
            in2 => \_gnd_net_\,
            in3 => \N__47706\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47213\,
            ce => \N__46857\,
            sr => \N__46701\
        );

    \phase_controller_inst1.stoper_tr.target_time_17_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43298\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47213\,
            ce => \N__46857\,
            sr => \N__46701\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_15_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__37885\,
            in1 => \N__38162\,
            in2 => \N__38044\,
            in3 => \N__37685\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47210\,
            ce => 'H',
            sr => \N__46708\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_12_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__37884\,
            in1 => \N__38161\,
            in2 => \N__38043\,
            in3 => \N__37661\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47210\,
            ce => 'H',
            sr => \N__46708\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_16_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__38160\,
            in1 => \N__38005\,
            in2 => \N__37901\,
            in3 => \N__37637\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47210\,
            ce => 'H',
            sr => \N__46708\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_4_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__41054\,
            in1 => \N__40630\,
            in2 => \N__40902\,
            in3 => \N__37613\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47210\,
            ce => 'H',
            sr => \N__46708\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_5_LC_15_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__40629\,
            in1 => \N__40872\,
            in2 => \N__41069\,
            in3 => \N__37580\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47210\,
            ce => 'H',
            sr => \N__46708\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_13_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__38159\,
            in1 => \N__38004\,
            in2 => \N__37900\,
            in3 => \N__37547\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47210\,
            ce => 'H',
            sr => \N__46708\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_9_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__37895\,
            in1 => \N__38178\,
            in2 => \N__38050\,
            in3 => \N__37523\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47207\,
            ce => 'H',
            sr => \N__46712\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_6_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__40632\,
            in1 => \N__40895\,
            in2 => \N__37499\,
            in3 => \N__41061\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47207\,
            ce => 'H',
            sr => \N__46712\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_14_LC_15_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__37893\,
            in1 => \N__38176\,
            in2 => \N__38048\,
            in3 => \N__38330\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47207\,
            ce => 'H',
            sr => \N__46712\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_1_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__40631\,
            in1 => \N__40894\,
            in2 => \N__38306\,
            in3 => \N__41060\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47207\,
            ce => 'H',
            sr => \N__46712\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_2_LC_15_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__41059\,
            in1 => \N__40633\,
            in2 => \N__40915\,
            in3 => \N__38264\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47207\,
            ce => 'H',
            sr => \N__46712\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_17_LC_15_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__38174\,
            in1 => \N__38037\,
            in2 => \N__38234\,
            in3 => \N__37896\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47207\,
            ce => 'H',
            sr => \N__46712\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_18_LC_15_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__37894\,
            in1 => \N__38177\,
            in2 => \N__38049\,
            in3 => \N__38204\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47207\,
            ce => 'H',
            sr => \N__46712\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_19_LC_15_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__38175\,
            in1 => \N__38038\,
            in2 => \N__37910\,
            in3 => \N__37897\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47207\,
            ce => 'H',
            sr => \N__46712\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_10_LC_15_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__41062\,
            in1 => \N__40635\,
            in2 => \N__40900\,
            in3 => \N__37742\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47203\,
            ce => 'H',
            sr => \N__46718\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_11_LC_15_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010100010"
        )
    port map (
            in0 => \N__37715\,
            in1 => \N__40861\,
            in2 => \N__40665\,
            in3 => \N__41065\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47203\,
            ce => 'H',
            sr => \N__46718\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_9_LC_15_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__41063\,
            in1 => \N__40636\,
            in2 => \N__40901\,
            in3 => \N__38519\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47203\,
            ce => 'H',
            sr => \N__46718\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_15_LC_15_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__40634\,
            in1 => \N__40862\,
            in2 => \N__38489\,
            in3 => \N__41064\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47203\,
            ce => 'H',
            sr => \N__46718\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_3_LC_16_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41824\,
            in2 => \_gnd_net_\,
            in3 => \N__41836\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.counter_0_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39031\,
            in1 => \N__38454\,
            in2 => \_gnd_net_\,
            in3 => \N__38438\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_16_7_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            clk => \N__47328\,
            ce => \N__38909\,
            sr => \N__46598\
        );

    \delay_measurement_inst.delay_hc_timer.counter_1_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39049\,
            in1 => \N__38433\,
            in2 => \_gnd_net_\,
            in3 => \N__38417\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            clk => \N__47328\,
            ce => \N__38909\,
            sr => \N__46598\
        );

    \delay_measurement_inst.delay_hc_timer.counter_2_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39032\,
            in1 => \N__38412\,
            in2 => \_gnd_net_\,
            in3 => \N__38393\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            clk => \N__47328\,
            ce => \N__38909\,
            sr => \N__46598\
        );

    \delay_measurement_inst.delay_hc_timer.counter_3_LC_16_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39050\,
            in1 => \N__38388\,
            in2 => \_gnd_net_\,
            in3 => \N__38369\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            clk => \N__47328\,
            ce => \N__38909\,
            sr => \N__46598\
        );

    \delay_measurement_inst.delay_hc_timer.counter_4_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39033\,
            in1 => \N__38366\,
            in2 => \_gnd_net_\,
            in3 => \N__38351\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            clk => \N__47328\,
            ce => \N__38909\,
            sr => \N__46598\
        );

    \delay_measurement_inst.delay_hc_timer.counter_5_LC_16_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39051\,
            in1 => \N__38348\,
            in2 => \_gnd_net_\,
            in3 => \N__38333\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            clk => \N__47328\,
            ce => \N__38909\,
            sr => \N__46598\
        );

    \delay_measurement_inst.delay_hc_timer.counter_6_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39034\,
            in1 => \N__38697\,
            in2 => \_gnd_net_\,
            in3 => \N__38678\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            clk => \N__47328\,
            ce => \N__38909\,
            sr => \N__46598\
        );

    \delay_measurement_inst.delay_hc_timer.counter_7_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39052\,
            in1 => \N__38673\,
            in2 => \_gnd_net_\,
            in3 => \N__38654\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            clk => \N__47328\,
            ce => \N__38909\,
            sr => \N__46598\
        );

    \delay_measurement_inst.delay_hc_timer.counter_8_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39056\,
            in1 => \N__38649\,
            in2 => \_gnd_net_\,
            in3 => \N__38630\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_16_8_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            clk => \N__47320\,
            ce => \N__38916\,
            sr => \N__46601\
        );

    \delay_measurement_inst.delay_hc_timer.counter_9_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39070\,
            in1 => \N__38625\,
            in2 => \_gnd_net_\,
            in3 => \N__38606\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            clk => \N__47320\,
            ce => \N__38916\,
            sr => \N__46601\
        );

    \delay_measurement_inst.delay_hc_timer.counter_10_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39053\,
            in1 => \N__38601\,
            in2 => \_gnd_net_\,
            in3 => \N__38582\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            clk => \N__47320\,
            ce => \N__38916\,
            sr => \N__46601\
        );

    \delay_measurement_inst.delay_hc_timer.counter_11_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39071\,
            in1 => \N__38577\,
            in2 => \_gnd_net_\,
            in3 => \N__38558\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            clk => \N__47320\,
            ce => \N__38916\,
            sr => \N__46601\
        );

    \delay_measurement_inst.delay_hc_timer.counter_12_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39054\,
            in1 => \N__38555\,
            in2 => \_gnd_net_\,
            in3 => \N__38540\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            clk => \N__47320\,
            ce => \N__38916\,
            sr => \N__46601\
        );

    \delay_measurement_inst.delay_hc_timer.counter_13_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39072\,
            in1 => \N__38537\,
            in2 => \_gnd_net_\,
            in3 => \N__38522\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            clk => \N__47320\,
            ce => \N__38916\,
            sr => \N__46601\
        );

    \delay_measurement_inst.delay_hc_timer.counter_14_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39055\,
            in1 => \N__38877\,
            in2 => \_gnd_net_\,
            in3 => \N__38858\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            clk => \N__47320\,
            ce => \N__38916\,
            sr => \N__46601\
        );

    \delay_measurement_inst.delay_hc_timer.counter_15_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39069\,
            in1 => \N__38853\,
            in2 => \_gnd_net_\,
            in3 => \N__38834\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            clk => \N__47320\,
            ce => \N__38916\,
            sr => \N__46601\
        );

    \delay_measurement_inst.delay_hc_timer.counter_16_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39057\,
            in1 => \N__38829\,
            in2 => \_gnd_net_\,
            in3 => \N__38810\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_16_9_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            clk => \N__47312\,
            ce => \N__38917\,
            sr => \N__46606\
        );

    \delay_measurement_inst.delay_hc_timer.counter_17_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39061\,
            in1 => \N__38805\,
            in2 => \_gnd_net_\,
            in3 => \N__38786\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            clk => \N__47312\,
            ce => \N__38917\,
            sr => \N__46606\
        );

    \delay_measurement_inst.delay_hc_timer.counter_18_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39058\,
            in1 => \N__38781\,
            in2 => \_gnd_net_\,
            in3 => \N__38762\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            clk => \N__47312\,
            ce => \N__38917\,
            sr => \N__46606\
        );

    \delay_measurement_inst.delay_hc_timer.counter_19_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39062\,
            in1 => \N__38757\,
            in2 => \_gnd_net_\,
            in3 => \N__38738\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            clk => \N__47312\,
            ce => \N__38917\,
            sr => \N__46606\
        );

    \delay_measurement_inst.delay_hc_timer.counter_20_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39059\,
            in1 => \N__38735\,
            in2 => \_gnd_net_\,
            in3 => \N__38720\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            clk => \N__47312\,
            ce => \N__38917\,
            sr => \N__46606\
        );

    \delay_measurement_inst.delay_hc_timer.counter_21_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39063\,
            in1 => \N__38717\,
            in2 => \_gnd_net_\,
            in3 => \N__38702\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            clk => \N__47312\,
            ce => \N__38917\,
            sr => \N__46606\
        );

    \delay_measurement_inst.delay_hc_timer.counter_22_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39060\,
            in1 => \N__39231\,
            in2 => \_gnd_net_\,
            in3 => \N__39212\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            clk => \N__47312\,
            ce => \N__38917\,
            sr => \N__46606\
        );

    \delay_measurement_inst.delay_hc_timer.counter_23_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39064\,
            in1 => \N__39207\,
            in2 => \_gnd_net_\,
            in3 => \N__39188\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            clk => \N__47312\,
            ce => \N__38917\,
            sr => \N__46606\
        );

    \delay_measurement_inst.delay_hc_timer.counter_24_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39065\,
            in1 => \N__39183\,
            in2 => \_gnd_net_\,
            in3 => \N__39164\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_16_10_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            clk => \N__47300\,
            ce => \N__38924\,
            sr => \N__46611\
        );

    \delay_measurement_inst.delay_hc_timer.counter_25_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39073\,
            in1 => \N__39159\,
            in2 => \_gnd_net_\,
            in3 => \N__39140\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            clk => \N__47300\,
            ce => \N__38924\,
            sr => \N__46611\
        );

    \delay_measurement_inst.delay_hc_timer.counter_26_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39066\,
            in1 => \N__39135\,
            in2 => \_gnd_net_\,
            in3 => \N__39116\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            clk => \N__47300\,
            ce => \N__38924\,
            sr => \N__46611\
        );

    \delay_measurement_inst.delay_hc_timer.counter_27_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39074\,
            in1 => \N__39111\,
            in2 => \_gnd_net_\,
            in3 => \N__39092\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            clk => \N__47300\,
            ce => \N__38924\,
            sr => \N__46611\
        );

    \delay_measurement_inst.delay_hc_timer.counter_28_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39067\,
            in1 => \N__39089\,
            in2 => \_gnd_net_\,
            in3 => \N__39077\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_28\,
            clk => \N__47300\,
            ce => \N__38924\,
            sr => \N__46611\
        );

    \delay_measurement_inst.delay_hc_timer.counter_29_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__38936\,
            in1 => \N__39068\,
            in2 => \_gnd_net_\,
            in3 => \N__38939\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47300\,
            ce => \N__38924\,
            sr => \N__46611\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43423\,
            lcout => \delay_measurement_inst.elapsed_time_tr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47291\,
            ce => \N__45718\,
            sr => \N__46615\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_9_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__42319\,
            in1 => \N__39401\,
            in2 => \N__42182\,
            in3 => \N__39351\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5PP_2_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__42796\,
            in1 => \N__47781\,
            in2 => \N__43402\,
            in3 => \N__44870\,
            lcout => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI200N_7_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__44662\,
            in1 => \N__44716\,
            in2 => \_gnd_net_\,
            in3 => \N__39446\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC3FA_2_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__39293\,
            in1 => \N__42770\,
            in2 => \N__39287\,
            in3 => \N__43523\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.N_375_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5KUTL_31_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__45802\,
            in1 => \N__39284\,
            in2 => \N__39272\,
            in3 => \N__39437\,
            lcout => \delay_measurement_inst.N_265_i\,
            ltout => \delay_measurement_inst.N_265_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICTS5M_31_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39269\,
            in3 => \N__46773\,
            lcout => \delay_measurement_inst.N_265_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39259\,
            lcout => \delay_measurement_inst.delay_tr_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4T357_15_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__45153\,
            in1 => \N__39536\,
            in2 => \_gnd_net_\,
            in3 => \N__43239\,
            lcout => \delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI43GB_6_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__44761\,
            in1 => \N__44655\,
            in2 => \_gnd_net_\,
            in3 => \N__44715\,
            lcout => \delay_measurement_inst.N_410\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI9IAF_1_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__40138\,
            in1 => \N__44812\,
            in2 => \N__44601\,
            in3 => \N__44760\,
            lcout => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ5M42_2_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100000000"
        )
    port map (
            in0 => \N__42797\,
            in1 => \N__44594\,
            in2 => \N__43403\,
            in3 => \N__42806\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_2_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__39431\,
            in1 => \N__43619\,
            in2 => \N__39440\,
            in3 => \N__39413\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_364\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI86841_4_LC_16_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__47780\,
            in1 => \N__44811\,
            in2 => \N__45160\,
            in3 => \N__44866\,
            lcout => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL5GJ7_15_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000010"
        )
    port map (
            in0 => \N__45155\,
            in1 => \N__42768\,
            in2 => \N__45801\,
            in3 => \N__43240\,
            lcout => \delay_measurement_inst.N_271_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO4MS_29_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45821\,
            in2 => \_gnd_net_\,
            in3 => \N__45875\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__45317\,
            in1 => \N__45356\,
            in2 => \N__45935\,
            in3 => \N__45392\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_6_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__45563\,
            in1 => \N__42812\,
            in2 => \N__39425\,
            in3 => \N__39422\,
            lcout => \delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20\,
            ltout => \delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI9DQM6_10_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39416\,
            in3 => \N__39535\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_409\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__45277\,
            in1 => \N__44488\,
            in2 => \N__45235\,
            in3 => \N__44542\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10\,
            ltout => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010001"
        )
    port map (
            in0 => \N__45154\,
            in1 => \N__47782\,
            in2 => \N__39524\,
            in3 => \N__44602\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.N_400_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111011100"
        )
    port map (
            in0 => \N__43241\,
            in1 => \N__45790\,
            in2 => \N__39521\,
            in3 => \N__42764\,
            lcout => \delay_measurement_inst.N_358\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_esr_9_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001101"
        )
    port map (
            in0 => \N__39515\,
            in1 => \N__44603\,
            in2 => \N__45803\,
            in3 => \N__43541\,
            lcout => measured_delay_tr_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47257\,
            ce => \N__43462\,
            sr => \N__46643\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110001"
        )
    port map (
            in0 => \N__47783\,
            in1 => \N__45161\,
            in2 => \N__42769\,
            in3 => \N__43242\,
            lcout => \delay_measurement_inst.N_394_1\,
            ltout => \delay_measurement_inst.N_394_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_esr_10_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45796\,
            in2 => \N__39518\,
            in3 => \N__44543\,
            lcout => measured_delay_tr_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47257\,
            ce => \N__43462\,
            sr => \N__46643\
        );

    \delay_measurement_inst.delay_tr_reg_esr_11_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__45794\,
            in1 => \N__39512\,
            in2 => \_gnd_net_\,
            in3 => \N__44492\,
            lcout => measured_delay_tr_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47257\,
            ce => \N__43462\,
            sr => \N__46643\
        );

    \delay_measurement_inst.delay_tr_reg_esr_12_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__39513\,
            in1 => \N__45797\,
            in2 => \_gnd_net_\,
            in3 => \N__45281\,
            lcout => measured_delay_tr_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47257\,
            ce => \N__43462\,
            sr => \N__46643\
        );

    \delay_measurement_inst.delay_tr_reg_esr_13_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__45795\,
            in1 => \N__39514\,
            in2 => \_gnd_net_\,
            in3 => \N__45236\,
            lcout => measured_delay_tr_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47257\,
            ce => \N__43462\,
            sr => \N__46643\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0_6_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__39489\,
            in1 => \N__41520\,
            in2 => \N__41991\,
            in3 => \N__39462\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_esr_6_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111100010011"
        )
    port map (
            in0 => \N__43544\,
            in1 => \N__43592\,
            in2 => \N__43648\,
            in3 => \N__44765\,
            lcout => measured_delay_tr_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47248\,
            ce => \N__43461\,
            sr => \N__46649\
        );

    \delay_measurement_inst.delay_tr_reg_ess_3_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010100010100000"
        )
    port map (
            in0 => \N__43401\,
            in1 => \N__43645\,
            in2 => \N__43602\,
            in3 => \N__43546\,
            lcout => measured_delay_tr_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47248\,
            ce => \N__43461\,
            sr => \N__46649\
        );

    \delay_measurement_inst.delay_tr_reg_esr_5_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010000000"
        )
    port map (
            in0 => \N__43543\,
            in1 => \N__43646\,
            in2 => \N__44819\,
            in3 => \N__43591\,
            lcout => measured_delay_tr_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47248\,
            ce => \N__43461\,
            sr => \N__46649\
        );

    \delay_measurement_inst.delay_tr_reg_esr_19_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__45785\,
            in1 => \N__44930\,
            in2 => \_gnd_net_\,
            in3 => \N__43253\,
            lcout => measured_delay_tr_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47248\,
            ce => \N__43461\,
            sr => \N__46649\
        );

    \delay_measurement_inst.delay_tr_reg_ess_1_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__43545\,
            in1 => \N__43593\,
            in2 => \N__43649\,
            in3 => \N__40139\,
            lcout => measured_delay_tr_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47248\,
            ce => \N__43461\,
            sr => \N__46649\
        );

    \delay_measurement_inst.delay_tr_reg_esr_2_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100010100000"
        )
    port map (
            in0 => \N__42789\,
            in1 => \N__43638\,
            in2 => \N__43601\,
            in3 => \N__43542\,
            lcout => measured_delay_tr_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47248\,
            ce => \N__43461\,
            sr => \N__46649\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_0_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__39568\,
            in1 => \N__39719\,
            in2 => \N__40019\,
            in3 => \N__40065\,
            lcout => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47241\,
            ce => \N__40518\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_1_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001010000"
        )
    port map (
            in0 => \N__40066\,
            in1 => \N__40011\,
            in2 => \N__39738\,
            in3 => \N__39569\,
            lcout => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47241\,
            ce => \N__40518\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_0_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__48028\,
            in1 => \N__48155\,
            in2 => \N__43344\,
            in3 => \N__47894\,
            lcout => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47241\,
            ce => \N__40518\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_1_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000110000"
        )
    port map (
            in0 => \N__48156\,
            in1 => \N__43334\,
            in2 => \N__47913\,
            in3 => \N__48029\,
            lcout => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47241\,
            ce => \N__40518\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__43333\,
            in1 => \N__43362\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.stoper_state_0_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__41021\,
            in1 => \N__40579\,
            in2 => \N__40919\,
            in3 => \N__40728\,
            lcout => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47241\,
            ce => \N__40518\,
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.target_time_17_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__44181\,
            in1 => \N__42347\,
            in2 => \_gnd_net_\,
            in3 => \N__43893\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47232\,
            ce => \N__43707\,
            sr => \N__46667\
        );

    \phase_controller_slave.stoper_hc.target_time_8_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__43896\,
            in1 => \N__44184\,
            in2 => \_gnd_net_\,
            in3 => \N__41767\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47232\,
            ce => \N__43707\,
            sr => \N__46667\
        );

    \phase_controller_slave.stoper_hc.target_time_16_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__44180\,
            in1 => \N__40454\,
            in2 => \_gnd_net_\,
            in3 => \N__43892\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47232\,
            ce => \N__43707\,
            sr => \N__46667\
        );

    \phase_controller_slave.stoper_hc.target_time_18_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__43894\,
            in1 => \N__44182\,
            in2 => \_gnd_net_\,
            in3 => \N__42190\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47232\,
            ce => \N__43707\,
            sr => \N__46667\
        );

    \phase_controller_slave.stoper_hc.target_time_19_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__44179\,
            in1 => \N__40394\,
            in2 => \_gnd_net_\,
            in3 => \N__41888\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47232\,
            ce => \N__43707\,
            sr => \N__46667\
        );

    \phase_controller_slave.stoper_hc.target_time_1_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110101000"
        )
    port map (
            in0 => \N__43895\,
            in1 => \N__40342\,
            in2 => \N__41275\,
            in3 => \N__44183\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47232\,
            ce => \N__43707\,
            sr => \N__46667\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41192\,
            in2 => \N__41201\,
            in3 => \N__45660\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_16_19_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41186\,
            in2 => \N__41180\,
            in3 => \N__45643\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41156\,
            in2 => \N__41171\,
            in3 => \N__45610\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41138\,
            in2 => \N__41150\,
            in3 => \N__46111\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41117\,
            in2 => \N__41132\,
            in3 => \N__46090\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41096\,
            in2 => \N__41111\,
            in3 => \N__46069\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__46048\,
            in1 => \N__41075\,
            in2 => \N__41090\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__46027\,
            in1 => \N__41369\,
            in2 => \N__41381\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41363\,
            in2 => \N__47363\,
            in3 => \N__48214\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_16_20_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__46003\,
            in1 => \N__41339\,
            in2 => \N__41357\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41333\,
            in2 => \N__41504\,
            in3 => \N__45982\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41309\,
            in2 => \N__41327\,
            in3 => \N__46291\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41303\,
            in2 => \N__41966\,
            in3 => \N__46270\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41288\,
            in2 => \N__41297\,
            in3 => \N__46249\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__46225\,
            in1 => \N__41282\,
            in2 => \N__41393\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41624\,
            in2 => \N__44357\,
            in3 => \N__46202\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_16_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41606\,
            in2 => \N__41618\,
            in3 => \N__46177\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_16_21_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41600\,
            in2 => \N__41585\,
            in3 => \N__46156\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41594\,
            in2 => \N__41540\,
            in3 => \N__46135\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41588\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_18_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43210\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47219\,
            ce => \N__46856\,
            sr => \N__46691\
        );

    \phase_controller_inst1.stoper_tr.target_time_19_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41567\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47219\,
            ce => \N__46856\,
            sr => \N__46691\
        );

    \phase_controller_inst1.stoper_tr.target_time_11_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47593\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41527\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47214\,
            ce => \N__46859\,
            sr => \N__46702\
        );

    \phase_controller_inst1.stoper_tr.target_time_15_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41491\,
            in2 => \_gnd_net_\,
            in3 => \N__47538\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47214\,
            ce => \N__46859\,
            sr => \N__46702\
        );

    \phase_controller_inst1.stoper_tr.target_time_13_LC_16_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47594\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41998\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47214\,
            ce => \N__46859\,
            sr => \N__46702\
        );

    \SB_DFF_inst_DELAY_HC1_LC_17_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41954\,
            lcout => delay_hc_d1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_DELAY_HC2_LC_17_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41945\,
            lcout => delay_hc_d2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_LC_17_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__41809\,
            in1 => \N__44291\,
            in2 => \N__42275\,
            in3 => \N__41894\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_25_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__42466\,
            in1 => \N__41837\,
            in2 => \_gnd_net_\,
            in3 => \N__42559\,
            lcout => measured_delay_hc_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47335\,
            ce => 'H',
            sr => \N__46595\
        );

    \delay_measurement_inst.delay_hc_reg_26_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__42560\,
            in1 => \N__41825\,
            in2 => \_gnd_net_\,
            in3 => \N__42467\,
            lcout => measured_delay_hc_26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47335\,
            ce => 'H',
            sr => \N__46595\
        );

    \delay_measurement_inst.delay_hc_reg_23_LC_17_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__42465\,
            in1 => \_gnd_net_\,
            in2 => \N__41813\,
            in3 => \N__42558\,
            lcout => measured_delay_hc_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47335\,
            ce => 'H',
            sr => \N__46595\
        );

    \delay_measurement_inst.delay_hc_reg_8_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__42104\,
            in1 => \N__41740\,
            in2 => \N__42651\,
            in3 => \N__41801\,
            lcout => measured_delay_hc_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47329\,
            ce => 'H',
            sr => \N__46599\
        );

    \delay_measurement_inst.delay_hc_reg_7_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__41648\,
            in1 => \N__42632\,
            in2 => \N__41708\,
            in3 => \N__42103\,
            lcout => measured_delay_hc_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47329\,
            ce => 'H',
            sr => \N__46599\
        );

    \delay_measurement_inst.delay_hc_reg_24_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__42446\,
            in1 => \N__42274\,
            in2 => \_gnd_net_\,
            in3 => \N__42630\,
            lcout => measured_delay_hc_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47329\,
            ce => 'H',
            sr => \N__46599\
        );

    \delay_measurement_inst.delay_hc_reg_0_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__42629\,
            in1 => \N__42233\,
            in2 => \_gnd_net_\,
            in3 => \N__42444\,
            lcout => measured_delay_hc_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47329\,
            ce => 'H',
            sr => \N__46599\
        );

    \delay_measurement_inst.delay_hc_reg_18_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111010111010"
        )
    port map (
            in0 => \N__42445\,
            in1 => \N__42631\,
            in2 => \N__42181\,
            in3 => \N__42209\,
            lcout => measured_delay_hc_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47329\,
            ce => 'H',
            sr => \N__46599\
        );

    \delay_measurement_inst.delay_hc_reg_30_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__42441\,
            in1 => \_gnd_net_\,
            in2 => \N__42653\,
            in3 => \N__44317\,
            lcout => measured_delay_hc_30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47321\,
            ce => 'H',
            sr => \N__46602\
        );

    \delay_measurement_inst.delay_hc_reg_29_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__44342\,
            in1 => \N__42640\,
            in2 => \_gnd_net_\,
            in3 => \N__42440\,
            lcout => measured_delay_hc_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47321\,
            ce => 'H',
            sr => \N__46602\
        );

    \delay_measurement_inst.delay_hc_reg_19_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011111111"
        )
    port map (
            in0 => \N__42048\,
            in1 => \N__42644\,
            in2 => \N__42134\,
            in3 => \N__42093\,
            lcout => measured_delay_hc_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47321\,
            ce => 'H',
            sr => \N__46602\
        );

    \delay_measurement_inst.delay_hc_reg_28_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__42439\,
            in1 => \_gnd_net_\,
            in2 => \N__42652\,
            in3 => \N__44330\,
            lcout => measured_delay_hc_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47321\,
            ce => 'H',
            sr => \N__46602\
        );

    \delay_measurement_inst.delay_hc_reg_27_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__44303\,
            in1 => \N__42636\,
            in2 => \_gnd_net_\,
            in3 => \N__42438\,
            lcout => measured_delay_hc_27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47321\,
            ce => 'H',
            sr => \N__46602\
        );

    \delay_measurement_inst.delay_hc_reg_21_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__42013\,
            in1 => \N__42645\,
            in2 => \_gnd_net_\,
            in3 => \N__42463\,
            lcout => measured_delay_hc_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47313\,
            ce => 'H',
            sr => \N__46607\
        );

    \delay_measurement_inst.delay_hc_reg_22_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__42667\,
            in1 => \N__42646\,
            in2 => \_gnd_net_\,
            in3 => \N__42464\,
            lcout => measured_delay_hc_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47313\,
            ce => 'H',
            sr => \N__46607\
        );

    \delay_measurement_inst.delay_hc_reg_17_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111100010"
        )
    port map (
            in0 => \N__42329\,
            in1 => \N__42647\,
            in2 => \N__42491\,
            in3 => \N__42462\,
            lcout => measured_delay_hc_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47313\,
            ce => 'H',
            sr => \N__46607\
        );

    \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42980\,
            in1 => \N__43419\,
            in2 => \_gnd_net_\,
            in3 => \N__42296\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_17_11_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            clk => \N__47301\,
            ce => \N__42857\,
            sr => \N__46612\
        );

    \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42961\,
            in1 => \N__44889\,
            in2 => \_gnd_net_\,
            in3 => \N__42293\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            clk => \N__47301\,
            ce => \N__42857\,
            sr => \N__46612\
        );

    \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42981\,
            in1 => \N__44835\,
            in2 => \_gnd_net_\,
            in3 => \N__42290\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            clk => \N__47301\,
            ce => \N__42857\,
            sr => \N__46612\
        );

    \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42962\,
            in1 => \N__44781\,
            in2 => \_gnd_net_\,
            in3 => \N__42287\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            clk => \N__47301\,
            ce => \N__42857\,
            sr => \N__46612\
        );

    \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42982\,
            in1 => \N__44731\,
            in2 => \_gnd_net_\,
            in3 => \N__42284\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            clk => \N__47301\,
            ce => \N__42857\,
            sr => \N__46612\
        );

    \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42963\,
            in1 => \N__44677\,
            in2 => \_gnd_net_\,
            in3 => \N__42281\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            clk => \N__47301\,
            ce => \N__42857\,
            sr => \N__46612\
        );

    \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42983\,
            in1 => \N__44625\,
            in2 => \_gnd_net_\,
            in3 => \N__42278\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            clk => \N__47301\,
            ce => \N__42857\,
            sr => \N__46612\
        );

    \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42964\,
            in1 => \N__44557\,
            in2 => \_gnd_net_\,
            in3 => \N__42710\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            clk => \N__47301\,
            ce => \N__42857\,
            sr => \N__46612\
        );

    \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42956\,
            in1 => \N__44511\,
            in2 => \_gnd_net_\,
            in3 => \N__42707\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_17_12_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            clk => \N__47292\,
            ce => \N__42856\,
            sr => \N__46616\
        );

    \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42968\,
            in1 => \N__45298\,
            in2 => \_gnd_net_\,
            in3 => \N__42704\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            clk => \N__47292\,
            ce => \N__42856\,
            sr => \N__46616\
        );

    \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42953\,
            in1 => \N__45252\,
            in2 => \_gnd_net_\,
            in3 => \N__42701\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            clk => \N__47292\,
            ce => \N__42856\,
            sr => \N__46616\
        );

    \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42965\,
            in1 => \N__45201\,
            in2 => \_gnd_net_\,
            in3 => \N__42698\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            clk => \N__47292\,
            ce => \N__42856\,
            sr => \N__46616\
        );

    \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42954\,
            in1 => \N__45175\,
            in2 => \_gnd_net_\,
            in3 => \N__42695\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            clk => \N__47292\,
            ce => \N__42856\,
            sr => \N__46616\
        );

    \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42966\,
            in1 => \N__45094\,
            in2 => \_gnd_net_\,
            in3 => \N__42692\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            clk => \N__47292\,
            ce => \N__42856\,
            sr => \N__46616\
        );

    \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42955\,
            in1 => \N__45051\,
            in2 => \_gnd_net_\,
            in3 => \N__42689\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            clk => \N__47292\,
            ce => \N__42856\,
            sr => \N__46616\
        );

    \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42967\,
            in1 => \N__44992\,
            in2 => \_gnd_net_\,
            in3 => \N__42686\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            clk => \N__47292\,
            ce => \N__42856\,
            sr => \N__46616\
        );

    \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42945\,
            in1 => \N__44949\,
            in2 => \_gnd_net_\,
            in3 => \N__42737\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_17_13_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            clk => \N__47284\,
            ce => \N__42849\,
            sr => \N__46619\
        );

    \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42949\,
            in1 => \N__45583\,
            in2 => \_gnd_net_\,
            in3 => \N__42734\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            clk => \N__47284\,
            ce => \N__42849\,
            sr => \N__46619\
        );

    \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42946\,
            in1 => \N__45537\,
            in2 => \_gnd_net_\,
            in3 => \N__42731\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            clk => \N__47284\,
            ce => \N__42849\,
            sr => \N__46619\
        );

    \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42950\,
            in1 => \N__45504\,
            in2 => \_gnd_net_\,
            in3 => \N__42728\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            clk => \N__47284\,
            ce => \N__42849\,
            sr => \N__46619\
        );

    \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42947\,
            in1 => \N__45471\,
            in2 => \_gnd_net_\,
            in3 => \N__42725\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            clk => \N__47284\,
            ce => \N__42849\,
            sr => \N__46619\
        );

    \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42951\,
            in1 => \N__45438\,
            in2 => \_gnd_net_\,
            in3 => \N__42722\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            clk => \N__47284\,
            ce => \N__42849\,
            sr => \N__46619\
        );

    \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42948\,
            in1 => \N__45408\,
            in2 => \_gnd_net_\,
            in3 => \N__42719\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            clk => \N__47284\,
            ce => \N__42849\,
            sr => \N__46619\
        );

    \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42952\,
            in1 => \N__45370\,
            in2 => \_gnd_net_\,
            in3 => \N__42716\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            clk => \N__47284\,
            ce => \N__42849\,
            sr => \N__46619\
        );

    \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42957\,
            in1 => \N__45336\,
            in2 => \_gnd_net_\,
            in3 => \N__42713\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_17_14_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            clk => \N__47277\,
            ce => \N__42839\,
            sr => \N__46631\
        );

    \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42969\,
            in1 => \N__45954\,
            in2 => \_gnd_net_\,
            in3 => \N__42995\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            clk => \N__47277\,
            ce => \N__42839\,
            sr => \N__46631\
        );

    \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42958\,
            in1 => \N__45891\,
            in2 => \_gnd_net_\,
            in3 => \N__42992\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            clk => \N__47277\,
            ce => \N__42839\,
            sr => \N__46631\
        );

    \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42970\,
            in1 => \N__45837\,
            in2 => \_gnd_net_\,
            in3 => \N__42989\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            clk => \N__47277\,
            ce => \N__42839\,
            sr => \N__46631\
        );

    \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42959\,
            in1 => \N__45913\,
            in2 => \_gnd_net_\,
            in3 => \N__42986\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_28\,
            clk => \N__47277\,
            ce => \N__42839\,
            sr => \N__46631\
        );

    \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__45859\,
            in1 => \N__42960\,
            in2 => \_gnd_net_\,
            in3 => \N__42860\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47277\,
            ce => \N__42839\,
            sr => \N__46631\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__45455\,
            in1 => \N__45488\,
            in2 => \N__45422\,
            in3 => \N__45515\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_7_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_0_16_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__44973\,
            in1 => \N__45024\,
            in2 => \N__44925\,
            in3 => \N__45075\,
            lcout => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44897\,
            lcout => \delay_measurement_inst.elapsed_time_tr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47265\,
            ce => \N__45725\,
            sr => \N__46636\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__45076\,
            in1 => \N__44974\,
            in2 => \N__44926\,
            in3 => \N__45025\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_esr_16_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__45080\,
            in1 => \N__45760\,
            in2 => \_gnd_net_\,
            in3 => \N__43254\,
            lcout => measured_delay_tr_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47258\,
            ce => \N__43463\,
            sr => \N__46644\
        );

    \delay_measurement_inst.delay_tr_reg_esr_17_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100001010"
        )
    port map (
            in0 => \N__43255\,
            in1 => \_gnd_net_\,
            in2 => \N__45786\,
            in3 => \N__45029\,
            lcout => measured_delay_tr_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47258\,
            ce => \N__43463\,
            sr => \N__46644\
        );

    \delay_measurement_inst.delay_tr_reg_esr_18_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__44978\,
            in1 => \N__45761\,
            in2 => \_gnd_net_\,
            in3 => \N__43256\,
            lcout => measured_delay_tr_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47258\,
            ce => \N__43463\,
            sr => \N__46644\
        );

    \phase_controller_inst1.state_RNI7NN7_0_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43050\,
            in2 => \_gnd_net_\,
            in3 => \N__43003\,
            lcout => \phase_controller_inst1.N_83\,
            ltout => \phase_controller_inst1.N_83_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_tr_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000010"
        )
    port map (
            in0 => \N__48157\,
            in1 => \N__43160\,
            in2 => \N__43127\,
            in3 => \N__43124\,
            lcout => \phase_controller_inst1.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47249\,
            ce => 'H',
            sr => \N__46650\
        );

    \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__48158\,
            in1 => \N__47998\,
            in2 => \_gnd_net_\,
            in3 => \N__47873\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.time_passed_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__43054\,
            in1 => \N__43366\,
            in2 => \N__43103\,
            in3 => \N__43346\,
            lcout => \phase_controller_inst1.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47249\,
            ce => 'H',
            sr => \N__46650\
        );

    \phase_controller_inst1.state_0_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111000001010"
        )
    port map (
            in0 => \N__43004\,
            in1 => \N__43096\,
            in2 => \N__43055\,
            in3 => \N__43040\,
            lcout => \phase_controller_inst1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47249\,
            ce => 'H',
            sr => \N__46650\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47997\,
            in2 => \_gnd_net_\,
            in3 => \N__47872\,
            lcout => \phase_controller_inst1.stoper_tr.time_passed11\,
            ltout => \phase_controller_inst1.stoper_tr.time_passed11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43301\,
            in3 => \N__43345\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__47889\,
            in1 => \N__48154\,
            in2 => \N__48066\,
            in3 => \N__46016\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47242\,
            ce => 'H',
            sr => \N__46659\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__48024\,
            in1 => \N__47890\,
            in2 => \N__48179\,
            in3 => \N__46187\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47242\,
            ce => 'H',
            sr => \N__46659\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__47888\,
            in1 => \N__48153\,
            in2 => \N__48065\,
            in3 => \N__46037\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47242\,
            ce => 'H',
            sr => \N__46659\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__48025\,
            in1 => \N__47891\,
            in2 => \N__48180\,
            in3 => \N__45632\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47242\,
            ce => 'H',
            sr => \N__46659\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__47886\,
            in1 => \N__48145\,
            in2 => \N__48063\,
            in3 => \N__45599\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47242\,
            ce => 'H',
            sr => \N__46659\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__48026\,
            in1 => \N__47892\,
            in2 => \N__48181\,
            in3 => \N__46100\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47242\,
            ce => 'H',
            sr => \N__46659\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__47887\,
            in1 => \N__48149\,
            in2 => \N__48064\,
            in3 => \N__46079\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47242\,
            ce => 'H',
            sr => \N__46659\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__48027\,
            in1 => \N__47893\,
            in2 => \N__48182\,
            in3 => \N__46058\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47242\,
            ce => 'H',
            sr => \N__46659\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100010001100"
        )
    port map (
            in0 => \N__47910\,
            in1 => \N__45992\,
            in2 => \N__48071\,
            in3 => \N__48173\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47233\,
            ce => 'H',
            sr => \N__46668\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__43367\,
            in1 => \N__45664\,
            in2 => \_gnd_net_\,
            in3 => \N__43343\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011010000"
        )
    port map (
            in0 => \N__48047\,
            in1 => \N__47933\,
            in2 => \N__43304\,
            in3 => \N__48178\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47233\,
            ce => 'H',
            sr => \N__46668\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__48174\,
            in1 => \N__48048\,
            in2 => \N__47946\,
            in3 => \N__45971\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47233\,
            ce => 'H',
            sr => \N__46668\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__47911\,
            in1 => \N__48175\,
            in2 => \N__48072\,
            in3 => \N__46280\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47233\,
            ce => 'H',
            sr => \N__46668\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__48176\,
            in1 => \N__48049\,
            in2 => \N__47947\,
            in3 => \N__46259\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47233\,
            ce => 'H',
            sr => \N__46668\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__47912\,
            in1 => \N__48177\,
            in2 => \N__48073\,
            in3 => \N__46238\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47233\,
            ce => 'H',
            sr => \N__46668\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__48059\,
            in1 => \N__48185\,
            in2 => \N__47948\,
            in3 => \N__46214\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47227\,
            ce => 'H',
            sr => \N__46677\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__47942\,
            in1 => \N__48061\,
            in2 => \N__48197\,
            in3 => \N__46121\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47227\,
            ce => 'H',
            sr => \N__46677\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100010001100"
        )
    port map (
            in0 => \N__47940\,
            in1 => \N__46166\,
            in2 => \N__48195\,
            in3 => \N__48062\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47227\,
            ce => 'H',
            sr => \N__46677\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__47941\,
            in1 => \N__48060\,
            in2 => \N__48196\,
            in3 => \N__46145\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47227\,
            ce => 'H',
            sr => \N__46677\
        );

    \phase_controller_slave.stoper_tr.target_time_16_LC_17_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44384\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47224\,
            ce => \N__44453\,
            sr => \N__46682\
        );

    \phase_controller_inst1.stoper_tr.target_time_16_LC_17_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44385\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47220\,
            ce => \N__46852\,
            sr => \N__46692\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_4_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__44341\,
            in1 => \N__44329\,
            in2 => \N__44318\,
            in3 => \N__44302\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.target_time_13_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__44154\,
            in1 => \N__44282\,
            in2 => \_gnd_net_\,
            in3 => \N__43897\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47322\,
            ce => \N__43712\,
            sr => \N__46603\
        );

    \phase_controller_slave.stoper_hc.target_time_5_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__44156\,
            in1 => \N__43957\,
            in2 => \_gnd_net_\,
            in3 => \N__43827\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47314\,
            ce => \N__43711\,
            sr => \N__46608\
        );

    \delay_measurement_inst.delay_tr_reg_esr_4_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100010100000"
        )
    port map (
            in0 => \N__44865\,
            in1 => \N__43647\,
            in2 => \N__43604\,
            in3 => \N__43550\,
            lcout => measured_delay_tr_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47302\,
            ce => \N__43451\,
            sr => \N__46613\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43424\,
            in2 => \N__44842\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.elapsed_time_tr_3\,
            ltout => OPEN,
            carryin => \bfn_18_13_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__47293\,
            ce => \N__45703\,
            sr => \N__46617\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_18_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44893\,
            in2 => \N__44788\,
            in3 => \N__44846\,
            lcout => \delay_measurement_inst.elapsed_time_tr_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__47293\,
            ce => \N__45703\,
            sr => \N__46617\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44737\,
            in2 => \N__44843\,
            in3 => \N__44792\,
            lcout => \delay_measurement_inst.elapsed_time_tr_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__47293\,
            ce => \N__45703\,
            sr => \N__46617\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44683\,
            in2 => \N__44789\,
            in3 => \N__44741\,
            lcout => \delay_measurement_inst.elapsed_time_tr_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__47293\,
            ce => \N__45703\,
            sr => \N__46617\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44738\,
            in2 => \N__44633\,
            in3 => \N__44687\,
            lcout => \delay_measurement_inst.elapsed_time_tr_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__47293\,
            ce => \N__45703\,
            sr => \N__46617\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44684\,
            in2 => \N__44569\,
            in3 => \N__44636\,
            lcout => \delay_measurement_inst.elapsed_time_tr_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__47293\,
            ce => \N__45703\,
            sr => \N__46617\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_18_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44629\,
            in2 => \N__44515\,
            in3 => \N__44573\,
            lcout => \delay_measurement_inst.elapsed_time_tr_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__47293\,
            ce => \N__45703\,
            sr => \N__46617\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_18_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45297\,
            in2 => \N__44570\,
            in3 => \N__44519\,
            lcout => \delay_measurement_inst.elapsed_time_tr_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__47293\,
            ce => \N__45703\,
            sr => \N__46617\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44516\,
            in2 => \N__45259\,
            in3 => \N__44474\,
            lcout => \delay_measurement_inst.elapsed_time_tr_11\,
            ltout => OPEN,
            carryin => \bfn_18_14_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__47285\,
            ce => \N__45727\,
            sr => \N__46620\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45302\,
            in2 => \N__45208\,
            in3 => \N__45263\,
            lcout => \delay_measurement_inst.elapsed_time_tr_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__47285\,
            ce => \N__45727\,
            sr => \N__46620\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45181\,
            in2 => \N__45260\,
            in3 => \N__45212\,
            lcout => \delay_measurement_inst.elapsed_time_tr_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__47285\,
            ce => \N__45727\,
            sr => \N__46620\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45100\,
            in2 => \N__45209\,
            in3 => \N__45185\,
            lcout => \delay_measurement_inst.elapsed_time_tr_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__47285\,
            ce => \N__45727\,
            sr => \N__46620\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45182\,
            in2 => \N__45059\,
            in3 => \N__45104\,
            lcout => \delay_measurement_inst.elapsed_time_tr_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__47285\,
            ce => \N__45727\,
            sr => \N__46620\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45101\,
            in2 => \N__45004\,
            in3 => \N__45062\,
            lcout => \delay_measurement_inst.elapsed_time_tr_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__47285\,
            ce => \N__45727\,
            sr => \N__46620\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45055\,
            in2 => \N__44953\,
            in3 => \N__45008\,
            lcout => \delay_measurement_inst.elapsed_time_tr_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__47285\,
            ce => \N__45727\,
            sr => \N__46620\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_18_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45579\,
            in2 => \N__45005\,
            in3 => \N__44960\,
            lcout => \delay_measurement_inst.elapsed_time_tr_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__47285\,
            ce => \N__45727\,
            sr => \N__46620\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44957\,
            in2 => \N__45548\,
            in3 => \N__44900\,
            lcout => \delay_measurement_inst.elapsed_time_tr_19\,
            ltout => OPEN,
            carryin => \bfn_18_15_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__47278\,
            ce => \N__45726\,
            sr => \N__46632\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45505\,
            in2 => \N__45590\,
            in3 => \N__45551\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__47278\,
            ce => \N__45726\,
            sr => \N__46632\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45547\,
            in2 => \N__45478\,
            in3 => \N__45509\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__47278\,
            ce => \N__45726\,
            sr => \N__46632\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45506\,
            in2 => \N__45445\,
            in3 => \N__45482\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__47278\,
            ce => \N__45726\,
            sr => \N__46632\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45409\,
            in2 => \N__45479\,
            in3 => \N__45449\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__47278\,
            ce => \N__45726\,
            sr => \N__46632\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45376\,
            in2 => \N__45446\,
            in3 => \N__45413\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__47278\,
            ce => \N__45726\,
            sr => \N__46632\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45410\,
            in2 => \N__45340\,
            in3 => \N__45380\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__47278\,
            ce => \N__45726\,
            sr => \N__46632\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_18_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45377\,
            in2 => \N__45958\,
            in3 => \N__45344\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__47278\,
            ce => \N__45726\,
            sr => \N__46632\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45341\,
            in2 => \N__45898\,
            in3 => \N__45305\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\,
            ltout => OPEN,
            carryin => \bfn_18_16_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__47266\,
            ce => \N__45731\,
            sr => \N__46637\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45962\,
            in2 => \N__45844\,
            in3 => \N__45920\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__47266\,
            ce => \N__45731\,
            sr => \N__46637\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45917\,
            in2 => \N__45899\,
            in3 => \N__45863\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__47266\,
            ce => \N__45731\,
            sr => \N__46637\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45860\,
            in2 => \N__45845\,
            in3 => \N__45809\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__47266\,
            ce => \N__45731\,
            sr => \N__46637\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45806\,
            lcout => \delay_measurement_inst.elapsed_time_tr_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47266\,
            ce => \N__45731\,
            sr => \N__46637\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45674\,
            in2 => \N__45668\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_17_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45644\,
            in2 => \_gnd_net_\,
            in3 => \N__45626\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45623\,
            in2 => \N__45614\,
            in3 => \N__45593\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__46115\,
            in3 => \N__46094\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46091\,
            in2 => \_gnd_net_\,
            in3 => \N__46073\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46070\,
            in2 => \_gnd_net_\,
            in3 => \N__46052\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46049\,
            in2 => \_gnd_net_\,
            in3 => \N__46031\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_18_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46028\,
            in2 => \_gnd_net_\,
            in3 => \N__46010\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_18_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48215\,
            in2 => \_gnd_net_\,
            in3 => \N__46007\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9\,
            ltout => OPEN,
            carryin => \bfn_18_18_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46004\,
            in2 => \_gnd_net_\,
            in3 => \N__45986\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45983\,
            in2 => \_gnd_net_\,
            in3 => \N__45965\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_18_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46292\,
            in2 => \_gnd_net_\,
            in3 => \N__46274\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46271\,
            in2 => \_gnd_net_\,
            in3 => \N__46253\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46250\,
            in2 => \_gnd_net_\,
            in3 => \N__46232\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_18_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46229\,
            in2 => \_gnd_net_\,
            in3 => \N__46205\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46201\,
            in2 => \_gnd_net_\,
            in3 => \N__46181\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_18_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46178\,
            in2 => \_gnd_net_\,
            in3 => \N__46160\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17\,
            ltout => OPEN,
            carryin => \bfn_18_19_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46157\,
            in2 => \_gnd_net_\,
            in3 => \N__46139\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_18_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46136\,
            in2 => \_gnd_net_\,
            in3 => \N__46124\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__47915\,
            in1 => \N__48184\,
            in2 => \N__48074\,
            in3 => \N__48224\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47234\,
            ce => 'H',
            sr => \N__46669\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_18_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__48183\,
            in1 => \N__48067\,
            in2 => \_gnd_net_\,
            in3 => \N__47914\,
            lcout => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_0_13_LC_18_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47530\,
            in2 => \_gnd_net_\,
            in3 => \N__47684\,
            lcout => \phase_controller_inst1.stoper_tr.N_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_14_LC_18_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011110000"
        )
    port map (
            in0 => \N__47810\,
            in1 => \N__47779\,
            in2 => \N__47694\,
            in3 => \N__47735\,
            lcout => measured_delay_tr_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47234\,
            ce => 'H',
            sr => \N__46669\
        );

    \phase_controller_slave.start_timer_hc_RNO_0_LC_18_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47666\,
            in2 => \_gnd_net_\,
            in3 => \N__47642\,
            lcout => \phase_controller_slave.N_211\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_9_LC_20_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010011110101"
        )
    port map (
            in0 => \N__47604\,
            in1 => \N__47540\,
            in2 => \N__47447\,
            in3 => \N__47402\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47250\,
            ce => \N__46826\,
            sr => \N__46670\
        );
end \INTERFACE\;
