// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jul 10 2025 20:22:24

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "MAIN" view "INTERFACE"

module MAIN (
    s3_phy,
    il_min_comp2,
    il_max_comp1,
    s1_phy,
    reset,
    il_min_comp1,
    delay_tr_input,
    s4_phy,
    rgb_g,
    start_stop,
    s2_phy,
    rgb_r,
    rgb_b,
    pwm_output,
    il_max_comp2,
    delay_hc_input);

    output s3_phy;
    input il_min_comp2;
    input il_max_comp1;
    output s1_phy;
    input reset;
    input il_min_comp1;
    input delay_tr_input;
    output s4_phy;
    output rgb_g;
    input start_stop;
    output s2_phy;
    output rgb_r;
    output rgb_b;
    output pwm_output;
    input il_max_comp2;
    input delay_hc_input;

    wire N__50761;
    wire N__50760;
    wire N__50759;
    wire N__50750;
    wire N__50749;
    wire N__50748;
    wire N__50741;
    wire N__50740;
    wire N__50739;
    wire N__50732;
    wire N__50731;
    wire N__50730;
    wire N__50723;
    wire N__50722;
    wire N__50721;
    wire N__50714;
    wire N__50713;
    wire N__50712;
    wire N__50705;
    wire N__50704;
    wire N__50703;
    wire N__50696;
    wire N__50695;
    wire N__50694;
    wire N__50687;
    wire N__50686;
    wire N__50685;
    wire N__50678;
    wire N__50677;
    wire N__50676;
    wire N__50669;
    wire N__50668;
    wire N__50667;
    wire N__50660;
    wire N__50659;
    wire N__50658;
    wire N__50651;
    wire N__50650;
    wire N__50649;
    wire N__50632;
    wire N__50631;
    wire N__50628;
    wire N__50625;
    wire N__50624;
    wire N__50619;
    wire N__50616;
    wire N__50613;
    wire N__50608;
    wire N__50605;
    wire N__50604;
    wire N__50601;
    wire N__50598;
    wire N__50597;
    wire N__50592;
    wire N__50589;
    wire N__50586;
    wire N__50581;
    wire N__50578;
    wire N__50577;
    wire N__50574;
    wire N__50571;
    wire N__50570;
    wire N__50565;
    wire N__50562;
    wire N__50559;
    wire N__50554;
    wire N__50551;
    wire N__50550;
    wire N__50547;
    wire N__50544;
    wire N__50541;
    wire N__50536;
    wire N__50533;
    wire N__50532;
    wire N__50531;
    wire N__50530;
    wire N__50529;
    wire N__50528;
    wire N__50527;
    wire N__50526;
    wire N__50525;
    wire N__50524;
    wire N__50523;
    wire N__50522;
    wire N__50521;
    wire N__50520;
    wire N__50519;
    wire N__50518;
    wire N__50517;
    wire N__50516;
    wire N__50515;
    wire N__50514;
    wire N__50513;
    wire N__50512;
    wire N__50511;
    wire N__50510;
    wire N__50509;
    wire N__50508;
    wire N__50507;
    wire N__50506;
    wire N__50505;
    wire N__50504;
    wire N__50499;
    wire N__50490;
    wire N__50481;
    wire N__50472;
    wire N__50463;
    wire N__50454;
    wire N__50445;
    wire N__50436;
    wire N__50427;
    wire N__50418;
    wire N__50413;
    wire N__50410;
    wire N__50407;
    wire N__50404;
    wire N__50403;
    wire N__50400;
    wire N__50397;
    wire N__50394;
    wire N__50389;
    wire N__50386;
    wire N__50385;
    wire N__50384;
    wire N__50383;
    wire N__50380;
    wire N__50377;
    wire N__50374;
    wire N__50371;
    wire N__50368;
    wire N__50365;
    wire N__50362;
    wire N__50359;
    wire N__50354;
    wire N__50351;
    wire N__50348;
    wire N__50345;
    wire N__50342;
    wire N__50339;
    wire N__50332;
    wire N__50329;
    wire N__50328;
    wire N__50325;
    wire N__50322;
    wire N__50321;
    wire N__50318;
    wire N__50315;
    wire N__50312;
    wire N__50305;
    wire N__50304;
    wire N__50301;
    wire N__50298;
    wire N__50295;
    wire N__50292;
    wire N__50287;
    wire N__50284;
    wire N__50281;
    wire N__50278;
    wire N__50277;
    wire N__50276;
    wire N__50275;
    wire N__50274;
    wire N__50273;
    wire N__50272;
    wire N__50271;
    wire N__50270;
    wire N__50269;
    wire N__50268;
    wire N__50267;
    wire N__50266;
    wire N__50265;
    wire N__50264;
    wire N__50263;
    wire N__50262;
    wire N__50261;
    wire N__50260;
    wire N__50259;
    wire N__50258;
    wire N__50257;
    wire N__50256;
    wire N__50255;
    wire N__50254;
    wire N__50253;
    wire N__50252;
    wire N__50251;
    wire N__50250;
    wire N__50249;
    wire N__50248;
    wire N__50247;
    wire N__50246;
    wire N__50245;
    wire N__50244;
    wire N__50243;
    wire N__50242;
    wire N__50241;
    wire N__50240;
    wire N__50239;
    wire N__50238;
    wire N__50237;
    wire N__50236;
    wire N__50235;
    wire N__50234;
    wire N__50233;
    wire N__50232;
    wire N__50231;
    wire N__50230;
    wire N__50229;
    wire N__50228;
    wire N__50227;
    wire N__50226;
    wire N__50225;
    wire N__50224;
    wire N__50223;
    wire N__50222;
    wire N__50221;
    wire N__50220;
    wire N__50219;
    wire N__50218;
    wire N__50217;
    wire N__50216;
    wire N__50215;
    wire N__50214;
    wire N__50213;
    wire N__50212;
    wire N__50211;
    wire N__50210;
    wire N__50209;
    wire N__50208;
    wire N__50207;
    wire N__50206;
    wire N__50205;
    wire N__50204;
    wire N__50203;
    wire N__50202;
    wire N__50201;
    wire N__50200;
    wire N__50199;
    wire N__50198;
    wire N__50197;
    wire N__50196;
    wire N__50195;
    wire N__50194;
    wire N__50193;
    wire N__50192;
    wire N__50191;
    wire N__50190;
    wire N__50189;
    wire N__50188;
    wire N__50187;
    wire N__50186;
    wire N__50185;
    wire N__50184;
    wire N__50183;
    wire N__50182;
    wire N__50181;
    wire N__50180;
    wire N__50179;
    wire N__50178;
    wire N__50177;
    wire N__50176;
    wire N__50175;
    wire N__50174;
    wire N__50173;
    wire N__50172;
    wire N__50171;
    wire N__50170;
    wire N__50169;
    wire N__50168;
    wire N__50167;
    wire N__50166;
    wire N__50165;
    wire N__50164;
    wire N__50163;
    wire N__50162;
    wire N__50161;
    wire N__50160;
    wire N__50159;
    wire N__50158;
    wire N__50157;
    wire N__50156;
    wire N__50155;
    wire N__50154;
    wire N__50153;
    wire N__50152;
    wire N__50151;
    wire N__50150;
    wire N__50149;
    wire N__50148;
    wire N__50147;
    wire N__50146;
    wire N__50145;
    wire N__50144;
    wire N__50143;
    wire N__50142;
    wire N__50141;
    wire N__50140;
    wire N__50139;
    wire N__50138;
    wire N__50137;
    wire N__50136;
    wire N__50135;
    wire N__50134;
    wire N__50133;
    wire N__50132;
    wire N__50131;
    wire N__50130;
    wire N__50129;
    wire N__50128;
    wire N__50127;
    wire N__50126;
    wire N__49819;
    wire N__49816;
    wire N__49815;
    wire N__49814;
    wire N__49813;
    wire N__49812;
    wire N__49811;
    wire N__49798;
    wire N__49795;
    wire N__49792;
    wire N__49791;
    wire N__49790;
    wire N__49789;
    wire N__49788;
    wire N__49787;
    wire N__49786;
    wire N__49783;
    wire N__49780;
    wire N__49777;
    wire N__49774;
    wire N__49771;
    wire N__49768;
    wire N__49765;
    wire N__49762;
    wire N__49759;
    wire N__49756;
    wire N__49753;
    wire N__49750;
    wire N__49747;
    wire N__49746;
    wire N__49745;
    wire N__49744;
    wire N__49743;
    wire N__49742;
    wire N__49741;
    wire N__49740;
    wire N__49739;
    wire N__49738;
    wire N__49737;
    wire N__49736;
    wire N__49735;
    wire N__49734;
    wire N__49733;
    wire N__49732;
    wire N__49731;
    wire N__49730;
    wire N__49729;
    wire N__49728;
    wire N__49727;
    wire N__49726;
    wire N__49725;
    wire N__49724;
    wire N__49723;
    wire N__49722;
    wire N__49721;
    wire N__49720;
    wire N__49719;
    wire N__49718;
    wire N__49717;
    wire N__49716;
    wire N__49715;
    wire N__49714;
    wire N__49713;
    wire N__49712;
    wire N__49711;
    wire N__49710;
    wire N__49709;
    wire N__49708;
    wire N__49707;
    wire N__49706;
    wire N__49705;
    wire N__49704;
    wire N__49703;
    wire N__49702;
    wire N__49701;
    wire N__49700;
    wire N__49699;
    wire N__49698;
    wire N__49697;
    wire N__49696;
    wire N__49695;
    wire N__49694;
    wire N__49693;
    wire N__49692;
    wire N__49691;
    wire N__49690;
    wire N__49689;
    wire N__49688;
    wire N__49687;
    wire N__49686;
    wire N__49685;
    wire N__49684;
    wire N__49683;
    wire N__49682;
    wire N__49681;
    wire N__49680;
    wire N__49679;
    wire N__49678;
    wire N__49677;
    wire N__49676;
    wire N__49675;
    wire N__49674;
    wire N__49673;
    wire N__49672;
    wire N__49671;
    wire N__49670;
    wire N__49669;
    wire N__49668;
    wire N__49667;
    wire N__49666;
    wire N__49665;
    wire N__49664;
    wire N__49663;
    wire N__49662;
    wire N__49661;
    wire N__49660;
    wire N__49657;
    wire N__49656;
    wire N__49655;
    wire N__49654;
    wire N__49653;
    wire N__49652;
    wire N__49651;
    wire N__49650;
    wire N__49649;
    wire N__49648;
    wire N__49647;
    wire N__49646;
    wire N__49645;
    wire N__49644;
    wire N__49643;
    wire N__49642;
    wire N__49641;
    wire N__49640;
    wire N__49639;
    wire N__49638;
    wire N__49637;
    wire N__49636;
    wire N__49633;
    wire N__49632;
    wire N__49631;
    wire N__49630;
    wire N__49629;
    wire N__49628;
    wire N__49627;
    wire N__49626;
    wire N__49625;
    wire N__49624;
    wire N__49623;
    wire N__49622;
    wire N__49621;
    wire N__49620;
    wire N__49619;
    wire N__49618;
    wire N__49617;
    wire N__49616;
    wire N__49615;
    wire N__49614;
    wire N__49613;
    wire N__49612;
    wire N__49611;
    wire N__49610;
    wire N__49609;
    wire N__49608;
    wire N__49607;
    wire N__49604;
    wire N__49603;
    wire N__49318;
    wire N__49315;
    wire N__49312;
    wire N__49311;
    wire N__49308;
    wire N__49305;
    wire N__49304;
    wire N__49299;
    wire N__49296;
    wire N__49293;
    wire N__49288;
    wire N__49285;
    wire N__49284;
    wire N__49281;
    wire N__49278;
    wire N__49275;
    wire N__49274;
    wire N__49269;
    wire N__49266;
    wire N__49263;
    wire N__49258;
    wire N__49255;
    wire N__49254;
    wire N__49251;
    wire N__49248;
    wire N__49243;
    wire N__49242;
    wire N__49239;
    wire N__49236;
    wire N__49233;
    wire N__49228;
    wire N__49225;
    wire N__49224;
    wire N__49221;
    wire N__49218;
    wire N__49213;
    wire N__49212;
    wire N__49209;
    wire N__49206;
    wire N__49203;
    wire N__49198;
    wire N__49195;
    wire N__49194;
    wire N__49189;
    wire N__49188;
    wire N__49185;
    wire N__49182;
    wire N__49179;
    wire N__49174;
    wire N__49171;
    wire N__49170;
    wire N__49165;
    wire N__49164;
    wire N__49161;
    wire N__49158;
    wire N__49155;
    wire N__49150;
    wire N__49147;
    wire N__49146;
    wire N__49143;
    wire N__49140;
    wire N__49139;
    wire N__49134;
    wire N__49131;
    wire N__49128;
    wire N__49123;
    wire N__49120;
    wire N__49119;
    wire N__49116;
    wire N__49113;
    wire N__49112;
    wire N__49107;
    wire N__49104;
    wire N__49101;
    wire N__49096;
    wire N__49093;
    wire N__49092;
    wire N__49089;
    wire N__49086;
    wire N__49085;
    wire N__49080;
    wire N__49077;
    wire N__49074;
    wire N__49069;
    wire N__49066;
    wire N__49065;
    wire N__49062;
    wire N__49061;
    wire N__49058;
    wire N__49055;
    wire N__49052;
    wire N__49047;
    wire N__49042;
    wire N__49039;
    wire N__49038;
    wire N__49037;
    wire N__49034;
    wire N__49031;
    wire N__49028;
    wire N__49023;
    wire N__49018;
    wire N__49015;
    wire N__49014;
    wire N__49011;
    wire N__49008;
    wire N__49007;
    wire N__49002;
    wire N__48999;
    wire N__48996;
    wire N__48991;
    wire N__48988;
    wire N__48987;
    wire N__48984;
    wire N__48981;
    wire N__48980;
    wire N__48975;
    wire N__48972;
    wire N__48969;
    wire N__48964;
    wire N__48961;
    wire N__48960;
    wire N__48955;
    wire N__48954;
    wire N__48951;
    wire N__48948;
    wire N__48945;
    wire N__48940;
    wire N__48937;
    wire N__48934;
    wire N__48933;
    wire N__48930;
    wire N__48927;
    wire N__48926;
    wire N__48921;
    wire N__48918;
    wire N__48915;
    wire N__48910;
    wire N__48907;
    wire N__48906;
    wire N__48903;
    wire N__48900;
    wire N__48895;
    wire N__48894;
    wire N__48891;
    wire N__48888;
    wire N__48885;
    wire N__48880;
    wire N__48877;
    wire N__48876;
    wire N__48875;
    wire N__48870;
    wire N__48867;
    wire N__48864;
    wire N__48859;
    wire N__48856;
    wire N__48853;
    wire N__48852;
    wire N__48849;
    wire N__48846;
    wire N__48845;
    wire N__48842;
    wire N__48839;
    wire N__48836;
    wire N__48833;
    wire N__48830;
    wire N__48827;
    wire N__48824;
    wire N__48819;
    wire N__48814;
    wire N__48811;
    wire N__48810;
    wire N__48807;
    wire N__48804;
    wire N__48801;
    wire N__48798;
    wire N__48797;
    wire N__48792;
    wire N__48789;
    wire N__48786;
    wire N__48781;
    wire N__48778;
    wire N__48775;
    wire N__48774;
    wire N__48771;
    wire N__48768;
    wire N__48765;
    wire N__48764;
    wire N__48761;
    wire N__48758;
    wire N__48755;
    wire N__48752;
    wire N__48745;
    wire N__48742;
    wire N__48741;
    wire N__48736;
    wire N__48735;
    wire N__48732;
    wire N__48729;
    wire N__48726;
    wire N__48721;
    wire N__48718;
    wire N__48717;
    wire N__48716;
    wire N__48711;
    wire N__48708;
    wire N__48705;
    wire N__48700;
    wire N__48697;
    wire N__48696;
    wire N__48693;
    wire N__48690;
    wire N__48689;
    wire N__48684;
    wire N__48681;
    wire N__48678;
    wire N__48673;
    wire N__48670;
    wire N__48667;
    wire N__48666;
    wire N__48663;
    wire N__48662;
    wire N__48659;
    wire N__48656;
    wire N__48653;
    wire N__48650;
    wire N__48647;
    wire N__48640;
    wire N__48637;
    wire N__48636;
    wire N__48635;
    wire N__48630;
    wire N__48627;
    wire N__48624;
    wire N__48619;
    wire N__48616;
    wire N__48615;
    wire N__48612;
    wire N__48609;
    wire N__48604;
    wire N__48603;
    wire N__48600;
    wire N__48597;
    wire N__48594;
    wire N__48589;
    wire N__48586;
    wire N__48583;
    wire N__48580;
    wire N__48579;
    wire N__48578;
    wire N__48575;
    wire N__48572;
    wire N__48569;
    wire N__48566;
    wire N__48563;
    wire N__48560;
    wire N__48559;
    wire N__48556;
    wire N__48551;
    wire N__48548;
    wire N__48541;
    wire N__48538;
    wire N__48537;
    wire N__48534;
    wire N__48531;
    wire N__48530;
    wire N__48529;
    wire N__48524;
    wire N__48521;
    wire N__48518;
    wire N__48515;
    wire N__48512;
    wire N__48505;
    wire N__48502;
    wire N__48499;
    wire N__48498;
    wire N__48497;
    wire N__48492;
    wire N__48489;
    wire N__48486;
    wire N__48485;
    wire N__48482;
    wire N__48479;
    wire N__48476;
    wire N__48469;
    wire N__48466;
    wire N__48465;
    wire N__48462;
    wire N__48459;
    wire N__48456;
    wire N__48455;
    wire N__48452;
    wire N__48451;
    wire N__48448;
    wire N__48445;
    wire N__48442;
    wire N__48439;
    wire N__48430;
    wire N__48427;
    wire N__48426;
    wire N__48423;
    wire N__48420;
    wire N__48419;
    wire N__48416;
    wire N__48413;
    wire N__48410;
    wire N__48407;
    wire N__48404;
    wire N__48403;
    wire N__48400;
    wire N__48395;
    wire N__48392;
    wire N__48385;
    wire N__48382;
    wire N__48381;
    wire N__48378;
    wire N__48375;
    wire N__48374;
    wire N__48373;
    wire N__48370;
    wire N__48367;
    wire N__48364;
    wire N__48361;
    wire N__48356;
    wire N__48353;
    wire N__48346;
    wire N__48343;
    wire N__48342;
    wire N__48341;
    wire N__48338;
    wire N__48333;
    wire N__48330;
    wire N__48327;
    wire N__48326;
    wire N__48323;
    wire N__48320;
    wire N__48317;
    wire N__48310;
    wire N__48307;
    wire N__48304;
    wire N__48303;
    wire N__48302;
    wire N__48299;
    wire N__48296;
    wire N__48293;
    wire N__48288;
    wire N__48285;
    wire N__48284;
    wire N__48279;
    wire N__48276;
    wire N__48271;
    wire N__48268;
    wire N__48267;
    wire N__48266;
    wire N__48265;
    wire N__48264;
    wire N__48263;
    wire N__48262;
    wire N__48261;
    wire N__48244;
    wire N__48241;
    wire N__48238;
    wire N__48235;
    wire N__48234;
    wire N__48233;
    wire N__48230;
    wire N__48227;
    wire N__48224;
    wire N__48221;
    wire N__48220;
    wire N__48217;
    wire N__48214;
    wire N__48211;
    wire N__48208;
    wire N__48203;
    wire N__48198;
    wire N__48193;
    wire N__48190;
    wire N__48189;
    wire N__48188;
    wire N__48185;
    wire N__48182;
    wire N__48179;
    wire N__48176;
    wire N__48175;
    wire N__48172;
    wire N__48169;
    wire N__48166;
    wire N__48163;
    wire N__48158;
    wire N__48153;
    wire N__48148;
    wire N__48145;
    wire N__48144;
    wire N__48143;
    wire N__48140;
    wire N__48137;
    wire N__48134;
    wire N__48133;
    wire N__48130;
    wire N__48127;
    wire N__48124;
    wire N__48121;
    wire N__48118;
    wire N__48115;
    wire N__48110;
    wire N__48103;
    wire N__48100;
    wire N__48099;
    wire N__48096;
    wire N__48093;
    wire N__48090;
    wire N__48087;
    wire N__48086;
    wire N__48085;
    wire N__48082;
    wire N__48079;
    wire N__48074;
    wire N__48067;
    wire N__48064;
    wire N__48061;
    wire N__48058;
    wire N__48057;
    wire N__48056;
    wire N__48053;
    wire N__48050;
    wire N__48049;
    wire N__48046;
    wire N__48043;
    wire N__48040;
    wire N__48037;
    wire N__48034;
    wire N__48027;
    wire N__48022;
    wire N__48019;
    wire N__48018;
    wire N__48017;
    wire N__48012;
    wire N__48009;
    wire N__48006;
    wire N__48005;
    wire N__48002;
    wire N__47999;
    wire N__47996;
    wire N__47989;
    wire N__47986;
    wire N__47985;
    wire N__47982;
    wire N__47981;
    wire N__47978;
    wire N__47973;
    wire N__47968;
    wire N__47967;
    wire N__47964;
    wire N__47961;
    wire N__47956;
    wire N__47953;
    wire N__47952;
    wire N__47949;
    wire N__47948;
    wire N__47945;
    wire N__47942;
    wire N__47939;
    wire N__47936;
    wire N__47933;
    wire N__47930;
    wire N__47927;
    wire N__47926;
    wire N__47923;
    wire N__47918;
    wire N__47915;
    wire N__47908;
    wire N__47905;
    wire N__47902;
    wire N__47901;
    wire N__47900;
    wire N__47897;
    wire N__47894;
    wire N__47893;
    wire N__47890;
    wire N__47885;
    wire N__47882;
    wire N__47879;
    wire N__47876;
    wire N__47873;
    wire N__47866;
    wire N__47863;
    wire N__47862;
    wire N__47861;
    wire N__47860;
    wire N__47855;
    wire N__47852;
    wire N__47849;
    wire N__47846;
    wire N__47841;
    wire N__47836;
    wire N__47833;
    wire N__47830;
    wire N__47829;
    wire N__47826;
    wire N__47823;
    wire N__47822;
    wire N__47821;
    wire N__47816;
    wire N__47811;
    wire N__47806;
    wire N__47803;
    wire N__47800;
    wire N__47797;
    wire N__47796;
    wire N__47795;
    wire N__47792;
    wire N__47789;
    wire N__47786;
    wire N__47785;
    wire N__47780;
    wire N__47777;
    wire N__47774;
    wire N__47771;
    wire N__47768;
    wire N__47765;
    wire N__47758;
    wire N__47755;
    wire N__47752;
    wire N__47751;
    wire N__47750;
    wire N__47747;
    wire N__47744;
    wire N__47741;
    wire N__47736;
    wire N__47733;
    wire N__47732;
    wire N__47729;
    wire N__47726;
    wire N__47723;
    wire N__47716;
    wire N__47713;
    wire N__47710;
    wire N__47709;
    wire N__47708;
    wire N__47705;
    wire N__47702;
    wire N__47701;
    wire N__47698;
    wire N__47693;
    wire N__47690;
    wire N__47687;
    wire N__47682;
    wire N__47677;
    wire N__47674;
    wire N__47673;
    wire N__47672;
    wire N__47669;
    wire N__47666;
    wire N__47665;
    wire N__47662;
    wire N__47659;
    wire N__47656;
    wire N__47653;
    wire N__47650;
    wire N__47643;
    wire N__47638;
    wire N__47635;
    wire N__47632;
    wire N__47631;
    wire N__47630;
    wire N__47627;
    wire N__47624;
    wire N__47621;
    wire N__47620;
    wire N__47617;
    wire N__47614;
    wire N__47611;
    wire N__47608;
    wire N__47603;
    wire N__47598;
    wire N__47593;
    wire N__47590;
    wire N__47587;
    wire N__47586;
    wire N__47585;
    wire N__47582;
    wire N__47579;
    wire N__47578;
    wire N__47575;
    wire N__47570;
    wire N__47567;
    wire N__47564;
    wire N__47559;
    wire N__47554;
    wire N__47551;
    wire N__47548;
    wire N__47545;
    wire N__47542;
    wire N__47539;
    wire N__47536;
    wire N__47533;
    wire N__47530;
    wire N__47527;
    wire N__47524;
    wire N__47521;
    wire N__47518;
    wire N__47517;
    wire N__47512;
    wire N__47509;
    wire N__47508;
    wire N__47507;
    wire N__47504;
    wire N__47501;
    wire N__47498;
    wire N__47495;
    wire N__47492;
    wire N__47489;
    wire N__47482;
    wire N__47479;
    wire N__47478;
    wire N__47477;
    wire N__47470;
    wire N__47469;
    wire N__47466;
    wire N__47463;
    wire N__47460;
    wire N__47457;
    wire N__47452;
    wire N__47449;
    wire N__47448;
    wire N__47447;
    wire N__47444;
    wire N__47441;
    wire N__47438;
    wire N__47437;
    wire N__47434;
    wire N__47431;
    wire N__47428;
    wire N__47425;
    wire N__47422;
    wire N__47415;
    wire N__47410;
    wire N__47407;
    wire N__47404;
    wire N__47401;
    wire N__47400;
    wire N__47399;
    wire N__47396;
    wire N__47393;
    wire N__47390;
    wire N__47383;
    wire N__47380;
    wire N__47377;
    wire N__47374;
    wire N__47371;
    wire N__47368;
    wire N__47365;
    wire N__47362;
    wire N__47359;
    wire N__47356;
    wire N__47353;
    wire N__47350;
    wire N__47347;
    wire N__47344;
    wire N__47341;
    wire N__47338;
    wire N__47335;
    wire N__47332;
    wire N__47329;
    wire N__47326;
    wire N__47323;
    wire N__47320;
    wire N__47317;
    wire N__47314;
    wire N__47313;
    wire N__47308;
    wire N__47305;
    wire N__47302;
    wire N__47301;
    wire N__47300;
    wire N__47297;
    wire N__47292;
    wire N__47287;
    wire N__47284;
    wire N__47281;
    wire N__47280;
    wire N__47279;
    wire N__47278;
    wire N__47277;
    wire N__47276;
    wire N__47275;
    wire N__47274;
    wire N__47273;
    wire N__47272;
    wire N__47271;
    wire N__47270;
    wire N__47269;
    wire N__47268;
    wire N__47267;
    wire N__47266;
    wire N__47265;
    wire N__47254;
    wire N__47251;
    wire N__47246;
    wire N__47241;
    wire N__47234;
    wire N__47227;
    wire N__47226;
    wire N__47225;
    wire N__47224;
    wire N__47223;
    wire N__47220;
    wire N__47219;
    wire N__47216;
    wire N__47215;
    wire N__47212;
    wire N__47203;
    wire N__47198;
    wire N__47193;
    wire N__47192;
    wire N__47189;
    wire N__47188;
    wire N__47185;
    wire N__47182;
    wire N__47179;
    wire N__47170;
    wire N__47167;
    wire N__47164;
    wire N__47161;
    wire N__47146;
    wire N__47145;
    wire N__47140;
    wire N__47137;
    wire N__47136;
    wire N__47133;
    wire N__47130;
    wire N__47125;
    wire N__47122;
    wire N__47119;
    wire N__47116;
    wire N__47113;
    wire N__47112;
    wire N__47111;
    wire N__47108;
    wire N__47105;
    wire N__47102;
    wire N__47095;
    wire N__47092;
    wire N__47089;
    wire N__47086;
    wire N__47083;
    wire N__47080;
    wire N__47079;
    wire N__47078;
    wire N__47073;
    wire N__47070;
    wire N__47067;
    wire N__47062;
    wire N__47059;
    wire N__47056;
    wire N__47053;
    wire N__47050;
    wire N__47047;
    wire N__47044;
    wire N__47041;
    wire N__47038;
    wire N__47035;
    wire N__47032;
    wire N__47029;
    wire N__47026;
    wire N__47023;
    wire N__47020;
    wire N__47017;
    wire N__47014;
    wire N__47011;
    wire N__47008;
    wire N__47005;
    wire N__47002;
    wire N__46999;
    wire N__46996;
    wire N__46995;
    wire N__46994;
    wire N__46993;
    wire N__46992;
    wire N__46991;
    wire N__46988;
    wire N__46981;
    wire N__46980;
    wire N__46979;
    wire N__46976;
    wire N__46975;
    wire N__46974;
    wire N__46973;
    wire N__46972;
    wire N__46971;
    wire N__46970;
    wire N__46969;
    wire N__46966;
    wire N__46965;
    wire N__46962;
    wire N__46959;
    wire N__46950;
    wire N__46937;
    wire N__46932;
    wire N__46931;
    wire N__46930;
    wire N__46929;
    wire N__46928;
    wire N__46927;
    wire N__46926;
    wire N__46925;
    wire N__46924;
    wire N__46921;
    wire N__46918;
    wire N__46915;
    wire N__46912;
    wire N__46909;
    wire N__46906;
    wire N__46903;
    wire N__46902;
    wire N__46901;
    wire N__46898;
    wire N__46897;
    wire N__46886;
    wire N__46881;
    wire N__46878;
    wire N__46873;
    wire N__46860;
    wire N__46849;
    wire N__46846;
    wire N__46843;
    wire N__46840;
    wire N__46837;
    wire N__46834;
    wire N__46831;
    wire N__46828;
    wire N__46825;
    wire N__46822;
    wire N__46819;
    wire N__46818;
    wire N__46817;
    wire N__46816;
    wire N__46815;
    wire N__46814;
    wire N__46813;
    wire N__46812;
    wire N__46811;
    wire N__46810;
    wire N__46809;
    wire N__46804;
    wire N__46803;
    wire N__46802;
    wire N__46801;
    wire N__46800;
    wire N__46799;
    wire N__46798;
    wire N__46797;
    wire N__46796;
    wire N__46791;
    wire N__46788;
    wire N__46785;
    wire N__46774;
    wire N__46773;
    wire N__46772;
    wire N__46771;
    wire N__46768;
    wire N__46765;
    wire N__46762;
    wire N__46759;
    wire N__46758;
    wire N__46757;
    wire N__46756;
    wire N__46753;
    wire N__46750;
    wire N__46749;
    wire N__46746;
    wire N__46745;
    wire N__46744;
    wire N__46743;
    wire N__46742;
    wire N__46741;
    wire N__46740;
    wire N__46739;
    wire N__46736;
    wire N__46733;
    wire N__46724;
    wire N__46717;
    wire N__46708;
    wire N__46707;
    wire N__46706;
    wire N__46705;
    wire N__46704;
    wire N__46703;
    wire N__46702;
    wire N__46701;
    wire N__46700;
    wire N__46699;
    wire N__46698;
    wire N__46697;
    wire N__46696;
    wire N__46695;
    wire N__46694;
    wire N__46693;
    wire N__46692;
    wire N__46691;
    wire N__46690;
    wire N__46689;
    wire N__46688;
    wire N__46687;
    wire N__46686;
    wire N__46685;
    wire N__46684;
    wire N__46683;
    wire N__46682;
    wire N__46681;
    wire N__46680;
    wire N__46679;
    wire N__46678;
    wire N__46671;
    wire N__46668;
    wire N__46665;
    wire N__46662;
    wire N__46659;
    wire N__46652;
    wire N__46651;
    wire N__46648;
    wire N__46647;
    wire N__46644;
    wire N__46639;
    wire N__46636;
    wire N__46633;
    wire N__46628;
    wire N__46625;
    wire N__46622;
    wire N__46617;
    wire N__46614;
    wire N__46609;
    wire N__46604;
    wire N__46593;
    wire N__46586;
    wire N__46577;
    wire N__46566;
    wire N__46561;
    wire N__46554;
    wire N__46551;
    wire N__46544;
    wire N__46539;
    wire N__46532;
    wire N__46531;
    wire N__46530;
    wire N__46529;
    wire N__46528;
    wire N__46527;
    wire N__46522;
    wire N__46517;
    wire N__46514;
    wire N__46507;
    wire N__46504;
    wire N__46501;
    wire N__46490;
    wire N__46485;
    wire N__46482;
    wire N__46477;
    wire N__46474;
    wire N__46467;
    wire N__46462;
    wire N__46457;
    wire N__46452;
    wire N__46443;
    wire N__46440;
    wire N__46423;
    wire N__46422;
    wire N__46421;
    wire N__46420;
    wire N__46419;
    wire N__46418;
    wire N__46415;
    wire N__46412;
    wire N__46409;
    wire N__46408;
    wire N__46407;
    wire N__46406;
    wire N__46403;
    wire N__46400;
    wire N__46397;
    wire N__46392;
    wire N__46389;
    wire N__46386;
    wire N__46383;
    wire N__46380;
    wire N__46379;
    wire N__46378;
    wire N__46377;
    wire N__46376;
    wire N__46375;
    wire N__46374;
    wire N__46373;
    wire N__46372;
    wire N__46371;
    wire N__46370;
    wire N__46369;
    wire N__46368;
    wire N__46367;
    wire N__46366;
    wire N__46363;
    wire N__46358;
    wire N__46353;
    wire N__46348;
    wire N__46345;
    wire N__46344;
    wire N__46343;
    wire N__46342;
    wire N__46341;
    wire N__46340;
    wire N__46339;
    wire N__46336;
    wire N__46335;
    wire N__46334;
    wire N__46333;
    wire N__46332;
    wire N__46331;
    wire N__46330;
    wire N__46329;
    wire N__46328;
    wire N__46327;
    wire N__46326;
    wire N__46325;
    wire N__46324;
    wire N__46323;
    wire N__46322;
    wire N__46321;
    wire N__46320;
    wire N__46319;
    wire N__46316;
    wire N__46315;
    wire N__46312;
    wire N__46309;
    wire N__46306;
    wire N__46305;
    wire N__46304;
    wire N__46303;
    wire N__46302;
    wire N__46301;
    wire N__46298;
    wire N__46297;
    wire N__46296;
    wire N__46295;
    wire N__46294;
    wire N__46293;
    wire N__46292;
    wire N__46291;
    wire N__46290;
    wire N__46287;
    wire N__46284;
    wire N__46283;
    wire N__46280;
    wire N__46277;
    wire N__46276;
    wire N__46275;
    wire N__46274;
    wire N__46273;
    wire N__46270;
    wire N__46267;
    wire N__46264;
    wire N__46261;
    wire N__46260;
    wire N__46259;
    wire N__46258;
    wire N__46257;
    wire N__46256;
    wire N__46255;
    wire N__46250;
    wire N__46243;
    wire N__46240;
    wire N__46237;
    wire N__46234;
    wire N__46233;
    wire N__46232;
    wire N__46231;
    wire N__46230;
    wire N__46229;
    wire N__46228;
    wire N__46225;
    wire N__46222;
    wire N__46219;
    wire N__46218;
    wire N__46217;
    wire N__46216;
    wire N__46215;
    wire N__46214;
    wire N__46213;
    wire N__46212;
    wire N__46211;
    wire N__46210;
    wire N__46209;
    wire N__46208;
    wire N__46205;
    wire N__46202;
    wire N__46199;
    wire N__46196;
    wire N__46193;
    wire N__46190;
    wire N__46187;
    wire N__46184;
    wire N__46181;
    wire N__46178;
    wire N__46175;
    wire N__46172;
    wire N__46169;
    wire N__46168;
    wire N__46165;
    wire N__46162;
    wire N__46159;
    wire N__46156;
    wire N__46153;
    wire N__46152;
    wire N__46149;
    wire N__46140;
    wire N__46137;
    wire N__46134;
    wire N__46131;
    wire N__46128;
    wire N__46123;
    wire N__46120;
    wire N__46117;
    wire N__46114;
    wire N__46111;
    wire N__46108;
    wire N__46105;
    wire N__46102;
    wire N__46099;
    wire N__46098;
    wire N__46095;
    wire N__46086;
    wire N__46083;
    wire N__46080;
    wire N__46077;
    wire N__46074;
    wire N__46065;
    wire N__46062;
    wire N__46059;
    wire N__46056;
    wire N__46053;
    wire N__46050;
    wire N__46047;
    wire N__46042;
    wire N__46039;
    wire N__46034;
    wire N__46027;
    wire N__46026;
    wire N__46023;
    wire N__46020;
    wire N__46019;
    wire N__46016;
    wire N__46011;
    wire N__46008;
    wire N__46007;
    wire N__46006;
    wire N__46003;
    wire N__46000;
    wire N__45999;
    wire N__45998;
    wire N__45997;
    wire N__45996;
    wire N__45995;
    wire N__45994;
    wire N__45993;
    wire N__45992;
    wire N__45991;
    wire N__45988;
    wire N__45985;
    wire N__45982;
    wire N__45981;
    wire N__45978;
    wire N__45975;
    wire N__45972;
    wire N__45971;
    wire N__45968;
    wire N__45967;
    wire N__45964;
    wire N__45963;
    wire N__45960;
    wire N__45959;
    wire N__45956;
    wire N__45949;
    wire N__45940;
    wire N__45931;
    wire N__45930;
    wire N__45929;
    wire N__45928;
    wire N__45927;
    wire N__45926;
    wire N__45925;
    wire N__45922;
    wire N__45921;
    wire N__45918;
    wire N__45913;
    wire N__45906;
    wire N__45903;
    wire N__45898;
    wire N__45889;
    wire N__45886;
    wire N__45877;
    wire N__45870;
    wire N__45865;
    wire N__45860;
    wire N__45851;
    wire N__45848;
    wire N__45841;
    wire N__45834;
    wire N__45825;
    wire N__45822;
    wire N__45817;
    wire N__45814;
    wire N__45811;
    wire N__45806;
    wire N__45801;
    wire N__45796;
    wire N__45793;
    wire N__45790;
    wire N__45787;
    wire N__45784;
    wire N__45781;
    wire N__45778;
    wire N__45775;
    wire N__45772;
    wire N__45769;
    wire N__45764;
    wire N__45753;
    wire N__45738;
    wire N__45729;
    wire N__45726;
    wire N__45723;
    wire N__45720;
    wire N__45717;
    wire N__45714;
    wire N__45711;
    wire N__45708;
    wire N__45703;
    wire N__45694;
    wire N__45673;
    wire N__45670;
    wire N__45667;
    wire N__45664;
    wire N__45661;
    wire N__45656;
    wire N__45649;
    wire N__45640;
    wire N__45631;
    wire N__45622;
    wire N__45615;
    wire N__45608;
    wire N__45599;
    wire N__45574;
    wire N__45571;
    wire N__45570;
    wire N__45567;
    wire N__45564;
    wire N__45563;
    wire N__45560;
    wire N__45557;
    wire N__45554;
    wire N__45547;
    wire N__45544;
    wire N__45541;
    wire N__45538;
    wire N__45535;
    wire N__45532;
    wire N__45529;
    wire N__45526;
    wire N__45523;
    wire N__45520;
    wire N__45517;
    wire N__45516;
    wire N__45513;
    wire N__45510;
    wire N__45507;
    wire N__45504;
    wire N__45503;
    wire N__45500;
    wire N__45497;
    wire N__45494;
    wire N__45487;
    wire N__45484;
    wire N__45481;
    wire N__45478;
    wire N__45475;
    wire N__45472;
    wire N__45469;
    wire N__45466;
    wire N__45463;
    wire N__45460;
    wire N__45457;
    wire N__45454;
    wire N__45451;
    wire N__45448;
    wire N__45445;
    wire N__45442;
    wire N__45441;
    wire N__45440;
    wire N__45437;
    wire N__45434;
    wire N__45431;
    wire N__45428;
    wire N__45425;
    wire N__45422;
    wire N__45419;
    wire N__45414;
    wire N__45409;
    wire N__45406;
    wire N__45403;
    wire N__45400;
    wire N__45397;
    wire N__45394;
    wire N__45391;
    wire N__45390;
    wire N__45387;
    wire N__45386;
    wire N__45383;
    wire N__45380;
    wire N__45377;
    wire N__45374;
    wire N__45367;
    wire N__45364;
    wire N__45361;
    wire N__45360;
    wire N__45357;
    wire N__45354;
    wire N__45351;
    wire N__45348;
    wire N__45343;
    wire N__45340;
    wire N__45339;
    wire N__45338;
    wire N__45335;
    wire N__45332;
    wire N__45329;
    wire N__45324;
    wire N__45323;
    wire N__45322;
    wire N__45321;
    wire N__45316;
    wire N__45311;
    wire N__45310;
    wire N__45309;
    wire N__45308;
    wire N__45307;
    wire N__45306;
    wire N__45305;
    wire N__45304;
    wire N__45303;
    wire N__45302;
    wire N__45301;
    wire N__45298;
    wire N__45297;
    wire N__45296;
    wire N__45291;
    wire N__45282;
    wire N__45281;
    wire N__45280;
    wire N__45279;
    wire N__45272;
    wire N__45265;
    wire N__45262;
    wire N__45257;
    wire N__45252;
    wire N__45251;
    wire N__45250;
    wire N__45249;
    wire N__45246;
    wire N__45243;
    wire N__45240;
    wire N__45239;
    wire N__45238;
    wire N__45237;
    wire N__45236;
    wire N__45235;
    wire N__45232;
    wire N__45229;
    wire N__45224;
    wire N__45223;
    wire N__45222;
    wire N__45219;
    wire N__45212;
    wire N__45211;
    wire N__45208;
    wire N__45205;
    wire N__45202;
    wire N__45191;
    wire N__45188;
    wire N__45183;
    wire N__45178;
    wire N__45173;
    wire N__45170;
    wire N__45163;
    wire N__45158;
    wire N__45155;
    wire N__45150;
    wire N__45139;
    wire N__45138;
    wire N__45137;
    wire N__45136;
    wire N__45135;
    wire N__45134;
    wire N__45133;
    wire N__45132;
    wire N__45131;
    wire N__45130;
    wire N__45127;
    wire N__45126;
    wire N__45125;
    wire N__45124;
    wire N__45123;
    wire N__45122;
    wire N__45121;
    wire N__45120;
    wire N__45119;
    wire N__45118;
    wire N__45117;
    wire N__45116;
    wire N__45113;
    wire N__45112;
    wire N__45105;
    wire N__45102;
    wire N__45099;
    wire N__45092;
    wire N__45085;
    wire N__45082;
    wire N__45077;
    wire N__45068;
    wire N__45067;
    wire N__45066;
    wire N__45065;
    wire N__45064;
    wire N__45063;
    wire N__45062;
    wire N__45061;
    wire N__45060;
    wire N__45057;
    wire N__45054;
    wire N__45051;
    wire N__45048;
    wire N__45047;
    wire N__45046;
    wire N__45043;
    wire N__45038;
    wire N__45033;
    wire N__45030;
    wire N__45027;
    wire N__45024;
    wire N__45021;
    wire N__45016;
    wire N__45005;
    wire N__45000;
    wire N__44995;
    wire N__44990;
    wire N__44983;
    wire N__44976;
    wire N__44973;
    wire N__44966;
    wire N__44963;
    wire N__44956;
    wire N__44947;
    wire N__44944;
    wire N__44941;
    wire N__44938;
    wire N__44935;
    wire N__44934;
    wire N__44933;
    wire N__44930;
    wire N__44927;
    wire N__44924;
    wire N__44923;
    wire N__44922;
    wire N__44921;
    wire N__44920;
    wire N__44919;
    wire N__44918;
    wire N__44917;
    wire N__44916;
    wire N__44915;
    wire N__44914;
    wire N__44913;
    wire N__44912;
    wire N__44911;
    wire N__44906;
    wire N__44903;
    wire N__44900;
    wire N__44897;
    wire N__44894;
    wire N__44891;
    wire N__44888;
    wire N__44885;
    wire N__44884;
    wire N__44883;
    wire N__44880;
    wire N__44877;
    wire N__44874;
    wire N__44871;
    wire N__44868;
    wire N__44867;
    wire N__44866;
    wire N__44865;
    wire N__44862;
    wire N__44859;
    wire N__44856;
    wire N__44853;
    wire N__44852;
    wire N__44849;
    wire N__44842;
    wire N__44837;
    wire N__44834;
    wire N__44833;
    wire N__44832;
    wire N__44829;
    wire N__44826;
    wire N__44823;
    wire N__44818;
    wire N__44815;
    wire N__44812;
    wire N__44811;
    wire N__44810;
    wire N__44809;
    wire N__44808;
    wire N__44807;
    wire N__44806;
    wire N__44803;
    wire N__44800;
    wire N__44799;
    wire N__44794;
    wire N__44789;
    wire N__44786;
    wire N__44783;
    wire N__44778;
    wire N__44775;
    wire N__44772;
    wire N__44769;
    wire N__44768;
    wire N__44765;
    wire N__44754;
    wire N__44751;
    wire N__44748;
    wire N__44745;
    wire N__44742;
    wire N__44739;
    wire N__44736;
    wire N__44731;
    wire N__44728;
    wire N__44721;
    wire N__44714;
    wire N__44711;
    wire N__44708;
    wire N__44705;
    wire N__44702;
    wire N__44699;
    wire N__44694;
    wire N__44689;
    wire N__44684;
    wire N__44675;
    wire N__44664;
    wire N__44653;
    wire N__44652;
    wire N__44651;
    wire N__44650;
    wire N__44647;
    wire N__44644;
    wire N__44641;
    wire N__44638;
    wire N__44635;
    wire N__44632;
    wire N__44629;
    wire N__44626;
    wire N__44625;
    wire N__44622;
    wire N__44619;
    wire N__44614;
    wire N__44611;
    wire N__44606;
    wire N__44603;
    wire N__44600;
    wire N__44593;
    wire N__44590;
    wire N__44587;
    wire N__44584;
    wire N__44581;
    wire N__44578;
    wire N__44577;
    wire N__44574;
    wire N__44573;
    wire N__44570;
    wire N__44567;
    wire N__44564;
    wire N__44563;
    wire N__44562;
    wire N__44559;
    wire N__44556;
    wire N__44553;
    wire N__44550;
    wire N__44547;
    wire N__44544;
    wire N__44533;
    wire N__44530;
    wire N__44527;
    wire N__44524;
    wire N__44521;
    wire N__44520;
    wire N__44517;
    wire N__44514;
    wire N__44513;
    wire N__44510;
    wire N__44507;
    wire N__44504;
    wire N__44501;
    wire N__44498;
    wire N__44495;
    wire N__44490;
    wire N__44489;
    wire N__44486;
    wire N__44483;
    wire N__44480;
    wire N__44473;
    wire N__44470;
    wire N__44467;
    wire N__44464;
    wire N__44461;
    wire N__44458;
    wire N__44455;
    wire N__44454;
    wire N__44453;
    wire N__44450;
    wire N__44447;
    wire N__44444;
    wire N__44443;
    wire N__44438;
    wire N__44435;
    wire N__44432;
    wire N__44431;
    wire N__44428;
    wire N__44425;
    wire N__44422;
    wire N__44419;
    wire N__44416;
    wire N__44407;
    wire N__44404;
    wire N__44401;
    wire N__44398;
    wire N__44395;
    wire N__44392;
    wire N__44389;
    wire N__44386;
    wire N__44383;
    wire N__44380;
    wire N__44377;
    wire N__44374;
    wire N__44371;
    wire N__44368;
    wire N__44365;
    wire N__44362;
    wire N__44359;
    wire N__44356;
    wire N__44353;
    wire N__44350;
    wire N__44347;
    wire N__44344;
    wire N__44341;
    wire N__44338;
    wire N__44335;
    wire N__44332;
    wire N__44331;
    wire N__44328;
    wire N__44327;
    wire N__44324;
    wire N__44321;
    wire N__44318;
    wire N__44311;
    wire N__44310;
    wire N__44307;
    wire N__44304;
    wire N__44303;
    wire N__44298;
    wire N__44295;
    wire N__44292;
    wire N__44289;
    wire N__44286;
    wire N__44281;
    wire N__44278;
    wire N__44275;
    wire N__44272;
    wire N__44269;
    wire N__44266;
    wire N__44265;
    wire N__44262;
    wire N__44259;
    wire N__44256;
    wire N__44253;
    wire N__44252;
    wire N__44249;
    wire N__44246;
    wire N__44243;
    wire N__44236;
    wire N__44233;
    wire N__44230;
    wire N__44227;
    wire N__44224;
    wire N__44221;
    wire N__44218;
    wire N__44215;
    wire N__44212;
    wire N__44209;
    wire N__44206;
    wire N__44203;
    wire N__44202;
    wire N__44201;
    wire N__44198;
    wire N__44195;
    wire N__44192;
    wire N__44189;
    wire N__44186;
    wire N__44183;
    wire N__44180;
    wire N__44179;
    wire N__44178;
    wire N__44173;
    wire N__44170;
    wire N__44167;
    wire N__44164;
    wire N__44161;
    wire N__44152;
    wire N__44149;
    wire N__44146;
    wire N__44143;
    wire N__44140;
    wire N__44139;
    wire N__44136;
    wire N__44135;
    wire N__44132;
    wire N__44127;
    wire N__44126;
    wire N__44123;
    wire N__44120;
    wire N__44119;
    wire N__44116;
    wire N__44111;
    wire N__44108;
    wire N__44105;
    wire N__44102;
    wire N__44095;
    wire N__44092;
    wire N__44089;
    wire N__44086;
    wire N__44083;
    wire N__44082;
    wire N__44081;
    wire N__44080;
    wire N__44079;
    wire N__44078;
    wire N__44077;
    wire N__44074;
    wire N__44073;
    wire N__44072;
    wire N__44071;
    wire N__44070;
    wire N__44069;
    wire N__44068;
    wire N__44067;
    wire N__44066;
    wire N__44063;
    wire N__44060;
    wire N__44057;
    wire N__44056;
    wire N__44055;
    wire N__44054;
    wire N__44053;
    wire N__44052;
    wire N__44051;
    wire N__44050;
    wire N__44049;
    wire N__44046;
    wire N__44043;
    wire N__44040;
    wire N__44037;
    wire N__44020;
    wire N__44019;
    wire N__44018;
    wire N__44017;
    wire N__44010;
    wire N__43999;
    wire N__43998;
    wire N__43997;
    wire N__43996;
    wire N__43993;
    wire N__43988;
    wire N__43987;
    wire N__43986;
    wire N__43985;
    wire N__43984;
    wire N__43983;
    wire N__43982;
    wire N__43981;
    wire N__43980;
    wire N__43977;
    wire N__43974;
    wire N__43967;
    wire N__43962;
    wire N__43959;
    wire N__43954;
    wire N__43949;
    wire N__43946;
    wire N__43941;
    wire N__43928;
    wire N__43923;
    wire N__43920;
    wire N__43913;
    wire N__43908;
    wire N__43901;
    wire N__43898;
    wire N__43891;
    wire N__43888;
    wire N__43885;
    wire N__43882;
    wire N__43873;
    wire N__43872;
    wire N__43869;
    wire N__43866;
    wire N__43863;
    wire N__43860;
    wire N__43859;
    wire N__43856;
    wire N__43853;
    wire N__43850;
    wire N__43845;
    wire N__43842;
    wire N__43837;
    wire N__43834;
    wire N__43831;
    wire N__43828;
    wire N__43825;
    wire N__43822;
    wire N__43819;
    wire N__43816;
    wire N__43813;
    wire N__43810;
    wire N__43807;
    wire N__43804;
    wire N__43801;
    wire N__43798;
    wire N__43797;
    wire N__43794;
    wire N__43793;
    wire N__43790;
    wire N__43789;
    wire N__43786;
    wire N__43785;
    wire N__43782;
    wire N__43779;
    wire N__43776;
    wire N__43773;
    wire N__43770;
    wire N__43767;
    wire N__43762;
    wire N__43757;
    wire N__43750;
    wire N__43747;
    wire N__43744;
    wire N__43741;
    wire N__43738;
    wire N__43735;
    wire N__43732;
    wire N__43729;
    wire N__43726;
    wire N__43723;
    wire N__43720;
    wire N__43717;
    wire N__43714;
    wire N__43711;
    wire N__43708;
    wire N__43705;
    wire N__43702;
    wire N__43701;
    wire N__43698;
    wire N__43695;
    wire N__43694;
    wire N__43689;
    wire N__43686;
    wire N__43681;
    wire N__43678;
    wire N__43675;
    wire N__43672;
    wire N__43669;
    wire N__43666;
    wire N__43663;
    wire N__43662;
    wire N__43661;
    wire N__43658;
    wire N__43657;
    wire N__43654;
    wire N__43651;
    wire N__43648;
    wire N__43645;
    wire N__43636;
    wire N__43633;
    wire N__43632;
    wire N__43629;
    wire N__43626;
    wire N__43625;
    wire N__43620;
    wire N__43617;
    wire N__43616;
    wire N__43613;
    wire N__43612;
    wire N__43609;
    wire N__43606;
    wire N__43603;
    wire N__43600;
    wire N__43591;
    wire N__43590;
    wire N__43589;
    wire N__43588;
    wire N__43585;
    wire N__43582;
    wire N__43579;
    wire N__43576;
    wire N__43573;
    wire N__43570;
    wire N__43569;
    wire N__43566;
    wire N__43563;
    wire N__43560;
    wire N__43557;
    wire N__43554;
    wire N__43551;
    wire N__43540;
    wire N__43537;
    wire N__43536;
    wire N__43535;
    wire N__43532;
    wire N__43529;
    wire N__43528;
    wire N__43527;
    wire N__43524;
    wire N__43521;
    wire N__43516;
    wire N__43513;
    wire N__43508;
    wire N__43505;
    wire N__43502;
    wire N__43495;
    wire N__43492;
    wire N__43489;
    wire N__43486;
    wire N__43483;
    wire N__43480;
    wire N__43477;
    wire N__43474;
    wire N__43471;
    wire N__43470;
    wire N__43469;
    wire N__43468;
    wire N__43465;
    wire N__43462;
    wire N__43459;
    wire N__43456;
    wire N__43453;
    wire N__43452;
    wire N__43447;
    wire N__43442;
    wire N__43439;
    wire N__43436;
    wire N__43429;
    wire N__43426;
    wire N__43423;
    wire N__43420;
    wire N__43417;
    wire N__43414;
    wire N__43411;
    wire N__43408;
    wire N__43405;
    wire N__43402;
    wire N__43399;
    wire N__43396;
    wire N__43393;
    wire N__43390;
    wire N__43387;
    wire N__43384;
    wire N__43381;
    wire N__43378;
    wire N__43375;
    wire N__43372;
    wire N__43371;
    wire N__43368;
    wire N__43365;
    wire N__43364;
    wire N__43359;
    wire N__43356;
    wire N__43351;
    wire N__43348;
    wire N__43345;
    wire N__43342;
    wire N__43339;
    wire N__43336;
    wire N__43333;
    wire N__43330;
    wire N__43327;
    wire N__43324;
    wire N__43321;
    wire N__43320;
    wire N__43317;
    wire N__43314;
    wire N__43313;
    wire N__43308;
    wire N__43305;
    wire N__43300;
    wire N__43297;
    wire N__43294;
    wire N__43291;
    wire N__43288;
    wire N__43287;
    wire N__43284;
    wire N__43281;
    wire N__43280;
    wire N__43277;
    wire N__43274;
    wire N__43271;
    wire N__43268;
    wire N__43263;
    wire N__43258;
    wire N__43255;
    wire N__43252;
    wire N__43249;
    wire N__43246;
    wire N__43243;
    wire N__43242;
    wire N__43241;
    wire N__43238;
    wire N__43233;
    wire N__43228;
    wire N__43225;
    wire N__43224;
    wire N__43221;
    wire N__43218;
    wire N__43217;
    wire N__43212;
    wire N__43209;
    wire N__43204;
    wire N__43201;
    wire N__43198;
    wire N__43195;
    wire N__43192;
    wire N__43189;
    wire N__43186;
    wire N__43183;
    wire N__43180;
    wire N__43177;
    wire N__43174;
    wire N__43171;
    wire N__43170;
    wire N__43167;
    wire N__43164;
    wire N__43163;
    wire N__43158;
    wire N__43155;
    wire N__43150;
    wire N__43147;
    wire N__43144;
    wire N__43141;
    wire N__43138;
    wire N__43135;
    wire N__43132;
    wire N__43129;
    wire N__43128;
    wire N__43127;
    wire N__43124;
    wire N__43119;
    wire N__43114;
    wire N__43111;
    wire N__43108;
    wire N__43107;
    wire N__43106;
    wire N__43103;
    wire N__43098;
    wire N__43093;
    wire N__43090;
    wire N__43089;
    wire N__43086;
    wire N__43083;
    wire N__43080;
    wire N__43077;
    wire N__43076;
    wire N__43071;
    wire N__43068;
    wire N__43063;
    wire N__43060;
    wire N__43057;
    wire N__43054;
    wire N__43053;
    wire N__43050;
    wire N__43047;
    wire N__43042;
    wire N__43041;
    wire N__43038;
    wire N__43035;
    wire N__43030;
    wire N__43027;
    wire N__43024;
    wire N__43021;
    wire N__43018;
    wire N__43017;
    wire N__43016;
    wire N__43013;
    wire N__43008;
    wire N__43003;
    wire N__43000;
    wire N__42999;
    wire N__42996;
    wire N__42993;
    wire N__42990;
    wire N__42987;
    wire N__42986;
    wire N__42981;
    wire N__42978;
    wire N__42973;
    wire N__42970;
    wire N__42967;
    wire N__42964;
    wire N__42961;
    wire N__42960;
    wire N__42959;
    wire N__42956;
    wire N__42953;
    wire N__42950;
    wire N__42943;
    wire N__42940;
    wire N__42937;
    wire N__42936;
    wire N__42933;
    wire N__42930;
    wire N__42929;
    wire N__42926;
    wire N__42923;
    wire N__42920;
    wire N__42913;
    wire N__42910;
    wire N__42907;
    wire N__42904;
    wire N__42901;
    wire N__42900;
    wire N__42899;
    wire N__42896;
    wire N__42893;
    wire N__42890;
    wire N__42883;
    wire N__42880;
    wire N__42877;
    wire N__42876;
    wire N__42873;
    wire N__42870;
    wire N__42869;
    wire N__42866;
    wire N__42863;
    wire N__42860;
    wire N__42853;
    wire N__42850;
    wire N__42847;
    wire N__42846;
    wire N__42843;
    wire N__42840;
    wire N__42839;
    wire N__42836;
    wire N__42833;
    wire N__42830;
    wire N__42823;
    wire N__42820;
    wire N__42819;
    wire N__42816;
    wire N__42813;
    wire N__42810;
    wire N__42807;
    wire N__42806;
    wire N__42801;
    wire N__42798;
    wire N__42793;
    wire N__42790;
    wire N__42787;
    wire N__42786;
    wire N__42785;
    wire N__42784;
    wire N__42783;
    wire N__42782;
    wire N__42781;
    wire N__42780;
    wire N__42779;
    wire N__42778;
    wire N__42777;
    wire N__42776;
    wire N__42775;
    wire N__42774;
    wire N__42773;
    wire N__42772;
    wire N__42771;
    wire N__42770;
    wire N__42769;
    wire N__42768;
    wire N__42767;
    wire N__42766;
    wire N__42765;
    wire N__42764;
    wire N__42763;
    wire N__42762;
    wire N__42761;
    wire N__42760;
    wire N__42759;
    wire N__42758;
    wire N__42749;
    wire N__42740;
    wire N__42731;
    wire N__42722;
    wire N__42713;
    wire N__42704;
    wire N__42699;
    wire N__42690;
    wire N__42687;
    wire N__42680;
    wire N__42671;
    wire N__42664;
    wire N__42661;
    wire N__42658;
    wire N__42655;
    wire N__42654;
    wire N__42651;
    wire N__42648;
    wire N__42645;
    wire N__42640;
    wire N__42639;
    wire N__42638;
    wire N__42635;
    wire N__42632;
    wire N__42629;
    wire N__42624;
    wire N__42623;
    wire N__42620;
    wire N__42617;
    wire N__42614;
    wire N__42607;
    wire N__42604;
    wire N__42601;
    wire N__42598;
    wire N__42595;
    wire N__42592;
    wire N__42591;
    wire N__42590;
    wire N__42583;
    wire N__42580;
    wire N__42577;
    wire N__42576;
    wire N__42575;
    wire N__42568;
    wire N__42565;
    wire N__42562;
    wire N__42559;
    wire N__42558;
    wire N__42555;
    wire N__42552;
    wire N__42551;
    wire N__42548;
    wire N__42545;
    wire N__42542;
    wire N__42535;
    wire N__42532;
    wire N__42529;
    wire N__42526;
    wire N__42525;
    wire N__42524;
    wire N__42519;
    wire N__42516;
    wire N__42513;
    wire N__42508;
    wire N__42505;
    wire N__42504;
    wire N__42503;
    wire N__42498;
    wire N__42495;
    wire N__42492;
    wire N__42487;
    wire N__42484;
    wire N__42483;
    wire N__42480;
    wire N__42477;
    wire N__42476;
    wire N__42471;
    wire N__42468;
    wire N__42465;
    wire N__42460;
    wire N__42457;
    wire N__42456;
    wire N__42453;
    wire N__42450;
    wire N__42449;
    wire N__42444;
    wire N__42441;
    wire N__42438;
    wire N__42433;
    wire N__42430;
    wire N__42429;
    wire N__42426;
    wire N__42425;
    wire N__42422;
    wire N__42419;
    wire N__42416;
    wire N__42411;
    wire N__42406;
    wire N__42403;
    wire N__42402;
    wire N__42399;
    wire N__42396;
    wire N__42393;
    wire N__42392;
    wire N__42387;
    wire N__42384;
    wire N__42381;
    wire N__42376;
    wire N__42373;
    wire N__42372;
    wire N__42369;
    wire N__42366;
    wire N__42365;
    wire N__42360;
    wire N__42357;
    wire N__42354;
    wire N__42349;
    wire N__42346;
    wire N__42345;
    wire N__42342;
    wire N__42339;
    wire N__42338;
    wire N__42333;
    wire N__42330;
    wire N__42327;
    wire N__42322;
    wire N__42319;
    wire N__42318;
    wire N__42315;
    wire N__42312;
    wire N__42309;
    wire N__42304;
    wire N__42301;
    wire N__42300;
    wire N__42295;
    wire N__42294;
    wire N__42291;
    wire N__42288;
    wire N__42285;
    wire N__42280;
    wire N__42277;
    wire N__42276;
    wire N__42275;
    wire N__42270;
    wire N__42267;
    wire N__42264;
    wire N__42259;
    wire N__42256;
    wire N__42255;
    wire N__42252;
    wire N__42249;
    wire N__42248;
    wire N__42243;
    wire N__42240;
    wire N__42237;
    wire N__42232;
    wire N__42229;
    wire N__42228;
    wire N__42225;
    wire N__42222;
    wire N__42221;
    wire N__42216;
    wire N__42213;
    wire N__42210;
    wire N__42205;
    wire N__42202;
    wire N__42201;
    wire N__42198;
    wire N__42195;
    wire N__42192;
    wire N__42191;
    wire N__42186;
    wire N__42183;
    wire N__42180;
    wire N__42175;
    wire N__42172;
    wire N__42171;
    wire N__42168;
    wire N__42167;
    wire N__42164;
    wire N__42161;
    wire N__42158;
    wire N__42153;
    wire N__42148;
    wire N__42145;
    wire N__42144;
    wire N__42141;
    wire N__42138;
    wire N__42137;
    wire N__42132;
    wire N__42129;
    wire N__42126;
    wire N__42121;
    wire N__42118;
    wire N__42117;
    wire N__42114;
    wire N__42111;
    wire N__42110;
    wire N__42105;
    wire N__42102;
    wire N__42099;
    wire N__42094;
    wire N__42091;
    wire N__42090;
    wire N__42087;
    wire N__42084;
    wire N__42083;
    wire N__42078;
    wire N__42075;
    wire N__42072;
    wire N__42067;
    wire N__42064;
    wire N__42063;
    wire N__42062;
    wire N__42057;
    wire N__42054;
    wire N__42051;
    wire N__42046;
    wire N__42043;
    wire N__42042;
    wire N__42037;
    wire N__42036;
    wire N__42033;
    wire N__42030;
    wire N__42027;
    wire N__42022;
    wire N__42019;
    wire N__42018;
    wire N__42015;
    wire N__42012;
    wire N__42011;
    wire N__42006;
    wire N__42003;
    wire N__42000;
    wire N__41995;
    wire N__41992;
    wire N__41991;
    wire N__41988;
    wire N__41985;
    wire N__41984;
    wire N__41979;
    wire N__41976;
    wire N__41973;
    wire N__41968;
    wire N__41965;
    wire N__41964;
    wire N__41961;
    wire N__41960;
    wire N__41957;
    wire N__41954;
    wire N__41951;
    wire N__41946;
    wire N__41941;
    wire N__41938;
    wire N__41937;
    wire N__41934;
    wire N__41931;
    wire N__41928;
    wire N__41927;
    wire N__41922;
    wire N__41919;
    wire N__41916;
    wire N__41911;
    wire N__41908;
    wire N__41907;
    wire N__41904;
    wire N__41901;
    wire N__41900;
    wire N__41895;
    wire N__41892;
    wire N__41889;
    wire N__41884;
    wire N__41881;
    wire N__41880;
    wire N__41877;
    wire N__41874;
    wire N__41873;
    wire N__41868;
    wire N__41865;
    wire N__41862;
    wire N__41857;
    wire N__41854;
    wire N__41851;
    wire N__41848;
    wire N__41845;
    wire N__41842;
    wire N__41841;
    wire N__41838;
    wire N__41835;
    wire N__41832;
    wire N__41829;
    wire N__41828;
    wire N__41825;
    wire N__41822;
    wire N__41819;
    wire N__41812;
    wire N__41809;
    wire N__41806;
    wire N__41803;
    wire N__41800;
    wire N__41799;
    wire N__41796;
    wire N__41793;
    wire N__41790;
    wire N__41789;
    wire N__41786;
    wire N__41783;
    wire N__41780;
    wire N__41779;
    wire N__41778;
    wire N__41775;
    wire N__41770;
    wire N__41767;
    wire N__41764;
    wire N__41757;
    wire N__41754;
    wire N__41751;
    wire N__41746;
    wire N__41743;
    wire N__41740;
    wire N__41739;
    wire N__41736;
    wire N__41733;
    wire N__41730;
    wire N__41729;
    wire N__41728;
    wire N__41725;
    wire N__41722;
    wire N__41719;
    wire N__41718;
    wire N__41715;
    wire N__41712;
    wire N__41709;
    wire N__41706;
    wire N__41703;
    wire N__41700;
    wire N__41691;
    wire N__41688;
    wire N__41685;
    wire N__41680;
    wire N__41677;
    wire N__41674;
    wire N__41671;
    wire N__41670;
    wire N__41667;
    wire N__41664;
    wire N__41663;
    wire N__41662;
    wire N__41659;
    wire N__41656;
    wire N__41651;
    wire N__41644;
    wire N__41641;
    wire N__41640;
    wire N__41637;
    wire N__41634;
    wire N__41629;
    wire N__41626;
    wire N__41623;
    wire N__41620;
    wire N__41617;
    wire N__41614;
    wire N__41611;
    wire N__41610;
    wire N__41607;
    wire N__41604;
    wire N__41603;
    wire N__41598;
    wire N__41595;
    wire N__41592;
    wire N__41587;
    wire N__41584;
    wire N__41581;
    wire N__41578;
    wire N__41575;
    wire N__41572;
    wire N__41571;
    wire N__41568;
    wire N__41565;
    wire N__41562;
    wire N__41559;
    wire N__41558;
    wire N__41555;
    wire N__41552;
    wire N__41549;
    wire N__41542;
    wire N__41539;
    wire N__41536;
    wire N__41533;
    wire N__41530;
    wire N__41527;
    wire N__41524;
    wire N__41523;
    wire N__41520;
    wire N__41519;
    wire N__41516;
    wire N__41515;
    wire N__41514;
    wire N__41509;
    wire N__41506;
    wire N__41501;
    wire N__41498;
    wire N__41495;
    wire N__41492;
    wire N__41489;
    wire N__41482;
    wire N__41479;
    wire N__41476;
    wire N__41473;
    wire N__41470;
    wire N__41467;
    wire N__41464;
    wire N__41461;
    wire N__41458;
    wire N__41455;
    wire N__41454;
    wire N__41453;
    wire N__41450;
    wire N__41447;
    wire N__41446;
    wire N__41443;
    wire N__41438;
    wire N__41435;
    wire N__41432;
    wire N__41429;
    wire N__41428;
    wire N__41425;
    wire N__41420;
    wire N__41417;
    wire N__41410;
    wire N__41407;
    wire N__41404;
    wire N__41401;
    wire N__41398;
    wire N__41395;
    wire N__41392;
    wire N__41391;
    wire N__41390;
    wire N__41387;
    wire N__41382;
    wire N__41379;
    wire N__41376;
    wire N__41373;
    wire N__41370;
    wire N__41365;
    wire N__41362;
    wire N__41359;
    wire N__41356;
    wire N__41353;
    wire N__41350;
    wire N__41347;
    wire N__41344;
    wire N__41341;
    wire N__41340;
    wire N__41339;
    wire N__41338;
    wire N__41335;
    wire N__41332;
    wire N__41329;
    wire N__41326;
    wire N__41323;
    wire N__41320;
    wire N__41319;
    wire N__41316;
    wire N__41313;
    wire N__41308;
    wire N__41305;
    wire N__41302;
    wire N__41299;
    wire N__41294;
    wire N__41291;
    wire N__41284;
    wire N__41281;
    wire N__41278;
    wire N__41275;
    wire N__41272;
    wire N__41269;
    wire N__41266;
    wire N__41263;
    wire N__41260;
    wire N__41257;
    wire N__41256;
    wire N__41253;
    wire N__41250;
    wire N__41245;
    wire N__41244;
    wire N__41241;
    wire N__41238;
    wire N__41233;
    wire N__41232;
    wire N__41229;
    wire N__41226;
    wire N__41221;
    wire N__41220;
    wire N__41219;
    wire N__41216;
    wire N__41215;
    wire N__41214;
    wire N__41213;
    wire N__41212;
    wire N__41211;
    wire N__41210;
    wire N__41209;
    wire N__41208;
    wire N__41207;
    wire N__41204;
    wire N__41203;
    wire N__41200;
    wire N__41199;
    wire N__41198;
    wire N__41197;
    wire N__41196;
    wire N__41195;
    wire N__41188;
    wire N__41187;
    wire N__41186;
    wire N__41185;
    wire N__41184;
    wire N__41183;
    wire N__41180;
    wire N__41177;
    wire N__41174;
    wire N__41171;
    wire N__41170;
    wire N__41169;
    wire N__41166;
    wire N__41163;
    wire N__41160;
    wire N__41159;
    wire N__41158;
    wire N__41157;
    wire N__41156;
    wire N__41155;
    wire N__41154;
    wire N__41153;
    wire N__41150;
    wire N__41143;
    wire N__41134;
    wire N__41131;
    wire N__41128;
    wire N__41119;
    wire N__41114;
    wire N__41105;
    wire N__41094;
    wire N__41083;
    wire N__41074;
    wire N__41071;
    wire N__41068;
    wire N__41065;
    wire N__41050;
    wire N__41049;
    wire N__41048;
    wire N__41047;
    wire N__41046;
    wire N__41043;
    wire N__41042;
    wire N__41041;
    wire N__41040;
    wire N__41039;
    wire N__41038;
    wire N__41037;
    wire N__41036;
    wire N__41035;
    wire N__41034;
    wire N__41033;
    wire N__41032;
    wire N__41025;
    wire N__41022;
    wire N__41021;
    wire N__41020;
    wire N__41019;
    wire N__41018;
    wire N__41017;
    wire N__41016;
    wire N__41015;
    wire N__41014;
    wire N__41013;
    wire N__41012;
    wire N__41009;
    wire N__41002;
    wire N__40993;
    wire N__40984;
    wire N__40983;
    wire N__40982;
    wire N__40981;
    wire N__40980;
    wire N__40979;
    wire N__40978;
    wire N__40975;
    wire N__40972;
    wire N__40959;
    wire N__40950;
    wire N__40947;
    wire N__40944;
    wire N__40939;
    wire N__40936;
    wire N__40925;
    wire N__40916;
    wire N__40903;
    wire N__40902;
    wire N__40899;
    wire N__40896;
    wire N__40891;
    wire N__40888;
    wire N__40885;
    wire N__40882;
    wire N__40881;
    wire N__40878;
    wire N__40877;
    wire N__40874;
    wire N__40873;
    wire N__40870;
    wire N__40867;
    wire N__40864;
    wire N__40861;
    wire N__40858;
    wire N__40855;
    wire N__40854;
    wire N__40851;
    wire N__40844;
    wire N__40841;
    wire N__40838;
    wire N__40833;
    wire N__40828;
    wire N__40825;
    wire N__40822;
    wire N__40819;
    wire N__40816;
    wire N__40813;
    wire N__40810;
    wire N__40807;
    wire N__40804;
    wire N__40801;
    wire N__40798;
    wire N__40795;
    wire N__40792;
    wire N__40789;
    wire N__40786;
    wire N__40783;
    wire N__40780;
    wire N__40777;
    wire N__40776;
    wire N__40773;
    wire N__40770;
    wire N__40765;
    wire N__40762;
    wire N__40759;
    wire N__40756;
    wire N__40753;
    wire N__40750;
    wire N__40747;
    wire N__40744;
    wire N__40741;
    wire N__40738;
    wire N__40735;
    wire N__40732;
    wire N__40729;
    wire N__40726;
    wire N__40723;
    wire N__40720;
    wire N__40717;
    wire N__40714;
    wire N__40711;
    wire N__40708;
    wire N__40705;
    wire N__40702;
    wire N__40699;
    wire N__40696;
    wire N__40693;
    wire N__40690;
    wire N__40687;
    wire N__40684;
    wire N__40681;
    wire N__40678;
    wire N__40675;
    wire N__40672;
    wire N__40669;
    wire N__40666;
    wire N__40663;
    wire N__40660;
    wire N__40657;
    wire N__40654;
    wire N__40651;
    wire N__40648;
    wire N__40645;
    wire N__40642;
    wire N__40639;
    wire N__40636;
    wire N__40633;
    wire N__40630;
    wire N__40627;
    wire N__40624;
    wire N__40621;
    wire N__40618;
    wire N__40615;
    wire N__40612;
    wire N__40609;
    wire N__40606;
    wire N__40603;
    wire N__40600;
    wire N__40597;
    wire N__40594;
    wire N__40591;
    wire N__40588;
    wire N__40585;
    wire N__40582;
    wire N__40579;
    wire N__40576;
    wire N__40573;
    wire N__40570;
    wire N__40567;
    wire N__40564;
    wire N__40561;
    wire N__40558;
    wire N__40555;
    wire N__40552;
    wire N__40549;
    wire N__40546;
    wire N__40543;
    wire N__40540;
    wire N__40537;
    wire N__40534;
    wire N__40531;
    wire N__40528;
    wire N__40525;
    wire N__40522;
    wire N__40519;
    wire N__40516;
    wire N__40513;
    wire N__40510;
    wire N__40507;
    wire N__40504;
    wire N__40501;
    wire N__40498;
    wire N__40495;
    wire N__40492;
    wire N__40489;
    wire N__40486;
    wire N__40483;
    wire N__40480;
    wire N__40477;
    wire N__40474;
    wire N__40471;
    wire N__40468;
    wire N__40465;
    wire N__40462;
    wire N__40459;
    wire N__40456;
    wire N__40453;
    wire N__40450;
    wire N__40447;
    wire N__40444;
    wire N__40441;
    wire N__40438;
    wire N__40435;
    wire N__40432;
    wire N__40429;
    wire N__40426;
    wire N__40425;
    wire N__40424;
    wire N__40421;
    wire N__40418;
    wire N__40417;
    wire N__40412;
    wire N__40409;
    wire N__40406;
    wire N__40403;
    wire N__40400;
    wire N__40397;
    wire N__40392;
    wire N__40387;
    wire N__40384;
    wire N__40381;
    wire N__40378;
    wire N__40375;
    wire N__40374;
    wire N__40373;
    wire N__40372;
    wire N__40365;
    wire N__40362;
    wire N__40357;
    wire N__40354;
    wire N__40351;
    wire N__40348;
    wire N__40345;
    wire N__40342;
    wire N__40339;
    wire N__40336;
    wire N__40333;
    wire N__40330;
    wire N__40327;
    wire N__40326;
    wire N__40325;
    wire N__40322;
    wire N__40319;
    wire N__40316;
    wire N__40313;
    wire N__40310;
    wire N__40307;
    wire N__40300;
    wire N__40297;
    wire N__40294;
    wire N__40291;
    wire N__40288;
    wire N__40285;
    wire N__40282;
    wire N__40279;
    wire N__40276;
    wire N__40273;
    wire N__40270;
    wire N__40269;
    wire N__40266;
    wire N__40263;
    wire N__40260;
    wire N__40259;
    wire N__40258;
    wire N__40255;
    wire N__40252;
    wire N__40249;
    wire N__40246;
    wire N__40241;
    wire N__40240;
    wire N__40237;
    wire N__40234;
    wire N__40231;
    wire N__40228;
    wire N__40225;
    wire N__40216;
    wire N__40213;
    wire N__40210;
    wire N__40207;
    wire N__40206;
    wire N__40205;
    wire N__40202;
    wire N__40199;
    wire N__40196;
    wire N__40195;
    wire N__40192;
    wire N__40189;
    wire N__40186;
    wire N__40183;
    wire N__40182;
    wire N__40179;
    wire N__40172;
    wire N__40169;
    wire N__40164;
    wire N__40159;
    wire N__40156;
    wire N__40153;
    wire N__40150;
    wire N__40149;
    wire N__40146;
    wire N__40143;
    wire N__40142;
    wire N__40141;
    wire N__40138;
    wire N__40135;
    wire N__40132;
    wire N__40129;
    wire N__40126;
    wire N__40123;
    wire N__40118;
    wire N__40117;
    wire N__40114;
    wire N__40109;
    wire N__40106;
    wire N__40099;
    wire N__40096;
    wire N__40093;
    wire N__40090;
    wire N__40087;
    wire N__40084;
    wire N__40081;
    wire N__40078;
    wire N__40075;
    wire N__40072;
    wire N__40069;
    wire N__40066;
    wire N__40063;
    wire N__40060;
    wire N__40057;
    wire N__40054;
    wire N__40051;
    wire N__40048;
    wire N__40045;
    wire N__40042;
    wire N__40039;
    wire N__40036;
    wire N__40033;
    wire N__40030;
    wire N__40027;
    wire N__40024;
    wire N__40021;
    wire N__40018;
    wire N__40015;
    wire N__40012;
    wire N__40009;
    wire N__40006;
    wire N__40003;
    wire N__40000;
    wire N__39997;
    wire N__39996;
    wire N__39993;
    wire N__39990;
    wire N__39989;
    wire N__39986;
    wire N__39985;
    wire N__39982;
    wire N__39979;
    wire N__39976;
    wire N__39973;
    wire N__39970;
    wire N__39963;
    wire N__39958;
    wire N__39955;
    wire N__39952;
    wire N__39949;
    wire N__39946;
    wire N__39943;
    wire N__39940;
    wire N__39939;
    wire N__39936;
    wire N__39935;
    wire N__39928;
    wire N__39925;
    wire N__39922;
    wire N__39919;
    wire N__39916;
    wire N__39913;
    wire N__39910;
    wire N__39907;
    wire N__39904;
    wire N__39901;
    wire N__39898;
    wire N__39895;
    wire N__39892;
    wire N__39889;
    wire N__39886;
    wire N__39883;
    wire N__39880;
    wire N__39877;
    wire N__39874;
    wire N__39871;
    wire N__39868;
    wire N__39865;
    wire N__39862;
    wire N__39859;
    wire N__39856;
    wire N__39853;
    wire N__39850;
    wire N__39847;
    wire N__39844;
    wire N__39841;
    wire N__39838;
    wire N__39835;
    wire N__39832;
    wire N__39829;
    wire N__39826;
    wire N__39823;
    wire N__39820;
    wire N__39817;
    wire N__39814;
    wire N__39811;
    wire N__39808;
    wire N__39805;
    wire N__39802;
    wire N__39799;
    wire N__39796;
    wire N__39793;
    wire N__39790;
    wire N__39787;
    wire N__39784;
    wire N__39781;
    wire N__39778;
    wire N__39775;
    wire N__39772;
    wire N__39769;
    wire N__39766;
    wire N__39763;
    wire N__39760;
    wire N__39757;
    wire N__39754;
    wire N__39751;
    wire N__39748;
    wire N__39745;
    wire N__39742;
    wire N__39739;
    wire N__39736;
    wire N__39733;
    wire N__39730;
    wire N__39727;
    wire N__39724;
    wire N__39721;
    wire N__39718;
    wire N__39715;
    wire N__39712;
    wire N__39709;
    wire N__39706;
    wire N__39703;
    wire N__39700;
    wire N__39697;
    wire N__39694;
    wire N__39691;
    wire N__39688;
    wire N__39685;
    wire N__39682;
    wire N__39679;
    wire N__39676;
    wire N__39673;
    wire N__39670;
    wire N__39667;
    wire N__39664;
    wire N__39661;
    wire N__39658;
    wire N__39655;
    wire N__39652;
    wire N__39649;
    wire N__39646;
    wire N__39643;
    wire N__39640;
    wire N__39637;
    wire N__39634;
    wire N__39631;
    wire N__39628;
    wire N__39625;
    wire N__39622;
    wire N__39619;
    wire N__39616;
    wire N__39613;
    wire N__39610;
    wire N__39607;
    wire N__39604;
    wire N__39601;
    wire N__39598;
    wire N__39595;
    wire N__39592;
    wire N__39589;
    wire N__39586;
    wire N__39583;
    wire N__39580;
    wire N__39577;
    wire N__39574;
    wire N__39571;
    wire N__39568;
    wire N__39565;
    wire N__39562;
    wire N__39559;
    wire N__39556;
    wire N__39553;
    wire N__39550;
    wire N__39547;
    wire N__39544;
    wire N__39541;
    wire N__39538;
    wire N__39535;
    wire N__39532;
    wire N__39529;
    wire N__39526;
    wire N__39523;
    wire N__39520;
    wire N__39517;
    wire N__39514;
    wire N__39511;
    wire N__39508;
    wire N__39505;
    wire N__39502;
    wire N__39499;
    wire N__39496;
    wire N__39493;
    wire N__39492;
    wire N__39491;
    wire N__39488;
    wire N__39485;
    wire N__39482;
    wire N__39479;
    wire N__39478;
    wire N__39475;
    wire N__39472;
    wire N__39469;
    wire N__39466;
    wire N__39465;
    wire N__39462;
    wire N__39455;
    wire N__39452;
    wire N__39449;
    wire N__39446;
    wire N__39443;
    wire N__39436;
    wire N__39433;
    wire N__39432;
    wire N__39429;
    wire N__39426;
    wire N__39425;
    wire N__39422;
    wire N__39419;
    wire N__39416;
    wire N__39413;
    wire N__39408;
    wire N__39403;
    wire N__39402;
    wire N__39399;
    wire N__39396;
    wire N__39393;
    wire N__39392;
    wire N__39389;
    wire N__39386;
    wire N__39383;
    wire N__39378;
    wire N__39377;
    wire N__39374;
    wire N__39371;
    wire N__39368;
    wire N__39361;
    wire N__39360;
    wire N__39357;
    wire N__39354;
    wire N__39353;
    wire N__39350;
    wire N__39347;
    wire N__39344;
    wire N__39343;
    wire N__39338;
    wire N__39335;
    wire N__39332;
    wire N__39331;
    wire N__39328;
    wire N__39325;
    wire N__39322;
    wire N__39319;
    wire N__39310;
    wire N__39309;
    wire N__39306;
    wire N__39303;
    wire N__39300;
    wire N__39297;
    wire N__39292;
    wire N__39289;
    wire N__39286;
    wire N__39285;
    wire N__39282;
    wire N__39279;
    wire N__39276;
    wire N__39273;
    wire N__39268;
    wire N__39265;
    wire N__39262;
    wire N__39259;
    wire N__39256;
    wire N__39253;
    wire N__39250;
    wire N__39247;
    wire N__39244;
    wire N__39241;
    wire N__39238;
    wire N__39235;
    wire N__39232;
    wire N__39229;
    wire N__39226;
    wire N__39223;
    wire N__39220;
    wire N__39217;
    wire N__39214;
    wire N__39211;
    wire N__39208;
    wire N__39207;
    wire N__39206;
    wire N__39203;
    wire N__39200;
    wire N__39197;
    wire N__39190;
    wire N__39189;
    wire N__39188;
    wire N__39187;
    wire N__39182;
    wire N__39179;
    wire N__39176;
    wire N__39169;
    wire N__39168;
    wire N__39167;
    wire N__39164;
    wire N__39161;
    wire N__39158;
    wire N__39151;
    wire N__39150;
    wire N__39147;
    wire N__39144;
    wire N__39139;
    wire N__39138;
    wire N__39135;
    wire N__39134;
    wire N__39131;
    wire N__39128;
    wire N__39125;
    wire N__39118;
    wire N__39117;
    wire N__39116;
    wire N__39115;
    wire N__39112;
    wire N__39107;
    wire N__39104;
    wire N__39097;
    wire N__39094;
    wire N__39091;
    wire N__39088;
    wire N__39085;
    wire N__39082;
    wire N__39079;
    wire N__39076;
    wire N__39073;
    wire N__39070;
    wire N__39067;
    wire N__39064;
    wire N__39061;
    wire N__39058;
    wire N__39055;
    wire N__39052;
    wire N__39049;
    wire N__39048;
    wire N__39047;
    wire N__39044;
    wire N__39041;
    wire N__39038;
    wire N__39035;
    wire N__39032;
    wire N__39029;
    wire N__39022;
    wire N__39019;
    wire N__39018;
    wire N__39017;
    wire N__39014;
    wire N__39011;
    wire N__39008;
    wire N__39005;
    wire N__39002;
    wire N__38999;
    wire N__38992;
    wire N__38991;
    wire N__38988;
    wire N__38985;
    wire N__38982;
    wire N__38979;
    wire N__38978;
    wire N__38975;
    wire N__38972;
    wire N__38969;
    wire N__38962;
    wire N__38961;
    wire N__38960;
    wire N__38957;
    wire N__38954;
    wire N__38951;
    wire N__38948;
    wire N__38945;
    wire N__38940;
    wire N__38935;
    wire N__38934;
    wire N__38931;
    wire N__38928;
    wire N__38925;
    wire N__38922;
    wire N__38919;
    wire N__38916;
    wire N__38911;
    wire N__38908;
    wire N__38905;
    wire N__38904;
    wire N__38901;
    wire N__38898;
    wire N__38897;
    wire N__38894;
    wire N__38891;
    wire N__38888;
    wire N__38881;
    wire N__38878;
    wire N__38877;
    wire N__38874;
    wire N__38871;
    wire N__38866;
    wire N__38863;
    wire N__38860;
    wire N__38859;
    wire N__38856;
    wire N__38853;
    wire N__38852;
    wire N__38849;
    wire N__38846;
    wire N__38843;
    wire N__38836;
    wire N__38833;
    wire N__38832;
    wire N__38831;
    wire N__38828;
    wire N__38825;
    wire N__38822;
    wire N__38817;
    wire N__38812;
    wire N__38811;
    wire N__38810;
    wire N__38809;
    wire N__38808;
    wire N__38797;
    wire N__38794;
    wire N__38791;
    wire N__38788;
    wire N__38785;
    wire N__38782;
    wire N__38779;
    wire N__38778;
    wire N__38777;
    wire N__38776;
    wire N__38773;
    wire N__38770;
    wire N__38767;
    wire N__38764;
    wire N__38757;
    wire N__38754;
    wire N__38751;
    wire N__38748;
    wire N__38745;
    wire N__38742;
    wire N__38737;
    wire N__38734;
    wire N__38731;
    wire N__38728;
    wire N__38725;
    wire N__38722;
    wire N__38719;
    wire N__38716;
    wire N__38713;
    wire N__38710;
    wire N__38707;
    wire N__38704;
    wire N__38701;
    wire N__38698;
    wire N__38695;
    wire N__38692;
    wire N__38689;
    wire N__38686;
    wire N__38683;
    wire N__38680;
    wire N__38677;
    wire N__38674;
    wire N__38671;
    wire N__38668;
    wire N__38665;
    wire N__38662;
    wire N__38659;
    wire N__38656;
    wire N__38653;
    wire N__38650;
    wire N__38647;
    wire N__38644;
    wire N__38641;
    wire N__38638;
    wire N__38635;
    wire N__38632;
    wire N__38629;
    wire N__38626;
    wire N__38623;
    wire N__38620;
    wire N__38617;
    wire N__38614;
    wire N__38611;
    wire N__38608;
    wire N__38605;
    wire N__38602;
    wire N__38599;
    wire N__38596;
    wire N__38593;
    wire N__38590;
    wire N__38587;
    wire N__38584;
    wire N__38581;
    wire N__38578;
    wire N__38575;
    wire N__38572;
    wire N__38569;
    wire N__38566;
    wire N__38563;
    wire N__38560;
    wire N__38557;
    wire N__38554;
    wire N__38551;
    wire N__38548;
    wire N__38545;
    wire N__38542;
    wire N__38539;
    wire N__38536;
    wire N__38533;
    wire N__38530;
    wire N__38527;
    wire N__38524;
    wire N__38521;
    wire N__38518;
    wire N__38515;
    wire N__38512;
    wire N__38509;
    wire N__38506;
    wire N__38503;
    wire N__38500;
    wire N__38497;
    wire N__38494;
    wire N__38491;
    wire N__38488;
    wire N__38485;
    wire N__38482;
    wire N__38479;
    wire N__38476;
    wire N__38473;
    wire N__38470;
    wire N__38467;
    wire N__38464;
    wire N__38461;
    wire N__38458;
    wire N__38455;
    wire N__38452;
    wire N__38449;
    wire N__38446;
    wire N__38443;
    wire N__38440;
    wire N__38437;
    wire N__38434;
    wire N__38431;
    wire N__38428;
    wire N__38425;
    wire N__38422;
    wire N__38419;
    wire N__38416;
    wire N__38413;
    wire N__38410;
    wire N__38407;
    wire N__38404;
    wire N__38401;
    wire N__38398;
    wire N__38395;
    wire N__38394;
    wire N__38393;
    wire N__38392;
    wire N__38391;
    wire N__38390;
    wire N__38389;
    wire N__38388;
    wire N__38387;
    wire N__38386;
    wire N__38385;
    wire N__38384;
    wire N__38383;
    wire N__38382;
    wire N__38381;
    wire N__38380;
    wire N__38379;
    wire N__38378;
    wire N__38377;
    wire N__38376;
    wire N__38375;
    wire N__38374;
    wire N__38373;
    wire N__38372;
    wire N__38369;
    wire N__38368;
    wire N__38367;
    wire N__38366;
    wire N__38365;
    wire N__38364;
    wire N__38363;
    wire N__38362;
    wire N__38355;
    wire N__38346;
    wire N__38343;
    wire N__38340;
    wire N__38339;
    wire N__38336;
    wire N__38333;
    wire N__38330;
    wire N__38327;
    wire N__38326;
    wire N__38323;
    wire N__38320;
    wire N__38317;
    wire N__38314;
    wire N__38311;
    wire N__38308;
    wire N__38305;
    wire N__38302;
    wire N__38299;
    wire N__38296;
    wire N__38295;
    wire N__38294;
    wire N__38293;
    wire N__38292;
    wire N__38291;
    wire N__38290;
    wire N__38289;
    wire N__38288;
    wire N__38287;
    wire N__38286;
    wire N__38285;
    wire N__38284;
    wire N__38283;
    wire N__38282;
    wire N__38281;
    wire N__38280;
    wire N__38279;
    wire N__38276;
    wire N__38269;
    wire N__38260;
    wire N__38255;
    wire N__38252;
    wire N__38247;
    wire N__38242;
    wire N__38231;
    wire N__38222;
    wire N__38213;
    wire N__38210;
    wire N__38207;
    wire N__38204;
    wire N__38201;
    wire N__38200;
    wire N__38197;
    wire N__38194;
    wire N__38191;
    wire N__38188;
    wire N__38185;
    wire N__38182;
    wire N__38179;
    wire N__38176;
    wire N__38173;
    wire N__38170;
    wire N__38167;
    wire N__38164;
    wire N__38163;
    wire N__38162;
    wire N__38159;
    wire N__38156;
    wire N__38151;
    wire N__38148;
    wire N__38143;
    wire N__38134;
    wire N__38127;
    wire N__38116;
    wire N__38113;
    wire N__38110;
    wire N__38103;
    wire N__38094;
    wire N__38091;
    wire N__38088;
    wire N__38087;
    wire N__38086;
    wire N__38083;
    wire N__38078;
    wire N__38073;
    wire N__38070;
    wire N__38065;
    wire N__38060;
    wire N__38055;
    wire N__38052;
    wire N__38049;
    wire N__38046;
    wire N__38043;
    wire N__38038;
    wire N__38035;
    wire N__38028;
    wire N__38023;
    wire N__38020;
    wire N__38015;
    wire N__38012;
    wire N__38001;
    wire N__37996;
    wire N__37993;
    wire N__37992;
    wire N__37989;
    wire N__37986;
    wire N__37983;
    wire N__37978;
    wire N__37975;
    wire N__37974;
    wire N__37971;
    wire N__37968;
    wire N__37965;
    wire N__37962;
    wire N__37959;
    wire N__37956;
    wire N__37951;
    wire N__37948;
    wire N__37945;
    wire N__37942;
    wire N__37939;
    wire N__37936;
    wire N__37935;
    wire N__37934;
    wire N__37933;
    wire N__37932;
    wire N__37931;
    wire N__37928;
    wire N__37927;
    wire N__37926;
    wire N__37923;
    wire N__37916;
    wire N__37913;
    wire N__37912;
    wire N__37911;
    wire N__37910;
    wire N__37909;
    wire N__37908;
    wire N__37905;
    wire N__37900;
    wire N__37897;
    wire N__37894;
    wire N__37881;
    wire N__37878;
    wire N__37873;
    wire N__37870;
    wire N__37867;
    wire N__37864;
    wire N__37861;
    wire N__37852;
    wire N__37849;
    wire N__37846;
    wire N__37845;
    wire N__37844;
    wire N__37843;
    wire N__37840;
    wire N__37837;
    wire N__37832;
    wire N__37827;
    wire N__37822;
    wire N__37819;
    wire N__37816;
    wire N__37813;
    wire N__37810;
    wire N__37807;
    wire N__37804;
    wire N__37801;
    wire N__37798;
    wire N__37795;
    wire N__37792;
    wire N__37789;
    wire N__37786;
    wire N__37783;
    wire N__37780;
    wire N__37777;
    wire N__37774;
    wire N__37771;
    wire N__37768;
    wire N__37765;
    wire N__37762;
    wire N__37759;
    wire N__37756;
    wire N__37753;
    wire N__37750;
    wire N__37747;
    wire N__37744;
    wire N__37741;
    wire N__37738;
    wire N__37737;
    wire N__37736;
    wire N__37733;
    wire N__37732;
    wire N__37731;
    wire N__37728;
    wire N__37725;
    wire N__37722;
    wire N__37717;
    wire N__37712;
    wire N__37705;
    wire N__37702;
    wire N__37699;
    wire N__37696;
    wire N__37695;
    wire N__37694;
    wire N__37693;
    wire N__37692;
    wire N__37687;
    wire N__37686;
    wire N__37683;
    wire N__37680;
    wire N__37677;
    wire N__37674;
    wire N__37669;
    wire N__37660;
    wire N__37657;
    wire N__37654;
    wire N__37651;
    wire N__37648;
    wire N__37647;
    wire N__37646;
    wire N__37643;
    wire N__37640;
    wire N__37637;
    wire N__37634;
    wire N__37629;
    wire N__37626;
    wire N__37623;
    wire N__37618;
    wire N__37615;
    wire N__37614;
    wire N__37611;
    wire N__37610;
    wire N__37607;
    wire N__37604;
    wire N__37601;
    wire N__37598;
    wire N__37595;
    wire N__37592;
    wire N__37589;
    wire N__37586;
    wire N__37583;
    wire N__37576;
    wire N__37573;
    wire N__37572;
    wire N__37571;
    wire N__37568;
    wire N__37565;
    wire N__37562;
    wire N__37559;
    wire N__37556;
    wire N__37553;
    wire N__37550;
    wire N__37547;
    wire N__37544;
    wire N__37537;
    wire N__37534;
    wire N__37533;
    wire N__37532;
    wire N__37529;
    wire N__37526;
    wire N__37523;
    wire N__37520;
    wire N__37517;
    wire N__37514;
    wire N__37511;
    wire N__37508;
    wire N__37505;
    wire N__37498;
    wire N__37495;
    wire N__37492;
    wire N__37489;
    wire N__37486;
    wire N__37485;
    wire N__37484;
    wire N__37483;
    wire N__37482;
    wire N__37481;
    wire N__37480;
    wire N__37475;
    wire N__37474;
    wire N__37465;
    wire N__37462;
    wire N__37459;
    wire N__37456;
    wire N__37451;
    wire N__37446;
    wire N__37443;
    wire N__37440;
    wire N__37435;
    wire N__37432;
    wire N__37431;
    wire N__37428;
    wire N__37425;
    wire N__37422;
    wire N__37419;
    wire N__37416;
    wire N__37413;
    wire N__37408;
    wire N__37405;
    wire N__37404;
    wire N__37401;
    wire N__37398;
    wire N__37395;
    wire N__37392;
    wire N__37389;
    wire N__37384;
    wire N__37381;
    wire N__37380;
    wire N__37377;
    wire N__37372;
    wire N__37371;
    wire N__37370;
    wire N__37369;
    wire N__37366;
    wire N__37363;
    wire N__37360;
    wire N__37357;
    wire N__37354;
    wire N__37349;
    wire N__37346;
    wire N__37343;
    wire N__37340;
    wire N__37337;
    wire N__37330;
    wire N__37327;
    wire N__37324;
    wire N__37323;
    wire N__37320;
    wire N__37317;
    wire N__37312;
    wire N__37309;
    wire N__37306;
    wire N__37303;
    wire N__37300;
    wire N__37299;
    wire N__37296;
    wire N__37293;
    wire N__37288;
    wire N__37285;
    wire N__37282;
    wire N__37279;
    wire N__37278;
    wire N__37275;
    wire N__37272;
    wire N__37269;
    wire N__37266;
    wire N__37261;
    wire N__37258;
    wire N__37257;
    wire N__37254;
    wire N__37251;
    wire N__37248;
    wire N__37245;
    wire N__37240;
    wire N__37237;
    wire N__37234;
    wire N__37233;
    wire N__37232;
    wire N__37229;
    wire N__37226;
    wire N__37223;
    wire N__37220;
    wire N__37217;
    wire N__37210;
    wire N__37207;
    wire N__37204;
    wire N__37201;
    wire N__37200;
    wire N__37199;
    wire N__37196;
    wire N__37193;
    wire N__37190;
    wire N__37185;
    wire N__37180;
    wire N__37177;
    wire N__37174;
    wire N__37173;
    wire N__37172;
    wire N__37169;
    wire N__37166;
    wire N__37163;
    wire N__37156;
    wire N__37153;
    wire N__37150;
    wire N__37147;
    wire N__37146;
    wire N__37143;
    wire N__37140;
    wire N__37137;
    wire N__37134;
    wire N__37133;
    wire N__37128;
    wire N__37125;
    wire N__37120;
    wire N__37117;
    wire N__37116;
    wire N__37115;
    wire N__37112;
    wire N__37109;
    wire N__37106;
    wire N__37103;
    wire N__37100;
    wire N__37099;
    wire N__37098;
    wire N__37095;
    wire N__37090;
    wire N__37085;
    wire N__37082;
    wire N__37075;
    wire N__37072;
    wire N__37069;
    wire N__37066;
    wire N__37065;
    wire N__37064;
    wire N__37061;
    wire N__37058;
    wire N__37055;
    wire N__37050;
    wire N__37045;
    wire N__37042;
    wire N__37039;
    wire N__37036;
    wire N__37035;
    wire N__37032;
    wire N__37031;
    wire N__37028;
    wire N__37025;
    wire N__37022;
    wire N__37019;
    wire N__37016;
    wire N__37013;
    wire N__37010;
    wire N__37007;
    wire N__37004;
    wire N__37001;
    wire N__36994;
    wire N__36993;
    wire N__36990;
    wire N__36987;
    wire N__36982;
    wire N__36979;
    wire N__36976;
    wire N__36973;
    wire N__36972;
    wire N__36969;
    wire N__36966;
    wire N__36961;
    wire N__36958;
    wire N__36955;
    wire N__36952;
    wire N__36951;
    wire N__36950;
    wire N__36947;
    wire N__36942;
    wire N__36939;
    wire N__36936;
    wire N__36931;
    wire N__36928;
    wire N__36927;
    wire N__36924;
    wire N__36921;
    wire N__36918;
    wire N__36915;
    wire N__36912;
    wire N__36911;
    wire N__36908;
    wire N__36907;
    wire N__36906;
    wire N__36903;
    wire N__36900;
    wire N__36897;
    wire N__36894;
    wire N__36891;
    wire N__36886;
    wire N__36877;
    wire N__36874;
    wire N__36871;
    wire N__36868;
    wire N__36865;
    wire N__36862;
    wire N__36861;
    wire N__36858;
    wire N__36855;
    wire N__36854;
    wire N__36851;
    wire N__36848;
    wire N__36845;
    wire N__36840;
    wire N__36837;
    wire N__36832;
    wire N__36831;
    wire N__36828;
    wire N__36827;
    wire N__36824;
    wire N__36821;
    wire N__36820;
    wire N__36819;
    wire N__36816;
    wire N__36813;
    wire N__36810;
    wire N__36807;
    wire N__36804;
    wire N__36801;
    wire N__36796;
    wire N__36793;
    wire N__36790;
    wire N__36787;
    wire N__36778;
    wire N__36775;
    wire N__36772;
    wire N__36771;
    wire N__36768;
    wire N__36765;
    wire N__36764;
    wire N__36761;
    wire N__36758;
    wire N__36755;
    wire N__36752;
    wire N__36749;
    wire N__36746;
    wire N__36739;
    wire N__36738;
    wire N__36735;
    wire N__36732;
    wire N__36729;
    wire N__36726;
    wire N__36725;
    wire N__36722;
    wire N__36719;
    wire N__36716;
    wire N__36709;
    wire N__36706;
    wire N__36703;
    wire N__36702;
    wire N__36699;
    wire N__36696;
    wire N__36691;
    wire N__36688;
    wire N__36685;
    wire N__36682;
    wire N__36679;
    wire N__36678;
    wire N__36677;
    wire N__36674;
    wire N__36671;
    wire N__36668;
    wire N__36665;
    wire N__36660;
    wire N__36655;
    wire N__36652;
    wire N__36649;
    wire N__36646;
    wire N__36643;
    wire N__36642;
    wire N__36639;
    wire N__36638;
    wire N__36635;
    wire N__36632;
    wire N__36629;
    wire N__36626;
    wire N__36621;
    wire N__36616;
    wire N__36613;
    wire N__36610;
    wire N__36609;
    wire N__36606;
    wire N__36603;
    wire N__36602;
    wire N__36599;
    wire N__36596;
    wire N__36593;
    wire N__36590;
    wire N__36585;
    wire N__36580;
    wire N__36577;
    wire N__36574;
    wire N__36571;
    wire N__36570;
    wire N__36567;
    wire N__36564;
    wire N__36561;
    wire N__36560;
    wire N__36557;
    wire N__36554;
    wire N__36551;
    wire N__36546;
    wire N__36543;
    wire N__36538;
    wire N__36535;
    wire N__36532;
    wire N__36531;
    wire N__36530;
    wire N__36527;
    wire N__36524;
    wire N__36521;
    wire N__36518;
    wire N__36517;
    wire N__36514;
    wire N__36511;
    wire N__36508;
    wire N__36505;
    wire N__36502;
    wire N__36499;
    wire N__36492;
    wire N__36487;
    wire N__36486;
    wire N__36483;
    wire N__36480;
    wire N__36479;
    wire N__36476;
    wire N__36473;
    wire N__36470;
    wire N__36465;
    wire N__36462;
    wire N__36457;
    wire N__36454;
    wire N__36451;
    wire N__36450;
    wire N__36447;
    wire N__36444;
    wire N__36441;
    wire N__36438;
    wire N__36437;
    wire N__36434;
    wire N__36431;
    wire N__36428;
    wire N__36421;
    wire N__36418;
    wire N__36415;
    wire N__36412;
    wire N__36411;
    wire N__36410;
    wire N__36409;
    wire N__36406;
    wire N__36403;
    wire N__36400;
    wire N__36399;
    wire N__36396;
    wire N__36395;
    wire N__36392;
    wire N__36389;
    wire N__36386;
    wire N__36383;
    wire N__36380;
    wire N__36377;
    wire N__36374;
    wire N__36371;
    wire N__36366;
    wire N__36363;
    wire N__36360;
    wire N__36357;
    wire N__36354;
    wire N__36351;
    wire N__36348;
    wire N__36345;
    wire N__36342;
    wire N__36339;
    wire N__36336;
    wire N__36331;
    wire N__36322;
    wire N__36321;
    wire N__36318;
    wire N__36315;
    wire N__36312;
    wire N__36311;
    wire N__36308;
    wire N__36305;
    wire N__36302;
    wire N__36299;
    wire N__36296;
    wire N__36293;
    wire N__36286;
    wire N__36283;
    wire N__36280;
    wire N__36277;
    wire N__36276;
    wire N__36273;
    wire N__36270;
    wire N__36269;
    wire N__36266;
    wire N__36263;
    wire N__36260;
    wire N__36257;
    wire N__36252;
    wire N__36247;
    wire N__36244;
    wire N__36241;
    wire N__36240;
    wire N__36237;
    wire N__36234;
    wire N__36233;
    wire N__36230;
    wire N__36227;
    wire N__36224;
    wire N__36219;
    wire N__36216;
    wire N__36211;
    wire N__36208;
    wire N__36205;
    wire N__36204;
    wire N__36201;
    wire N__36198;
    wire N__36197;
    wire N__36194;
    wire N__36191;
    wire N__36188;
    wire N__36183;
    wire N__36180;
    wire N__36175;
    wire N__36172;
    wire N__36169;
    wire N__36168;
    wire N__36165;
    wire N__36162;
    wire N__36161;
    wire N__36158;
    wire N__36155;
    wire N__36152;
    wire N__36149;
    wire N__36144;
    wire N__36139;
    wire N__36136;
    wire N__36133;
    wire N__36132;
    wire N__36127;
    wire N__36126;
    wire N__36123;
    wire N__36120;
    wire N__36117;
    wire N__36112;
    wire N__36109;
    wire N__36106;
    wire N__36103;
    wire N__36100;
    wire N__36099;
    wire N__36096;
    wire N__36093;
    wire N__36090;
    wire N__36089;
    wire N__36084;
    wire N__36081;
    wire N__36078;
    wire N__36073;
    wire N__36070;
    wire N__36067;
    wire N__36064;
    wire N__36063;
    wire N__36060;
    wire N__36057;
    wire N__36054;
    wire N__36051;
    wire N__36050;
    wire N__36045;
    wire N__36042;
    wire N__36039;
    wire N__36034;
    wire N__36031;
    wire N__36028;
    wire N__36025;
    wire N__36024;
    wire N__36021;
    wire N__36020;
    wire N__36017;
    wire N__36014;
    wire N__36011;
    wire N__36006;
    wire N__36001;
    wire N__35998;
    wire N__35995;
    wire N__35994;
    wire N__35991;
    wire N__35988;
    wire N__35985;
    wire N__35980;
    wire N__35977;
    wire N__35974;
    wire N__35971;
    wire N__35970;
    wire N__35967;
    wire N__35966;
    wire N__35963;
    wire N__35960;
    wire N__35957;
    wire N__35952;
    wire N__35947;
    wire N__35944;
    wire N__35943;
    wire N__35940;
    wire N__35937;
    wire N__35934;
    wire N__35929;
    wire N__35926;
    wire N__35923;
    wire N__35920;
    wire N__35917;
    wire N__35914;
    wire N__35911;
    wire N__35910;
    wire N__35907;
    wire N__35904;
    wire N__35899;
    wire N__35896;
    wire N__35893;
    wire N__35890;
    wire N__35887;
    wire N__35884;
    wire N__35883;
    wire N__35878;
    wire N__35877;
    wire N__35874;
    wire N__35871;
    wire N__35868;
    wire N__35863;
    wire N__35860;
    wire N__35859;
    wire N__35856;
    wire N__35853;
    wire N__35850;
    wire N__35847;
    wire N__35846;
    wire N__35841;
    wire N__35838;
    wire N__35835;
    wire N__35830;
    wire N__35827;
    wire N__35826;
    wire N__35823;
    wire N__35820;
    wire N__35817;
    wire N__35814;
    wire N__35813;
    wire N__35808;
    wire N__35805;
    wire N__35802;
    wire N__35797;
    wire N__35796;
    wire N__35793;
    wire N__35790;
    wire N__35787;
    wire N__35782;
    wire N__35779;
    wire N__35778;
    wire N__35775;
    wire N__35774;
    wire N__35771;
    wire N__35768;
    wire N__35765;
    wire N__35760;
    wire N__35755;
    wire N__35754;
    wire N__35749;
    wire N__35746;
    wire N__35743;
    wire N__35742;
    wire N__35739;
    wire N__35738;
    wire N__35735;
    wire N__35732;
    wire N__35729;
    wire N__35724;
    wire N__35719;
    wire N__35718;
    wire N__35713;
    wire N__35710;
    wire N__35707;
    wire N__35706;
    wire N__35703;
    wire N__35700;
    wire N__35695;
    wire N__35694;
    wire N__35691;
    wire N__35688;
    wire N__35685;
    wire N__35680;
    wire N__35677;
    wire N__35674;
    wire N__35671;
    wire N__35670;
    wire N__35667;
    wire N__35664;
    wire N__35663;
    wire N__35658;
    wire N__35655;
    wire N__35652;
    wire N__35647;
    wire N__35644;
    wire N__35641;
    wire N__35638;
    wire N__35637;
    wire N__35632;
    wire N__35631;
    wire N__35628;
    wire N__35625;
    wire N__35622;
    wire N__35617;
    wire N__35614;
    wire N__35611;
    wire N__35608;
    wire N__35605;
    wire N__35604;
    wire N__35601;
    wire N__35598;
    wire N__35593;
    wire N__35592;
    wire N__35589;
    wire N__35586;
    wire N__35583;
    wire N__35578;
    wire N__35577;
    wire N__35574;
    wire N__35571;
    wire N__35568;
    wire N__35565;
    wire N__35564;
    wire N__35561;
    wire N__35558;
    wire N__35555;
    wire N__35548;
    wire N__35545;
    wire N__35544;
    wire N__35541;
    wire N__35540;
    wire N__35537;
    wire N__35534;
    wire N__35531;
    wire N__35526;
    wire N__35521;
    wire N__35518;
    wire N__35517;
    wire N__35516;
    wire N__35513;
    wire N__35510;
    wire N__35507;
    wire N__35502;
    wire N__35497;
    wire N__35494;
    wire N__35491;
    wire N__35490;
    wire N__35487;
    wire N__35484;
    wire N__35483;
    wire N__35478;
    wire N__35475;
    wire N__35472;
    wire N__35467;
    wire N__35466;
    wire N__35463;
    wire N__35460;
    wire N__35459;
    wire N__35456;
    wire N__35453;
    wire N__35450;
    wire N__35445;
    wire N__35440;
    wire N__35437;
    wire N__35436;
    wire N__35433;
    wire N__35432;
    wire N__35429;
    wire N__35426;
    wire N__35423;
    wire N__35418;
    wire N__35413;
    wire N__35412;
    wire N__35409;
    wire N__35406;
    wire N__35403;
    wire N__35402;
    wire N__35399;
    wire N__35396;
    wire N__35393;
    wire N__35390;
    wire N__35383;
    wire N__35380;
    wire N__35379;
    wire N__35376;
    wire N__35375;
    wire N__35372;
    wire N__35369;
    wire N__35366;
    wire N__35361;
    wire N__35356;
    wire N__35353;
    wire N__35350;
    wire N__35349;
    wire N__35348;
    wire N__35347;
    wire N__35344;
    wire N__35339;
    wire N__35336;
    wire N__35329;
    wire N__35326;
    wire N__35325;
    wire N__35322;
    wire N__35319;
    wire N__35314;
    wire N__35313;
    wire N__35310;
    wire N__35307;
    wire N__35304;
    wire N__35299;
    wire N__35298;
    wire N__35295;
    wire N__35294;
    wire N__35293;
    wire N__35290;
    wire N__35287;
    wire N__35284;
    wire N__35279;
    wire N__35272;
    wire N__35269;
    wire N__35268;
    wire N__35265;
    wire N__35262;
    wire N__35261;
    wire N__35256;
    wire N__35253;
    wire N__35250;
    wire N__35245;
    wire N__35242;
    wire N__35241;
    wire N__35236;
    wire N__35235;
    wire N__35232;
    wire N__35229;
    wire N__35226;
    wire N__35221;
    wire N__35218;
    wire N__35215;
    wire N__35212;
    wire N__35209;
    wire N__35206;
    wire N__35203;
    wire N__35202;
    wire N__35201;
    wire N__35198;
    wire N__35195;
    wire N__35192;
    wire N__35185;
    wire N__35184;
    wire N__35183;
    wire N__35180;
    wire N__35175;
    wire N__35170;
    wire N__35167;
    wire N__35166;
    wire N__35163;
    wire N__35162;
    wire N__35159;
    wire N__35156;
    wire N__35153;
    wire N__35148;
    wire N__35143;
    wire N__35140;
    wire N__35137;
    wire N__35136;
    wire N__35135;
    wire N__35132;
    wire N__35127;
    wire N__35122;
    wire N__35119;
    wire N__35118;
    wire N__35115;
    wire N__35114;
    wire N__35111;
    wire N__35108;
    wire N__35105;
    wire N__35100;
    wire N__35095;
    wire N__35092;
    wire N__35091;
    wire N__35090;
    wire N__35089;
    wire N__35086;
    wire N__35079;
    wire N__35074;
    wire N__35071;
    wire N__35070;
    wire N__35067;
    wire N__35064;
    wire N__35059;
    wire N__35058;
    wire N__35055;
    wire N__35052;
    wire N__35049;
    wire N__35044;
    wire N__35041;
    wire N__35040;
    wire N__35039;
    wire N__35038;
    wire N__35035;
    wire N__35032;
    wire N__35029;
    wire N__35026;
    wire N__35017;
    wire N__35014;
    wire N__35013;
    wire N__35010;
    wire N__35007;
    wire N__35004;
    wire N__35003;
    wire N__34998;
    wire N__34995;
    wire N__34992;
    wire N__34987;
    wire N__34986;
    wire N__34983;
    wire N__34982;
    wire N__34979;
    wire N__34976;
    wire N__34973;
    wire N__34972;
    wire N__34969;
    wire N__34966;
    wire N__34963;
    wire N__34960;
    wire N__34957;
    wire N__34948;
    wire N__34945;
    wire N__34944;
    wire N__34939;
    wire N__34938;
    wire N__34935;
    wire N__34932;
    wire N__34929;
    wire N__34924;
    wire N__34921;
    wire N__34920;
    wire N__34917;
    wire N__34916;
    wire N__34913;
    wire N__34912;
    wire N__34909;
    wire N__34906;
    wire N__34901;
    wire N__34894;
    wire N__34891;
    wire N__34888;
    wire N__34885;
    wire N__34882;
    wire N__34879;
    wire N__34876;
    wire N__34873;
    wire N__34870;
    wire N__34869;
    wire N__34868;
    wire N__34867;
    wire N__34866;
    wire N__34865;
    wire N__34864;
    wire N__34863;
    wire N__34862;
    wire N__34861;
    wire N__34860;
    wire N__34859;
    wire N__34858;
    wire N__34857;
    wire N__34856;
    wire N__34855;
    wire N__34854;
    wire N__34853;
    wire N__34852;
    wire N__34851;
    wire N__34850;
    wire N__34849;
    wire N__34840;
    wire N__34831;
    wire N__34826;
    wire N__34825;
    wire N__34824;
    wire N__34823;
    wire N__34822;
    wire N__34821;
    wire N__34820;
    wire N__34819;
    wire N__34818;
    wire N__34809;
    wire N__34800;
    wire N__34791;
    wire N__34784;
    wire N__34775;
    wire N__34766;
    wire N__34759;
    wire N__34756;
    wire N__34747;
    wire N__34744;
    wire N__34741;
    wire N__34740;
    wire N__34739;
    wire N__34736;
    wire N__34733;
    wire N__34730;
    wire N__34727;
    wire N__34726;
    wire N__34721;
    wire N__34718;
    wire N__34715;
    wire N__34712;
    wire N__34707;
    wire N__34702;
    wire N__34699;
    wire N__34696;
    wire N__34693;
    wire N__34690;
    wire N__34687;
    wire N__34684;
    wire N__34681;
    wire N__34678;
    wire N__34675;
    wire N__34672;
    wire N__34669;
    wire N__34666;
    wire N__34663;
    wire N__34660;
    wire N__34657;
    wire N__34654;
    wire N__34651;
    wire N__34648;
    wire N__34645;
    wire N__34642;
    wire N__34639;
    wire N__34636;
    wire N__34633;
    wire N__34630;
    wire N__34627;
    wire N__34624;
    wire N__34621;
    wire N__34618;
    wire N__34615;
    wire N__34612;
    wire N__34609;
    wire N__34606;
    wire N__34603;
    wire N__34600;
    wire N__34597;
    wire N__34594;
    wire N__34591;
    wire N__34588;
    wire N__34585;
    wire N__34582;
    wire N__34579;
    wire N__34576;
    wire N__34573;
    wire N__34570;
    wire N__34567;
    wire N__34564;
    wire N__34561;
    wire N__34558;
    wire N__34555;
    wire N__34552;
    wire N__34549;
    wire N__34546;
    wire N__34543;
    wire N__34540;
    wire N__34537;
    wire N__34534;
    wire N__34531;
    wire N__34528;
    wire N__34525;
    wire N__34522;
    wire N__34519;
    wire N__34516;
    wire N__34513;
    wire N__34510;
    wire N__34507;
    wire N__34504;
    wire N__34501;
    wire N__34498;
    wire N__34495;
    wire N__34492;
    wire N__34489;
    wire N__34486;
    wire N__34483;
    wire N__34480;
    wire N__34477;
    wire N__34474;
    wire N__34471;
    wire N__34468;
    wire N__34465;
    wire N__34462;
    wire N__34459;
    wire N__34456;
    wire N__34453;
    wire N__34450;
    wire N__34447;
    wire N__34444;
    wire N__34441;
    wire N__34438;
    wire N__34435;
    wire N__34432;
    wire N__34429;
    wire N__34426;
    wire N__34423;
    wire N__34420;
    wire N__34417;
    wire N__34414;
    wire N__34411;
    wire N__34408;
    wire N__34405;
    wire N__34402;
    wire N__34399;
    wire N__34396;
    wire N__34393;
    wire N__34390;
    wire N__34387;
    wire N__34386;
    wire N__34381;
    wire N__34378;
    wire N__34375;
    wire N__34372;
    wire N__34369;
    wire N__34366;
    wire N__34363;
    wire N__34360;
    wire N__34357;
    wire N__34356;
    wire N__34353;
    wire N__34350;
    wire N__34347;
    wire N__34342;
    wire N__34339;
    wire N__34336;
    wire N__34333;
    wire N__34330;
    wire N__34327;
    wire N__34324;
    wire N__34321;
    wire N__34318;
    wire N__34315;
    wire N__34312;
    wire N__34309;
    wire N__34306;
    wire N__34303;
    wire N__34300;
    wire N__34297;
    wire N__34294;
    wire N__34291;
    wire N__34288;
    wire N__34285;
    wire N__34282;
    wire N__34279;
    wire N__34276;
    wire N__34273;
    wire N__34270;
    wire N__34267;
    wire N__34264;
    wire N__34261;
    wire N__34258;
    wire N__34255;
    wire N__34252;
    wire N__34249;
    wire N__34246;
    wire N__34243;
    wire N__34240;
    wire N__34237;
    wire N__34234;
    wire N__34231;
    wire N__34228;
    wire N__34225;
    wire N__34222;
    wire N__34219;
    wire N__34216;
    wire N__34213;
    wire N__34210;
    wire N__34207;
    wire N__34204;
    wire N__34201;
    wire N__34198;
    wire N__34195;
    wire N__34192;
    wire N__34189;
    wire N__34186;
    wire N__34183;
    wire N__34180;
    wire N__34177;
    wire N__34174;
    wire N__34171;
    wire N__34168;
    wire N__34165;
    wire N__34162;
    wire N__34159;
    wire N__34156;
    wire N__34153;
    wire N__34150;
    wire N__34147;
    wire N__34144;
    wire N__34141;
    wire N__34138;
    wire N__34135;
    wire N__34132;
    wire N__34129;
    wire N__34126;
    wire N__34123;
    wire N__34120;
    wire N__34117;
    wire N__34114;
    wire N__34111;
    wire N__34108;
    wire N__34105;
    wire N__34102;
    wire N__34099;
    wire N__34096;
    wire N__34093;
    wire N__34090;
    wire N__34087;
    wire N__34084;
    wire N__34081;
    wire N__34078;
    wire N__34075;
    wire N__34072;
    wire N__34069;
    wire N__34066;
    wire N__34063;
    wire N__34060;
    wire N__34057;
    wire N__34054;
    wire N__34051;
    wire N__34048;
    wire N__34047;
    wire N__34046;
    wire N__34045;
    wire N__34044;
    wire N__34043;
    wire N__34042;
    wire N__34035;
    wire N__34030;
    wire N__34027;
    wire N__34026;
    wire N__34025;
    wire N__34022;
    wire N__34021;
    wire N__34016;
    wire N__34013;
    wire N__34010;
    wire N__34007;
    wire N__34004;
    wire N__34001;
    wire N__33996;
    wire N__33985;
    wire N__33984;
    wire N__33983;
    wire N__33980;
    wire N__33975;
    wire N__33972;
    wire N__33969;
    wire N__33968;
    wire N__33967;
    wire N__33966;
    wire N__33963;
    wire N__33960;
    wire N__33957;
    wire N__33952;
    wire N__33943;
    wire N__33940;
    wire N__33937;
    wire N__33934;
    wire N__33931;
    wire N__33928;
    wire N__33927;
    wire N__33926;
    wire N__33925;
    wire N__33922;
    wire N__33921;
    wire N__33918;
    wire N__33917;
    wire N__33914;
    wire N__33911;
    wire N__33908;
    wire N__33905;
    wire N__33902;
    wire N__33899;
    wire N__33896;
    wire N__33893;
    wire N__33890;
    wire N__33887;
    wire N__33884;
    wire N__33879;
    wire N__33876;
    wire N__33871;
    wire N__33862;
    wire N__33859;
    wire N__33856;
    wire N__33853;
    wire N__33850;
    wire N__33847;
    wire N__33844;
    wire N__33841;
    wire N__33838;
    wire N__33835;
    wire N__33834;
    wire N__33831;
    wire N__33828;
    wire N__33823;
    wire N__33820;
    wire N__33817;
    wire N__33814;
    wire N__33811;
    wire N__33808;
    wire N__33805;
    wire N__33802;
    wire N__33799;
    wire N__33796;
    wire N__33793;
    wire N__33790;
    wire N__33787;
    wire N__33784;
    wire N__33781;
    wire N__33778;
    wire N__33775;
    wire N__33772;
    wire N__33769;
    wire N__33766;
    wire N__33763;
    wire N__33760;
    wire N__33757;
    wire N__33754;
    wire N__33751;
    wire N__33748;
    wire N__33745;
    wire N__33742;
    wire N__33739;
    wire N__33736;
    wire N__33733;
    wire N__33730;
    wire N__33727;
    wire N__33724;
    wire N__33721;
    wire N__33718;
    wire N__33715;
    wire N__33712;
    wire N__33709;
    wire N__33706;
    wire N__33703;
    wire N__33700;
    wire N__33697;
    wire N__33694;
    wire N__33691;
    wire N__33688;
    wire N__33685;
    wire N__33682;
    wire N__33679;
    wire N__33676;
    wire N__33673;
    wire N__33670;
    wire N__33667;
    wire N__33664;
    wire N__33661;
    wire N__33658;
    wire N__33655;
    wire N__33652;
    wire N__33649;
    wire N__33646;
    wire N__33643;
    wire N__33640;
    wire N__33637;
    wire N__33634;
    wire N__33631;
    wire N__33628;
    wire N__33625;
    wire N__33622;
    wire N__33619;
    wire N__33616;
    wire N__33613;
    wire N__33610;
    wire N__33607;
    wire N__33604;
    wire N__33601;
    wire N__33598;
    wire N__33595;
    wire N__33592;
    wire N__33589;
    wire N__33586;
    wire N__33583;
    wire N__33580;
    wire N__33577;
    wire N__33574;
    wire N__33571;
    wire N__33568;
    wire N__33565;
    wire N__33562;
    wire N__33559;
    wire N__33556;
    wire N__33553;
    wire N__33550;
    wire N__33547;
    wire N__33544;
    wire N__33541;
    wire N__33538;
    wire N__33535;
    wire N__33532;
    wire N__33529;
    wire N__33526;
    wire N__33523;
    wire N__33520;
    wire N__33517;
    wire N__33514;
    wire N__33511;
    wire N__33508;
    wire N__33505;
    wire N__33502;
    wire N__33499;
    wire N__33496;
    wire N__33493;
    wire N__33490;
    wire N__33487;
    wire N__33484;
    wire N__33481;
    wire N__33478;
    wire N__33475;
    wire N__33472;
    wire N__33469;
    wire N__33466;
    wire N__33463;
    wire N__33460;
    wire N__33457;
    wire N__33454;
    wire N__33451;
    wire N__33450;
    wire N__33447;
    wire N__33444;
    wire N__33441;
    wire N__33438;
    wire N__33435;
    wire N__33432;
    wire N__33427;
    wire N__33424;
    wire N__33421;
    wire N__33420;
    wire N__33417;
    wire N__33414;
    wire N__33411;
    wire N__33408;
    wire N__33403;
    wire N__33400;
    wire N__33397;
    wire N__33394;
    wire N__33391;
    wire N__33388;
    wire N__33385;
    wire N__33382;
    wire N__33379;
    wire N__33376;
    wire N__33373;
    wire N__33370;
    wire N__33367;
    wire N__33364;
    wire N__33361;
    wire N__33358;
    wire N__33355;
    wire N__33352;
    wire N__33349;
    wire N__33346;
    wire N__33343;
    wire N__33340;
    wire N__33337;
    wire N__33334;
    wire N__33331;
    wire N__33328;
    wire N__33325;
    wire N__33322;
    wire N__33319;
    wire N__33318;
    wire N__33317;
    wire N__33316;
    wire N__33313;
    wire N__33310;
    wire N__33307;
    wire N__33304;
    wire N__33295;
    wire N__33292;
    wire N__33289;
    wire N__33286;
    wire N__33285;
    wire N__33280;
    wire N__33277;
    wire N__33274;
    wire N__33271;
    wire N__33268;
    wire N__33265;
    wire N__33262;
    wire N__33259;
    wire N__33258;
    wire N__33255;
    wire N__33252;
    wire N__33247;
    wire N__33244;
    wire N__33241;
    wire N__33238;
    wire N__33237;
    wire N__33234;
    wire N__33231;
    wire N__33228;
    wire N__33225;
    wire N__33220;
    wire N__33217;
    wire N__33214;
    wire N__33211;
    wire N__33208;
    wire N__33205;
    wire N__33202;
    wire N__33199;
    wire N__33198;
    wire N__33195;
    wire N__33192;
    wire N__33189;
    wire N__33184;
    wire N__33181;
    wire N__33178;
    wire N__33177;
    wire N__33176;
    wire N__33175;
    wire N__33172;
    wire N__33169;
    wire N__33166;
    wire N__33163;
    wire N__33154;
    wire N__33151;
    wire N__33148;
    wire N__33145;
    wire N__33142;
    wire N__33139;
    wire N__33136;
    wire N__33135;
    wire N__33134;
    wire N__33131;
    wire N__33128;
    wire N__33125;
    wire N__33122;
    wire N__33119;
    wire N__33116;
    wire N__33113;
    wire N__33110;
    wire N__33103;
    wire N__33100;
    wire N__33097;
    wire N__33094;
    wire N__33091;
    wire N__33088;
    wire N__33085;
    wire N__33082;
    wire N__33079;
    wire N__33076;
    wire N__33075;
    wire N__33072;
    wire N__33069;
    wire N__33068;
    wire N__33067;
    wire N__33062;
    wire N__33059;
    wire N__33056;
    wire N__33053;
    wire N__33050;
    wire N__33043;
    wire N__33042;
    wire N__33041;
    wire N__33038;
    wire N__33033;
    wire N__33028;
    wire N__33027;
    wire N__33026;
    wire N__33025;
    wire N__33022;
    wire N__33021;
    wire N__33018;
    wire N__33015;
    wire N__33010;
    wire N__33007;
    wire N__33004;
    wire N__32999;
    wire N__32996;
    wire N__32993;
    wire N__32990;
    wire N__32983;
    wire N__32982;
    wire N__32981;
    wire N__32978;
    wire N__32975;
    wire N__32974;
    wire N__32971;
    wire N__32966;
    wire N__32963;
    wire N__32960;
    wire N__32957;
    wire N__32954;
    wire N__32947;
    wire N__32946;
    wire N__32943;
    wire N__32940;
    wire N__32939;
    wire N__32938;
    wire N__32935;
    wire N__32932;
    wire N__32929;
    wire N__32926;
    wire N__32923;
    wire N__32918;
    wire N__32911;
    wire N__32910;
    wire N__32909;
    wire N__32904;
    wire N__32901;
    wire N__32898;
    wire N__32893;
    wire N__32892;
    wire N__32891;
    wire N__32890;
    wire N__32889;
    wire N__32886;
    wire N__32883;
    wire N__32880;
    wire N__32877;
    wire N__32874;
    wire N__32871;
    wire N__32868;
    wire N__32865;
    wire N__32862;
    wire N__32859;
    wire N__32856;
    wire N__32851;
    wire N__32848;
    wire N__32839;
    wire N__32836;
    wire N__32835;
    wire N__32834;
    wire N__32831;
    wire N__32828;
    wire N__32827;
    wire N__32824;
    wire N__32823;
    wire N__32818;
    wire N__32815;
    wire N__32812;
    wire N__32809;
    wire N__32802;
    wire N__32797;
    wire N__32796;
    wire N__32793;
    wire N__32790;
    wire N__32787;
    wire N__32784;
    wire N__32779;
    wire N__32778;
    wire N__32777;
    wire N__32774;
    wire N__32771;
    wire N__32768;
    wire N__32763;
    wire N__32758;
    wire N__32755;
    wire N__32752;
    wire N__32749;
    wire N__32746;
    wire N__32743;
    wire N__32742;
    wire N__32737;
    wire N__32734;
    wire N__32731;
    wire N__32730;
    wire N__32727;
    wire N__32724;
    wire N__32721;
    wire N__32718;
    wire N__32717;
    wire N__32714;
    wire N__32711;
    wire N__32708;
    wire N__32701;
    wire N__32698;
    wire N__32695;
    wire N__32692;
    wire N__32691;
    wire N__32690;
    wire N__32687;
    wire N__32684;
    wire N__32679;
    wire N__32674;
    wire N__32673;
    wire N__32672;
    wire N__32669;
    wire N__32666;
    wire N__32663;
    wire N__32660;
    wire N__32657;
    wire N__32656;
    wire N__32653;
    wire N__32650;
    wire N__32647;
    wire N__32644;
    wire N__32635;
    wire N__32632;
    wire N__32629;
    wire N__32626;
    wire N__32623;
    wire N__32620;
    wire N__32617;
    wire N__32614;
    wire N__32611;
    wire N__32608;
    wire N__32605;
    wire N__32602;
    wire N__32599;
    wire N__32596;
    wire N__32593;
    wire N__32590;
    wire N__32587;
    wire N__32584;
    wire N__32581;
    wire N__32578;
    wire N__32575;
    wire N__32572;
    wire N__32569;
    wire N__32566;
    wire N__32563;
    wire N__32560;
    wire N__32557;
    wire N__32554;
    wire N__32551;
    wire N__32548;
    wire N__32545;
    wire N__32542;
    wire N__32539;
    wire N__32536;
    wire N__32533;
    wire N__32530;
    wire N__32527;
    wire N__32524;
    wire N__32521;
    wire N__32518;
    wire N__32515;
    wire N__32512;
    wire N__32509;
    wire N__32506;
    wire N__32503;
    wire N__32500;
    wire N__32497;
    wire N__32494;
    wire N__32491;
    wire N__32488;
    wire N__32485;
    wire N__32482;
    wire N__32479;
    wire N__32476;
    wire N__32473;
    wire N__32470;
    wire N__32467;
    wire N__32464;
    wire N__32461;
    wire N__32458;
    wire N__32455;
    wire N__32452;
    wire N__32449;
    wire N__32446;
    wire N__32443;
    wire N__32440;
    wire N__32437;
    wire N__32434;
    wire N__32431;
    wire N__32428;
    wire N__32425;
    wire N__32422;
    wire N__32419;
    wire N__32416;
    wire N__32413;
    wire N__32410;
    wire N__32407;
    wire N__32404;
    wire N__32401;
    wire N__32398;
    wire N__32395;
    wire N__32392;
    wire N__32389;
    wire N__32386;
    wire N__32383;
    wire N__32380;
    wire N__32377;
    wire N__32374;
    wire N__32371;
    wire N__32368;
    wire N__32365;
    wire N__32362;
    wire N__32359;
    wire N__32356;
    wire N__32353;
    wire N__32350;
    wire N__32347;
    wire N__32344;
    wire N__32341;
    wire N__32338;
    wire N__32335;
    wire N__32332;
    wire N__32329;
    wire N__32326;
    wire N__32323;
    wire N__32320;
    wire N__32317;
    wire N__32314;
    wire N__32311;
    wire N__32308;
    wire N__32305;
    wire N__32302;
    wire N__32299;
    wire N__32296;
    wire N__32293;
    wire N__32290;
    wire N__32287;
    wire N__32284;
    wire N__32281;
    wire N__32278;
    wire N__32275;
    wire N__32272;
    wire N__32269;
    wire N__32266;
    wire N__32263;
    wire N__32260;
    wire N__32257;
    wire N__32254;
    wire N__32251;
    wire N__32248;
    wire N__32245;
    wire N__32242;
    wire N__32239;
    wire N__32236;
    wire N__32233;
    wire N__32230;
    wire N__32227;
    wire N__32224;
    wire N__32221;
    wire N__32218;
    wire N__32215;
    wire N__32212;
    wire N__32211;
    wire N__32208;
    wire N__32205;
    wire N__32202;
    wire N__32201;
    wire N__32198;
    wire N__32195;
    wire N__32192;
    wire N__32191;
    wire N__32188;
    wire N__32183;
    wire N__32180;
    wire N__32177;
    wire N__32174;
    wire N__32167;
    wire N__32166;
    wire N__32163;
    wire N__32160;
    wire N__32155;
    wire N__32154;
    wire N__32151;
    wire N__32148;
    wire N__32147;
    wire N__32144;
    wire N__32141;
    wire N__32138;
    wire N__32135;
    wire N__32132;
    wire N__32129;
    wire N__32126;
    wire N__32123;
    wire N__32122;
    wire N__32121;
    wire N__32120;
    wire N__32117;
    wire N__32112;
    wire N__32109;
    wire N__32104;
    wire N__32101;
    wire N__32096;
    wire N__32089;
    wire N__32086;
    wire N__32083;
    wire N__32082;
    wire N__32079;
    wire N__32076;
    wire N__32075;
    wire N__32072;
    wire N__32069;
    wire N__32066;
    wire N__32059;
    wire N__32056;
    wire N__32053;
    wire N__32050;
    wire N__32047;
    wire N__32044;
    wire N__32041;
    wire N__32038;
    wire N__32037;
    wire N__32036;
    wire N__32035;
    wire N__32034;
    wire N__32031;
    wire N__32028;
    wire N__32025;
    wire N__32020;
    wire N__32017;
    wire N__32014;
    wire N__32009;
    wire N__32002;
    wire N__32001;
    wire N__32000;
    wire N__31997;
    wire N__31996;
    wire N__31993;
    wire N__31992;
    wire N__31987;
    wire N__31984;
    wire N__31981;
    wire N__31978;
    wire N__31975;
    wire N__31972;
    wire N__31969;
    wire N__31964;
    wire N__31957;
    wire N__31954;
    wire N__31953;
    wire N__31952;
    wire N__31951;
    wire N__31948;
    wire N__31945;
    wire N__31942;
    wire N__31941;
    wire N__31938;
    wire N__31935;
    wire N__31932;
    wire N__31929;
    wire N__31926;
    wire N__31923;
    wire N__31920;
    wire N__31915;
    wire N__31912;
    wire N__31903;
    wire N__31902;
    wire N__31901;
    wire N__31898;
    wire N__31897;
    wire N__31894;
    wire N__31891;
    wire N__31888;
    wire N__31885;
    wire N__31880;
    wire N__31879;
    wire N__31876;
    wire N__31873;
    wire N__31870;
    wire N__31867;
    wire N__31864;
    wire N__31859;
    wire N__31852;
    wire N__31851;
    wire N__31850;
    wire N__31849;
    wire N__31848;
    wire N__31845;
    wire N__31842;
    wire N__31839;
    wire N__31836;
    wire N__31833;
    wire N__31830;
    wire N__31825;
    wire N__31822;
    wire N__31819;
    wire N__31812;
    wire N__31807;
    wire N__31806;
    wire N__31803;
    wire N__31800;
    wire N__31795;
    wire N__31794;
    wire N__31791;
    wire N__31788;
    wire N__31783;
    wire N__31782;
    wire N__31779;
    wire N__31776;
    wire N__31773;
    wire N__31768;
    wire N__31765;
    wire N__31762;
    wire N__31759;
    wire N__31756;
    wire N__31755;
    wire N__31754;
    wire N__31753;
    wire N__31752;
    wire N__31751;
    wire N__31750;
    wire N__31749;
    wire N__31748;
    wire N__31747;
    wire N__31746;
    wire N__31745;
    wire N__31744;
    wire N__31743;
    wire N__31742;
    wire N__31741;
    wire N__31740;
    wire N__31739;
    wire N__31738;
    wire N__31737;
    wire N__31736;
    wire N__31735;
    wire N__31734;
    wire N__31733;
    wire N__31732;
    wire N__31731;
    wire N__31720;
    wire N__31719;
    wire N__31718;
    wire N__31717;
    wire N__31716;
    wire N__31715;
    wire N__31704;
    wire N__31689;
    wire N__31678;
    wire N__31669;
    wire N__31668;
    wire N__31667;
    wire N__31666;
    wire N__31665;
    wire N__31664;
    wire N__31663;
    wire N__31662;
    wire N__31659;
    wire N__31648;
    wire N__31643;
    wire N__31638;
    wire N__31629;
    wire N__31622;
    wire N__31609;
    wire N__31606;
    wire N__31603;
    wire N__31600;
    wire N__31597;
    wire N__31594;
    wire N__31591;
    wire N__31588;
    wire N__31585;
    wire N__31584;
    wire N__31583;
    wire N__31582;
    wire N__31579;
    wire N__31576;
    wire N__31573;
    wire N__31570;
    wire N__31561;
    wire N__31560;
    wire N__31559;
    wire N__31558;
    wire N__31555;
    wire N__31552;
    wire N__31551;
    wire N__31546;
    wire N__31543;
    wire N__31540;
    wire N__31537;
    wire N__31534;
    wire N__31525;
    wire N__31524;
    wire N__31523;
    wire N__31522;
    wire N__31521;
    wire N__31520;
    wire N__31517;
    wire N__31514;
    wire N__31513;
    wire N__31512;
    wire N__31511;
    wire N__31510;
    wire N__31509;
    wire N__31508;
    wire N__31507;
    wire N__31506;
    wire N__31503;
    wire N__31502;
    wire N__31501;
    wire N__31500;
    wire N__31499;
    wire N__31498;
    wire N__31497;
    wire N__31494;
    wire N__31493;
    wire N__31492;
    wire N__31489;
    wire N__31486;
    wire N__31485;
    wire N__31484;
    wire N__31483;
    wire N__31482;
    wire N__31481;
    wire N__31480;
    wire N__31479;
    wire N__31478;
    wire N__31467;
    wire N__31456;
    wire N__31441;
    wire N__31440;
    wire N__31437;
    wire N__31428;
    wire N__31421;
    wire N__31410;
    wire N__31405;
    wire N__31402;
    wire N__31401;
    wire N__31400;
    wire N__31397;
    wire N__31396;
    wire N__31395;
    wire N__31394;
    wire N__31393;
    wire N__31392;
    wire N__31391;
    wire N__31390;
    wire N__31389;
    wire N__31384;
    wire N__31379;
    wire N__31374;
    wire N__31371;
    wire N__31358;
    wire N__31349;
    wire N__31346;
    wire N__31343;
    wire N__31340;
    wire N__31327;
    wire N__31326;
    wire N__31325;
    wire N__31322;
    wire N__31319;
    wire N__31318;
    wire N__31317;
    wire N__31314;
    wire N__31311;
    wire N__31308;
    wire N__31305;
    wire N__31302;
    wire N__31299;
    wire N__31294;
    wire N__31291;
    wire N__31282;
    wire N__31281;
    wire N__31280;
    wire N__31279;
    wire N__31278;
    wire N__31275;
    wire N__31272;
    wire N__31269;
    wire N__31264;
    wire N__31261;
    wire N__31258;
    wire N__31253;
    wire N__31246;
    wire N__31245;
    wire N__31244;
    wire N__31241;
    wire N__31240;
    wire N__31239;
    wire N__31236;
    wire N__31233;
    wire N__31230;
    wire N__31225;
    wire N__31222;
    wire N__31219;
    wire N__31216;
    wire N__31213;
    wire N__31204;
    wire N__31203;
    wire N__31202;
    wire N__31201;
    wire N__31198;
    wire N__31197;
    wire N__31192;
    wire N__31189;
    wire N__31186;
    wire N__31183;
    wire N__31180;
    wire N__31177;
    wire N__31170;
    wire N__31165;
    wire N__31164;
    wire N__31163;
    wire N__31160;
    wire N__31157;
    wire N__31156;
    wire N__31153;
    wire N__31152;
    wire N__31147;
    wire N__31144;
    wire N__31141;
    wire N__31138;
    wire N__31135;
    wire N__31130;
    wire N__31123;
    wire N__31120;
    wire N__31117;
    wire N__31114;
    wire N__31111;
    wire N__31108;
    wire N__31107;
    wire N__31106;
    wire N__31105;
    wire N__31104;
    wire N__31103;
    wire N__31102;
    wire N__31101;
    wire N__31100;
    wire N__31099;
    wire N__31098;
    wire N__31097;
    wire N__31096;
    wire N__31095;
    wire N__31094;
    wire N__31093;
    wire N__31090;
    wire N__31087;
    wire N__31084;
    wire N__31081;
    wire N__31080;
    wire N__31079;
    wire N__31078;
    wire N__31077;
    wire N__31074;
    wire N__31071;
    wire N__31068;
    wire N__31065;
    wire N__31062;
    wire N__31059;
    wire N__31056;
    wire N__31053;
    wire N__31050;
    wire N__31047;
    wire N__31044;
    wire N__31027;
    wire N__31026;
    wire N__31023;
    wire N__31022;
    wire N__31013;
    wire N__31004;
    wire N__30999;
    wire N__30996;
    wire N__30993;
    wire N__30990;
    wire N__30989;
    wire N__30984;
    wire N__30979;
    wire N__30976;
    wire N__30973;
    wire N__30972;
    wire N__30967;
    wire N__30964;
    wire N__30959;
    wire N__30954;
    wire N__30951;
    wire N__30948;
    wire N__30945;
    wire N__30942;
    wire N__30937;
    wire N__30934;
    wire N__30925;
    wire N__30924;
    wire N__30923;
    wire N__30922;
    wire N__30919;
    wire N__30916;
    wire N__30913;
    wire N__30910;
    wire N__30909;
    wire N__30908;
    wire N__30907;
    wire N__30906;
    wire N__30905;
    wire N__30904;
    wire N__30903;
    wire N__30902;
    wire N__30901;
    wire N__30900;
    wire N__30899;
    wire N__30898;
    wire N__30897;
    wire N__30896;
    wire N__30895;
    wire N__30894;
    wire N__30893;
    wire N__30892;
    wire N__30883;
    wire N__30880;
    wire N__30863;
    wire N__30854;
    wire N__30851;
    wire N__30848;
    wire N__30845;
    wire N__30844;
    wire N__30843;
    wire N__30838;
    wire N__30829;
    wire N__30826;
    wire N__30821;
    wire N__30816;
    wire N__30811;
    wire N__30806;
    wire N__30799;
    wire N__30798;
    wire N__30797;
    wire N__30796;
    wire N__30795;
    wire N__30794;
    wire N__30793;
    wire N__30792;
    wire N__30791;
    wire N__30788;
    wire N__30771;
    wire N__30770;
    wire N__30769;
    wire N__30768;
    wire N__30767;
    wire N__30766;
    wire N__30765;
    wire N__30764;
    wire N__30763;
    wire N__30762;
    wire N__30761;
    wire N__30760;
    wire N__30759;
    wire N__30758;
    wire N__30757;
    wire N__30752;
    wire N__30749;
    wire N__30746;
    wire N__30741;
    wire N__30724;
    wire N__30721;
    wire N__30718;
    wire N__30717;
    wire N__30712;
    wire N__30709;
    wire N__30702;
    wire N__30697;
    wire N__30692;
    wire N__30689;
    wire N__30682;
    wire N__30681;
    wire N__30678;
    wire N__30675;
    wire N__30670;
    wire N__30667;
    wire N__30664;
    wire N__30661;
    wire N__30658;
    wire N__30655;
    wire N__30652;
    wire N__30649;
    wire N__30646;
    wire N__30643;
    wire N__30640;
    wire N__30637;
    wire N__30634;
    wire N__30631;
    wire N__30628;
    wire N__30625;
    wire N__30622;
    wire N__30619;
    wire N__30616;
    wire N__30613;
    wire N__30612;
    wire N__30611;
    wire N__30608;
    wire N__30605;
    wire N__30602;
    wire N__30599;
    wire N__30596;
    wire N__30595;
    wire N__30592;
    wire N__30589;
    wire N__30586;
    wire N__30583;
    wire N__30580;
    wire N__30577;
    wire N__30574;
    wire N__30571;
    wire N__30562;
    wire N__30559;
    wire N__30556;
    wire N__30553;
    wire N__30552;
    wire N__30551;
    wire N__30550;
    wire N__30549;
    wire N__30546;
    wire N__30545;
    wire N__30544;
    wire N__30543;
    wire N__30540;
    wire N__30533;
    wire N__30530;
    wire N__30523;
    wire N__30520;
    wire N__30517;
    wire N__30508;
    wire N__30505;
    wire N__30502;
    wire N__30499;
    wire N__30498;
    wire N__30497;
    wire N__30496;
    wire N__30493;
    wire N__30490;
    wire N__30487;
    wire N__30484;
    wire N__30481;
    wire N__30478;
    wire N__30469;
    wire N__30466;
    wire N__30463;
    wire N__30460;
    wire N__30457;
    wire N__30454;
    wire N__30451;
    wire N__30448;
    wire N__30447;
    wire N__30446;
    wire N__30445;
    wire N__30444;
    wire N__30443;
    wire N__30442;
    wire N__30441;
    wire N__30440;
    wire N__30439;
    wire N__30438;
    wire N__30437;
    wire N__30436;
    wire N__30435;
    wire N__30430;
    wire N__30429;
    wire N__30428;
    wire N__30427;
    wire N__30426;
    wire N__30425;
    wire N__30424;
    wire N__30423;
    wire N__30422;
    wire N__30405;
    wire N__30402;
    wire N__30397;
    wire N__30394;
    wire N__30391;
    wire N__30390;
    wire N__30389;
    wire N__30372;
    wire N__30369;
    wire N__30366;
    wire N__30361;
    wire N__30358;
    wire N__30353;
    wire N__30346;
    wire N__30343;
    wire N__30340;
    wire N__30331;
    wire N__30328;
    wire N__30327;
    wire N__30326;
    wire N__30325;
    wire N__30324;
    wire N__30323;
    wire N__30322;
    wire N__30321;
    wire N__30320;
    wire N__30319;
    wire N__30318;
    wire N__30317;
    wire N__30316;
    wire N__30315;
    wire N__30310;
    wire N__30309;
    wire N__30308;
    wire N__30307;
    wire N__30304;
    wire N__30301;
    wire N__30298;
    wire N__30295;
    wire N__30294;
    wire N__30293;
    wire N__30292;
    wire N__30291;
    wire N__30274;
    wire N__30271;
    wire N__30268;
    wire N__30265;
    wire N__30262;
    wire N__30261;
    wire N__30260;
    wire N__30243;
    wire N__30240;
    wire N__30239;
    wire N__30234;
    wire N__30229;
    wire N__30224;
    wire N__30221;
    wire N__30218;
    wire N__30215;
    wire N__30212;
    wire N__30199;
    wire N__30198;
    wire N__30197;
    wire N__30196;
    wire N__30195;
    wire N__30194;
    wire N__30193;
    wire N__30192;
    wire N__30191;
    wire N__30190;
    wire N__30189;
    wire N__30188;
    wire N__30187;
    wire N__30186;
    wire N__30185;
    wire N__30184;
    wire N__30183;
    wire N__30182;
    wire N__30181;
    wire N__30180;
    wire N__30179;
    wire N__30176;
    wire N__30173;
    wire N__30170;
    wire N__30167;
    wire N__30166;
    wire N__30149;
    wire N__30148;
    wire N__30143;
    wire N__30140;
    wire N__30139;
    wire N__30134;
    wire N__30117;
    wire N__30114;
    wire N__30111;
    wire N__30108;
    wire N__30105;
    wire N__30100;
    wire N__30097;
    wire N__30092;
    wire N__30085;
    wire N__30076;
    wire N__30075;
    wire N__30072;
    wire N__30069;
    wire N__30066;
    wire N__30065;
    wire N__30062;
    wire N__30061;
    wire N__30058;
    wire N__30055;
    wire N__30052;
    wire N__30049;
    wire N__30040;
    wire N__30037;
    wire N__30034;
    wire N__30033;
    wire N__30032;
    wire N__30031;
    wire N__30028;
    wire N__30021;
    wire N__30020;
    wire N__30019;
    wire N__30016;
    wire N__30013;
    wire N__30008;
    wire N__30001;
    wire N__29998;
    wire N__29995;
    wire N__29994;
    wire N__29993;
    wire N__29992;
    wire N__29991;
    wire N__29990;
    wire N__29989;
    wire N__29984;
    wire N__29983;
    wire N__29982;
    wire N__29981;
    wire N__29978;
    wire N__29975;
    wire N__29972;
    wire N__29969;
    wire N__29966;
    wire N__29965;
    wire N__29964;
    wire N__29963;
    wire N__29960;
    wire N__29959;
    wire N__29958;
    wire N__29957;
    wire N__29956;
    wire N__29955;
    wire N__29942;
    wire N__29931;
    wire N__29928;
    wire N__29927;
    wire N__29926;
    wire N__29923;
    wire N__29920;
    wire N__29917;
    wire N__29914;
    wire N__29911;
    wire N__29910;
    wire N__29909;
    wire N__29908;
    wire N__29907;
    wire N__29900;
    wire N__29895;
    wire N__29892;
    wire N__29877;
    wire N__29874;
    wire N__29869;
    wire N__29860;
    wire N__29859;
    wire N__29858;
    wire N__29855;
    wire N__29852;
    wire N__29849;
    wire N__29848;
    wire N__29845;
    wire N__29840;
    wire N__29837;
    wire N__29836;
    wire N__29835;
    wire N__29830;
    wire N__29827;
    wire N__29822;
    wire N__29815;
    wire N__29814;
    wire N__29813;
    wire N__29812;
    wire N__29811;
    wire N__29810;
    wire N__29809;
    wire N__29808;
    wire N__29807;
    wire N__29806;
    wire N__29805;
    wire N__29804;
    wire N__29803;
    wire N__29802;
    wire N__29801;
    wire N__29800;
    wire N__29799;
    wire N__29798;
    wire N__29797;
    wire N__29794;
    wire N__29779;
    wire N__29766;
    wire N__29755;
    wire N__29754;
    wire N__29753;
    wire N__29752;
    wire N__29747;
    wire N__29742;
    wire N__29735;
    wire N__29734;
    wire N__29733;
    wire N__29726;
    wire N__29723;
    wire N__29720;
    wire N__29717;
    wire N__29714;
    wire N__29711;
    wire N__29708;
    wire N__29701;
    wire N__29700;
    wire N__29699;
    wire N__29698;
    wire N__29697;
    wire N__29696;
    wire N__29695;
    wire N__29694;
    wire N__29693;
    wire N__29692;
    wire N__29691;
    wire N__29690;
    wire N__29689;
    wire N__29686;
    wire N__29671;
    wire N__29660;
    wire N__29659;
    wire N__29658;
    wire N__29657;
    wire N__29656;
    wire N__29655;
    wire N__29654;
    wire N__29653;
    wire N__29652;
    wire N__29651;
    wire N__29646;
    wire N__29643;
    wire N__29640;
    wire N__29635;
    wire N__29622;
    wire N__29613;
    wire N__29612;
    wire N__29611;
    wire N__29608;
    wire N__29605;
    wire N__29600;
    wire N__29597;
    wire N__29594;
    wire N__29587;
    wire N__29584;
    wire N__29581;
    wire N__29578;
    wire N__29575;
    wire N__29572;
    wire N__29569;
    wire N__29566;
    wire N__29563;
    wire N__29560;
    wire N__29557;
    wire N__29554;
    wire N__29551;
    wire N__29548;
    wire N__29545;
    wire N__29542;
    wire N__29539;
    wire N__29536;
    wire N__29533;
    wire N__29530;
    wire N__29527;
    wire N__29524;
    wire N__29521;
    wire N__29518;
    wire N__29515;
    wire N__29512;
    wire N__29509;
    wire N__29506;
    wire N__29503;
    wire N__29500;
    wire N__29497;
    wire N__29496;
    wire N__29491;
    wire N__29490;
    wire N__29489;
    wire N__29488;
    wire N__29487;
    wire N__29484;
    wire N__29475;
    wire N__29470;
    wire N__29467;
    wire N__29464;
    wire N__29461;
    wire N__29458;
    wire N__29457;
    wire N__29456;
    wire N__29453;
    wire N__29450;
    wire N__29447;
    wire N__29444;
    wire N__29443;
    wire N__29440;
    wire N__29437;
    wire N__29434;
    wire N__29431;
    wire N__29426;
    wire N__29419;
    wire N__29418;
    wire N__29417;
    wire N__29414;
    wire N__29411;
    wire N__29408;
    wire N__29407;
    wire N__29404;
    wire N__29399;
    wire N__29396;
    wire N__29391;
    wire N__29386;
    wire N__29385;
    wire N__29384;
    wire N__29383;
    wire N__29376;
    wire N__29375;
    wire N__29374;
    wire N__29373;
    wire N__29370;
    wire N__29367;
    wire N__29362;
    wire N__29359;
    wire N__29358;
    wire N__29357;
    wire N__29354;
    wire N__29347;
    wire N__29342;
    wire N__29335;
    wire N__29334;
    wire N__29333;
    wire N__29330;
    wire N__29329;
    wire N__29326;
    wire N__29323;
    wire N__29320;
    wire N__29317;
    wire N__29314;
    wire N__29309;
    wire N__29306;
    wire N__29301;
    wire N__29296;
    wire N__29293;
    wire N__29290;
    wire N__29289;
    wire N__29288;
    wire N__29287;
    wire N__29284;
    wire N__29281;
    wire N__29278;
    wire N__29275;
    wire N__29266;
    wire N__29263;
    wire N__29260;
    wire N__29257;
    wire N__29254;
    wire N__29251;
    wire N__29248;
    wire N__29247;
    wire N__29244;
    wire N__29241;
    wire N__29236;
    wire N__29233;
    wire N__29230;
    wire N__29227;
    wire N__29224;
    wire N__29223;
    wire N__29218;
    wire N__29215;
    wire N__29214;
    wire N__29213;
    wire N__29212;
    wire N__29211;
    wire N__29210;
    wire N__29209;
    wire N__29204;
    wire N__29195;
    wire N__29192;
    wire N__29185;
    wire N__29182;
    wire N__29179;
    wire N__29176;
    wire N__29173;
    wire N__29170;
    wire N__29167;
    wire N__29166;
    wire N__29163;
    wire N__29162;
    wire N__29159;
    wire N__29156;
    wire N__29153;
    wire N__29146;
    wire N__29143;
    wire N__29140;
    wire N__29137;
    wire N__29134;
    wire N__29131;
    wire N__29128;
    wire N__29125;
    wire N__29122;
    wire N__29119;
    wire N__29116;
    wire N__29113;
    wire N__29110;
    wire N__29107;
    wire N__29104;
    wire N__29101;
    wire N__29098;
    wire N__29097;
    wire N__29092;
    wire N__29089;
    wire N__29086;
    wire N__29083;
    wire N__29080;
    wire N__29077;
    wire N__29074;
    wire N__29071;
    wire N__29068;
    wire N__29065;
    wire N__29062;
    wire N__29059;
    wire N__29056;
    wire N__29055;
    wire N__29054;
    wire N__29053;
    wire N__29052;
    wire N__29051;
    wire N__29048;
    wire N__29045;
    wire N__29042;
    wire N__29039;
    wire N__29030;
    wire N__29029;
    wire N__29028;
    wire N__29023;
    wire N__29020;
    wire N__29017;
    wire N__29014;
    wire N__29005;
    wire N__29002;
    wire N__28999;
    wire N__28996;
    wire N__28993;
    wire N__28990;
    wire N__28987;
    wire N__28984;
    wire N__28981;
    wire N__28978;
    wire N__28975;
    wire N__28972;
    wire N__28969;
    wire N__28966;
    wire N__28963;
    wire N__28960;
    wire N__28957;
    wire N__28954;
    wire N__28951;
    wire N__28948;
    wire N__28945;
    wire N__28942;
    wire N__28939;
    wire N__28936;
    wire N__28933;
    wire N__28930;
    wire N__28927;
    wire N__28924;
    wire N__28921;
    wire N__28918;
    wire N__28915;
    wire N__28912;
    wire N__28909;
    wire N__28906;
    wire N__28903;
    wire N__28900;
    wire N__28897;
    wire N__28894;
    wire N__28891;
    wire N__28888;
    wire N__28885;
    wire N__28882;
    wire N__28879;
    wire N__28876;
    wire N__28873;
    wire N__28870;
    wire N__28867;
    wire N__28864;
    wire N__28861;
    wire N__28858;
    wire N__28855;
    wire N__28852;
    wire N__28849;
    wire N__28846;
    wire N__28843;
    wire N__28840;
    wire N__28837;
    wire N__28834;
    wire N__28831;
    wire N__28830;
    wire N__28829;
    wire N__28828;
    wire N__28825;
    wire N__28818;
    wire N__28815;
    wire N__28812;
    wire N__28807;
    wire N__28806;
    wire N__28803;
    wire N__28800;
    wire N__28795;
    wire N__28792;
    wire N__28789;
    wire N__28786;
    wire N__28783;
    wire N__28780;
    wire N__28777;
    wire N__28774;
    wire N__28771;
    wire N__28768;
    wire N__28765;
    wire N__28762;
    wire N__28759;
    wire N__28756;
    wire N__28753;
    wire N__28750;
    wire N__28747;
    wire N__28744;
    wire N__28741;
    wire N__28738;
    wire N__28735;
    wire N__28732;
    wire N__28729;
    wire N__28726;
    wire N__28723;
    wire N__28720;
    wire N__28717;
    wire N__28714;
    wire N__28711;
    wire N__28708;
    wire N__28705;
    wire N__28702;
    wire N__28699;
    wire N__28696;
    wire N__28693;
    wire N__28690;
    wire N__28687;
    wire N__28684;
    wire N__28681;
    wire N__28678;
    wire N__28675;
    wire N__28672;
    wire N__28669;
    wire N__28666;
    wire N__28663;
    wire N__28662;
    wire N__28659;
    wire N__28656;
    wire N__28651;
    wire N__28648;
    wire N__28645;
    wire N__28642;
    wire N__28639;
    wire N__28636;
    wire N__28633;
    wire N__28632;
    wire N__28629;
    wire N__28626;
    wire N__28623;
    wire N__28618;
    wire N__28615;
    wire N__28612;
    wire N__28609;
    wire N__28608;
    wire N__28605;
    wire N__28602;
    wire N__28599;
    wire N__28594;
    wire N__28591;
    wire N__28588;
    wire N__28585;
    wire N__28582;
    wire N__28581;
    wire N__28578;
    wire N__28575;
    wire N__28572;
    wire N__28567;
    wire N__28564;
    wire N__28561;
    wire N__28558;
    wire N__28557;
    wire N__28554;
    wire N__28551;
    wire N__28548;
    wire N__28543;
    wire N__28540;
    wire N__28537;
    wire N__28534;
    wire N__28531;
    wire N__28530;
    wire N__28527;
    wire N__28524;
    wire N__28519;
    wire N__28516;
    wire N__28513;
    wire N__28510;
    wire N__28509;
    wire N__28506;
    wire N__28503;
    wire N__28498;
    wire N__28495;
    wire N__28492;
    wire N__28489;
    wire N__28486;
    wire N__28485;
    wire N__28482;
    wire N__28479;
    wire N__28474;
    wire N__28471;
    wire N__28468;
    wire N__28465;
    wire N__28462;
    wire N__28461;
    wire N__28458;
    wire N__28455;
    wire N__28450;
    wire N__28447;
    wire N__28444;
    wire N__28441;
    wire N__28440;
    wire N__28437;
    wire N__28434;
    wire N__28429;
    wire N__28426;
    wire N__28423;
    wire N__28420;
    wire N__28417;
    wire N__28416;
    wire N__28413;
    wire N__28410;
    wire N__28405;
    wire N__28402;
    wire N__28399;
    wire N__28396;
    wire N__28395;
    wire N__28392;
    wire N__28389;
    wire N__28384;
    wire N__28381;
    wire N__28378;
    wire N__28375;
    wire N__28372;
    wire N__28371;
    wire N__28368;
    wire N__28365;
    wire N__28360;
    wire N__28357;
    wire N__28354;
    wire N__28351;
    wire N__28350;
    wire N__28347;
    wire N__28344;
    wire N__28339;
    wire N__28336;
    wire N__28333;
    wire N__28330;
    wire N__28327;
    wire N__28324;
    wire N__28323;
    wire N__28320;
    wire N__28317;
    wire N__28312;
    wire N__28309;
    wire N__28306;
    wire N__28303;
    wire N__28300;
    wire N__28297;
    wire N__28296;
    wire N__28293;
    wire N__28290;
    wire N__28285;
    wire N__28282;
    wire N__28279;
    wire N__28276;
    wire N__28273;
    wire N__28270;
    wire N__28267;
    wire N__28264;
    wire N__28261;
    wire N__28260;
    wire N__28259;
    wire N__28256;
    wire N__28253;
    wire N__28250;
    wire N__28247;
    wire N__28244;
    wire N__28237;
    wire N__28236;
    wire N__28233;
    wire N__28230;
    wire N__28225;
    wire N__28222;
    wire N__28219;
    wire N__28216;
    wire N__28213;
    wire N__28210;
    wire N__28207;
    wire N__28204;
    wire N__28203;
    wire N__28202;
    wire N__28199;
    wire N__28196;
    wire N__28193;
    wire N__28186;
    wire N__28183;
    wire N__28180;
    wire N__28179;
    wire N__28178;
    wire N__28175;
    wire N__28172;
    wire N__28169;
    wire N__28162;
    wire N__28159;
    wire N__28158;
    wire N__28155;
    wire N__28154;
    wire N__28151;
    wire N__28148;
    wire N__28145;
    wire N__28142;
    wire N__28135;
    wire N__28132;
    wire N__28131;
    wire N__28128;
    wire N__28127;
    wire N__28124;
    wire N__28121;
    wire N__28118;
    wire N__28115;
    wire N__28108;
    wire N__28105;
    wire N__28102;
    wire N__28101;
    wire N__28100;
    wire N__28099;
    wire N__28096;
    wire N__28093;
    wire N__28088;
    wire N__28081;
    wire N__28080;
    wire N__28077;
    wire N__28074;
    wire N__28071;
    wire N__28068;
    wire N__28067;
    wire N__28066;
    wire N__28061;
    wire N__28058;
    wire N__28055;
    wire N__28052;
    wire N__28045;
    wire N__28042;
    wire N__28039;
    wire N__28036;
    wire N__28033;
    wire N__28030;
    wire N__28029;
    wire N__28026;
    wire N__28023;
    wire N__28020;
    wire N__28019;
    wire N__28016;
    wire N__28013;
    wire N__28010;
    wire N__28007;
    wire N__28000;
    wire N__27999;
    wire N__27996;
    wire N__27993;
    wire N__27990;
    wire N__27989;
    wire N__27988;
    wire N__27985;
    wire N__27982;
    wire N__27979;
    wire N__27976;
    wire N__27971;
    wire N__27968;
    wire N__27961;
    wire N__27958;
    wire N__27955;
    wire N__27952;
    wire N__27949;
    wire N__27948;
    wire N__27945;
    wire N__27942;
    wire N__27941;
    wire N__27938;
    wire N__27935;
    wire N__27932;
    wire N__27929;
    wire N__27926;
    wire N__27919;
    wire N__27916;
    wire N__27915;
    wire N__27912;
    wire N__27909;
    wire N__27908;
    wire N__27905;
    wire N__27902;
    wire N__27899;
    wire N__27896;
    wire N__27893;
    wire N__27886;
    wire N__27883;
    wire N__27882;
    wire N__27881;
    wire N__27878;
    wire N__27875;
    wire N__27872;
    wire N__27867;
    wire N__27864;
    wire N__27861;
    wire N__27856;
    wire N__27853;
    wire N__27850;
    wire N__27849;
    wire N__27848;
    wire N__27845;
    wire N__27842;
    wire N__27839;
    wire N__27834;
    wire N__27829;
    wire N__27828;
    wire N__27825;
    wire N__27822;
    wire N__27821;
    wire N__27818;
    wire N__27815;
    wire N__27812;
    wire N__27809;
    wire N__27804;
    wire N__27799;
    wire N__27796;
    wire N__27793;
    wire N__27792;
    wire N__27789;
    wire N__27786;
    wire N__27783;
    wire N__27780;
    wire N__27775;
    wire N__27772;
    wire N__27771;
    wire N__27770;
    wire N__27767;
    wire N__27766;
    wire N__27765;
    wire N__27760;
    wire N__27757;
    wire N__27752;
    wire N__27749;
    wire N__27742;
    wire N__27739;
    wire N__27736;
    wire N__27733;
    wire N__27730;
    wire N__27727;
    wire N__27724;
    wire N__27721;
    wire N__27718;
    wire N__27715;
    wire N__27712;
    wire N__27711;
    wire N__27710;
    wire N__27707;
    wire N__27706;
    wire N__27703;
    wire N__27700;
    wire N__27697;
    wire N__27694;
    wire N__27691;
    wire N__27688;
    wire N__27685;
    wire N__27680;
    wire N__27673;
    wire N__27670;
    wire N__27667;
    wire N__27664;
    wire N__27661;
    wire N__27658;
    wire N__27655;
    wire N__27652;
    wire N__27649;
    wire N__27646;
    wire N__27643;
    wire N__27642;
    wire N__27639;
    wire N__27636;
    wire N__27635;
    wire N__27630;
    wire N__27627;
    wire N__27624;
    wire N__27619;
    wire N__27616;
    wire N__27613;
    wire N__27610;
    wire N__27607;
    wire N__27604;
    wire N__27601;
    wire N__27598;
    wire N__27595;
    wire N__27592;
    wire N__27589;
    wire N__27586;
    wire N__27583;
    wire N__27580;
    wire N__27577;
    wire N__27574;
    wire N__27571;
    wire N__27568;
    wire N__27567;
    wire N__27566;
    wire N__27563;
    wire N__27562;
    wire N__27559;
    wire N__27556;
    wire N__27553;
    wire N__27550;
    wire N__27547;
    wire N__27542;
    wire N__27539;
    wire N__27534;
    wire N__27531;
    wire N__27526;
    wire N__27523;
    wire N__27520;
    wire N__27517;
    wire N__27514;
    wire N__27511;
    wire N__27508;
    wire N__27505;
    wire N__27502;
    wire N__27501;
    wire N__27498;
    wire N__27495;
    wire N__27490;
    wire N__27487;
    wire N__27484;
    wire N__27481;
    wire N__27480;
    wire N__27477;
    wire N__27474;
    wire N__27469;
    wire N__27466;
    wire N__27463;
    wire N__27460;
    wire N__27459;
    wire N__27456;
    wire N__27453;
    wire N__27448;
    wire N__27445;
    wire N__27442;
    wire N__27439;
    wire N__27438;
    wire N__27435;
    wire N__27432;
    wire N__27429;
    wire N__27424;
    wire N__27421;
    wire N__27418;
    wire N__27415;
    wire N__27412;
    wire N__27409;
    wire N__27406;
    wire N__27403;
    wire N__27400;
    wire N__27397;
    wire N__27394;
    wire N__27393;
    wire N__27392;
    wire N__27389;
    wire N__27386;
    wire N__27385;
    wire N__27382;
    wire N__27379;
    wire N__27376;
    wire N__27373;
    wire N__27364;
    wire N__27363;
    wire N__27360;
    wire N__27359;
    wire N__27356;
    wire N__27353;
    wire N__27350;
    wire N__27343;
    wire N__27342;
    wire N__27339;
    wire N__27336;
    wire N__27331;
    wire N__27328;
    wire N__27325;
    wire N__27322;
    wire N__27319;
    wire N__27318;
    wire N__27315;
    wire N__27312;
    wire N__27307;
    wire N__27304;
    wire N__27301;
    wire N__27298;
    wire N__27295;
    wire N__27292;
    wire N__27291;
    wire N__27288;
    wire N__27285;
    wire N__27280;
    wire N__27277;
    wire N__27274;
    wire N__27271;
    wire N__27268;
    wire N__27267;
    wire N__27264;
    wire N__27261;
    wire N__27258;
    wire N__27253;
    wire N__27250;
    wire N__27247;
    wire N__27244;
    wire N__27243;
    wire N__27240;
    wire N__27237;
    wire N__27234;
    wire N__27229;
    wire N__27226;
    wire N__27223;
    wire N__27220;
    wire N__27219;
    wire N__27216;
    wire N__27213;
    wire N__27210;
    wire N__27205;
    wire N__27202;
    wire N__27199;
    wire N__27196;
    wire N__27195;
    wire N__27192;
    wire N__27189;
    wire N__27186;
    wire N__27181;
    wire N__27178;
    wire N__27175;
    wire N__27172;
    wire N__27171;
    wire N__27168;
    wire N__27165;
    wire N__27162;
    wire N__27157;
    wire N__27154;
    wire N__27151;
    wire N__27148;
    wire N__27145;
    wire N__27142;
    wire N__27141;
    wire N__27138;
    wire N__27135;
    wire N__27132;
    wire N__27129;
    wire N__27128;
    wire N__27123;
    wire N__27120;
    wire N__27115;
    wire N__27114;
    wire N__27111;
    wire N__27108;
    wire N__27103;
    wire N__27100;
    wire N__27097;
    wire N__27094;
    wire N__27091;
    wire N__27088;
    wire N__27085;
    wire N__27084;
    wire N__27081;
    wire N__27078;
    wire N__27073;
    wire N__27070;
    wire N__27067;
    wire N__27064;
    wire N__27063;
    wire N__27060;
    wire N__27057;
    wire N__27052;
    wire N__27049;
    wire N__27046;
    wire N__27043;
    wire N__27042;
    wire N__27039;
    wire N__27036;
    wire N__27031;
    wire N__27028;
    wire N__27025;
    wire N__27022;
    wire N__27021;
    wire N__27018;
    wire N__27015;
    wire N__27010;
    wire N__27007;
    wire N__27004;
    wire N__27001;
    wire N__27000;
    wire N__26997;
    wire N__26994;
    wire N__26989;
    wire N__26986;
    wire N__26983;
    wire N__26980;
    wire N__26977;
    wire N__26974;
    wire N__26971;
    wire N__26968;
    wire N__26965;
    wire N__26962;
    wire N__26959;
    wire N__26956;
    wire N__26953;
    wire N__26950;
    wire N__26947;
    wire N__26944;
    wire N__26941;
    wire N__26938;
    wire N__26935;
    wire N__26932;
    wire N__26929;
    wire N__26926;
    wire N__26923;
    wire N__26920;
    wire N__26917;
    wire N__26914;
    wire N__26911;
    wire N__26908;
    wire N__26905;
    wire N__26902;
    wire N__26899;
    wire N__26896;
    wire N__26893;
    wire N__26890;
    wire N__26887;
    wire N__26884;
    wire N__26881;
    wire N__26878;
    wire N__26875;
    wire N__26872;
    wire N__26869;
    wire N__26866;
    wire N__26863;
    wire N__26860;
    wire N__26857;
    wire N__26854;
    wire N__26851;
    wire N__26848;
    wire N__26845;
    wire N__26842;
    wire N__26839;
    wire N__26836;
    wire N__26833;
    wire N__26830;
    wire N__26827;
    wire N__26824;
    wire N__26821;
    wire N__26818;
    wire N__26815;
    wire N__26812;
    wire N__26809;
    wire N__26806;
    wire N__26803;
    wire N__26800;
    wire N__26797;
    wire N__26794;
    wire N__26791;
    wire N__26788;
    wire N__26785;
    wire N__26782;
    wire N__26779;
    wire N__26776;
    wire N__26773;
    wire N__26770;
    wire N__26767;
    wire N__26764;
    wire N__26761;
    wire N__26760;
    wire N__26759;
    wire N__26756;
    wire N__26755;
    wire N__26754;
    wire N__26751;
    wire N__26750;
    wire N__26749;
    wire N__26746;
    wire N__26733;
    wire N__26732;
    wire N__26731;
    wire N__26730;
    wire N__26729;
    wire N__26728;
    wire N__26725;
    wire N__26722;
    wire N__26719;
    wire N__26718;
    wire N__26717;
    wire N__26716;
    wire N__26715;
    wire N__26706;
    wire N__26699;
    wire N__26690;
    wire N__26683;
    wire N__26680;
    wire N__26677;
    wire N__26676;
    wire N__26675;
    wire N__26674;
    wire N__26673;
    wire N__26672;
    wire N__26671;
    wire N__26670;
    wire N__26667;
    wire N__26658;
    wire N__26655;
    wire N__26652;
    wire N__26649;
    wire N__26648;
    wire N__26641;
    wire N__26640;
    wire N__26639;
    wire N__26638;
    wire N__26631;
    wire N__26628;
    wire N__26621;
    wire N__26614;
    wire N__26611;
    wire N__26608;
    wire N__26605;
    wire N__26602;
    wire N__26599;
    wire N__26596;
    wire N__26593;
    wire N__26590;
    wire N__26587;
    wire N__26584;
    wire N__26581;
    wire N__26578;
    wire N__26577;
    wire N__26574;
    wire N__26571;
    wire N__26566;
    wire N__26563;
    wire N__26562;
    wire N__26557;
    wire N__26556;
    wire N__26555;
    wire N__26552;
    wire N__26547;
    wire N__26542;
    wire N__26539;
    wire N__26536;
    wire N__26533;
    wire N__26530;
    wire N__26527;
    wire N__26524;
    wire N__26521;
    wire N__26518;
    wire N__26515;
    wire N__26512;
    wire N__26509;
    wire N__26506;
    wire N__26503;
    wire N__26500;
    wire N__26497;
    wire N__26494;
    wire N__26491;
    wire N__26488;
    wire N__26485;
    wire N__26482;
    wire N__26479;
    wire N__26476;
    wire N__26473;
    wire N__26470;
    wire N__26467;
    wire N__26464;
    wire N__26461;
    wire N__26460;
    wire N__26459;
    wire N__26458;
    wire N__26457;
    wire N__26454;
    wire N__26447;
    wire N__26446;
    wire N__26443;
    wire N__26442;
    wire N__26441;
    wire N__26440;
    wire N__26439;
    wire N__26436;
    wire N__26433;
    wire N__26430;
    wire N__26419;
    wire N__26410;
    wire N__26407;
    wire N__26404;
    wire N__26401;
    wire N__26400;
    wire N__26397;
    wire N__26394;
    wire N__26389;
    wire N__26386;
    wire N__26385;
    wire N__26384;
    wire N__26381;
    wire N__26378;
    wire N__26375;
    wire N__26372;
    wire N__26367;
    wire N__26364;
    wire N__26361;
    wire N__26358;
    wire N__26353;
    wire N__26350;
    wire N__26347;
    wire N__26344;
    wire N__26341;
    wire N__26338;
    wire N__26335;
    wire N__26332;
    wire N__26329;
    wire N__26326;
    wire N__26323;
    wire N__26320;
    wire N__26317;
    wire N__26314;
    wire N__26311;
    wire N__26308;
    wire N__26305;
    wire N__26302;
    wire N__26299;
    wire N__26296;
    wire N__26293;
    wire N__26290;
    wire N__26287;
    wire N__26284;
    wire N__26281;
    wire N__26278;
    wire N__26275;
    wire N__26272;
    wire N__26269;
    wire N__26266;
    wire N__26263;
    wire N__26260;
    wire N__26257;
    wire N__26254;
    wire N__26251;
    wire N__26248;
    wire N__26245;
    wire N__26242;
    wire N__26239;
    wire N__26236;
    wire N__26233;
    wire N__26230;
    wire N__26227;
    wire N__26224;
    wire N__26221;
    wire N__26218;
    wire N__26217;
    wire N__26216;
    wire N__26215;
    wire N__26212;
    wire N__26211;
    wire N__26208;
    wire N__26207;
    wire N__26204;
    wire N__26191;
    wire N__26188;
    wire N__26185;
    wire N__26182;
    wire N__26179;
    wire N__26178;
    wire N__26177;
    wire N__26174;
    wire N__26171;
    wire N__26168;
    wire N__26161;
    wire N__26158;
    wire N__26155;
    wire N__26152;
    wire N__26149;
    wire N__26146;
    wire N__26143;
    wire N__26140;
    wire N__26137;
    wire N__26134;
    wire N__26131;
    wire N__26128;
    wire N__26125;
    wire N__26122;
    wire N__26119;
    wire N__26116;
    wire N__26113;
    wire N__26110;
    wire N__26107;
    wire N__26104;
    wire N__26103;
    wire N__26100;
    wire N__26097;
    wire N__26096;
    wire N__26095;
    wire N__26092;
    wire N__26087;
    wire N__26084;
    wire N__26079;
    wire N__26074;
    wire N__26071;
    wire N__26068;
    wire N__26065;
    wire N__26062;
    wire N__26061;
    wire N__26058;
    wire N__26055;
    wire N__26052;
    wire N__26051;
    wire N__26048;
    wire N__26045;
    wire N__26042;
    wire N__26041;
    wire N__26038;
    wire N__26035;
    wire N__26032;
    wire N__26029;
    wire N__26020;
    wire N__26017;
    wire N__26014;
    wire N__26011;
    wire N__26008;
    wire N__26005;
    wire N__26002;
    wire N__25999;
    wire N__25996;
    wire N__25993;
    wire N__25990;
    wire N__25987;
    wire N__25984;
    wire N__25983;
    wire N__25978;
    wire N__25977;
    wire N__25976;
    wire N__25975;
    wire N__25974;
    wire N__25971;
    wire N__25968;
    wire N__25961;
    wire N__25954;
    wire N__25951;
    wire N__25948;
    wire N__25945;
    wire N__25942;
    wire N__25939;
    wire N__25936;
    wire N__25933;
    wire N__25930;
    wire N__25927;
    wire N__25924;
    wire N__25921;
    wire N__25918;
    wire N__25915;
    wire N__25912;
    wire N__25909;
    wire N__25906;
    wire N__25903;
    wire N__25900;
    wire N__25897;
    wire N__25894;
    wire N__25891;
    wire N__25888;
    wire N__25885;
    wire N__25882;
    wire N__25879;
    wire N__25876;
    wire N__25873;
    wire N__25870;
    wire N__25867;
    wire N__25864;
    wire N__25861;
    wire N__25858;
    wire N__25855;
    wire N__25852;
    wire N__25849;
    wire N__25846;
    wire N__25843;
    wire N__25840;
    wire N__25837;
    wire N__25834;
    wire N__25831;
    wire N__25828;
    wire N__25825;
    wire N__25822;
    wire N__25819;
    wire N__25816;
    wire N__25815;
    wire N__25814;
    wire N__25809;
    wire N__25808;
    wire N__25807;
    wire N__25806;
    wire N__25803;
    wire N__25800;
    wire N__25797;
    wire N__25792;
    wire N__25783;
    wire N__25782;
    wire N__25779;
    wire N__25778;
    wire N__25775;
    wire N__25774;
    wire N__25771;
    wire N__25768;
    wire N__25763;
    wire N__25758;
    wire N__25755;
    wire N__25750;
    wire N__25747;
    wire N__25744;
    wire N__25741;
    wire N__25738;
    wire N__25737;
    wire N__25734;
    wire N__25731;
    wire N__25730;
    wire N__25725;
    wire N__25722;
    wire N__25719;
    wire N__25714;
    wire N__25711;
    wire N__25708;
    wire N__25705;
    wire N__25704;
    wire N__25701;
    wire N__25698;
    wire N__25695;
    wire N__25690;
    wire N__25687;
    wire N__25684;
    wire N__25681;
    wire N__25680;
    wire N__25677;
    wire N__25674;
    wire N__25671;
    wire N__25668;
    wire N__25663;
    wire N__25662;
    wire N__25661;
    wire N__25660;
    wire N__25659;
    wire N__25658;
    wire N__25657;
    wire N__25656;
    wire N__25655;
    wire N__25654;
    wire N__25653;
    wire N__25652;
    wire N__25645;
    wire N__25644;
    wire N__25643;
    wire N__25642;
    wire N__25641;
    wire N__25640;
    wire N__25639;
    wire N__25638;
    wire N__25637;
    wire N__25634;
    wire N__25633;
    wire N__25632;
    wire N__25631;
    wire N__25626;
    wire N__25613;
    wire N__25610;
    wire N__25593;
    wire N__25588;
    wire N__25587;
    wire N__25582;
    wire N__25577;
    wire N__25574;
    wire N__25569;
    wire N__25566;
    wire N__25555;
    wire N__25554;
    wire N__25553;
    wire N__25552;
    wire N__25551;
    wire N__25550;
    wire N__25549;
    wire N__25548;
    wire N__25547;
    wire N__25544;
    wire N__25541;
    wire N__25538;
    wire N__25535;
    wire N__25534;
    wire N__25533;
    wire N__25532;
    wire N__25531;
    wire N__25530;
    wire N__25529;
    wire N__25524;
    wire N__25517;
    wire N__25516;
    wire N__25515;
    wire N__25514;
    wire N__25513;
    wire N__25512;
    wire N__25511;
    wire N__25510;
    wire N__25509;
    wire N__25500;
    wire N__25487;
    wire N__25482;
    wire N__25477;
    wire N__25476;
    wire N__25471;
    wire N__25462;
    wire N__25455;
    wire N__25452;
    wire N__25449;
    wire N__25438;
    wire N__25437;
    wire N__25436;
    wire N__25435;
    wire N__25434;
    wire N__25433;
    wire N__25432;
    wire N__25431;
    wire N__25430;
    wire N__25429;
    wire N__25428;
    wire N__25427;
    wire N__25424;
    wire N__25421;
    wire N__25420;
    wire N__25419;
    wire N__25418;
    wire N__25417;
    wire N__25414;
    wire N__25411;
    wire N__25408;
    wire N__25405;
    wire N__25402;
    wire N__25399;
    wire N__25396;
    wire N__25393;
    wire N__25390;
    wire N__25389;
    wire N__25388;
    wire N__25387;
    wire N__25386;
    wire N__25385;
    wire N__25382;
    wire N__25375;
    wire N__25374;
    wire N__25373;
    wire N__25360;
    wire N__25355;
    wire N__25338;
    wire N__25333;
    wire N__25330;
    wire N__25325;
    wire N__25324;
    wire N__25321;
    wire N__25314;
    wire N__25309;
    wire N__25306;
    wire N__25301;
    wire N__25298;
    wire N__25291;
    wire N__25288;
    wire N__25285;
    wire N__25282;
    wire N__25279;
    wire N__25276;
    wire N__25275;
    wire N__25272;
    wire N__25269;
    wire N__25264;
    wire N__25261;
    wire N__25258;
    wire N__25255;
    wire N__25252;
    wire N__25249;
    wire N__25246;
    wire N__25243;
    wire N__25240;
    wire N__25237;
    wire N__25234;
    wire N__25231;
    wire N__25228;
    wire N__25225;
    wire N__25222;
    wire N__25219;
    wire N__25216;
    wire N__25213;
    wire N__25210;
    wire N__25207;
    wire N__25204;
    wire N__25201;
    wire N__25198;
    wire N__25195;
    wire N__25192;
    wire N__25191;
    wire N__25190;
    wire N__25189;
    wire N__25186;
    wire N__25183;
    wire N__25180;
    wire N__25177;
    wire N__25176;
    wire N__25173;
    wire N__25170;
    wire N__25167;
    wire N__25164;
    wire N__25161;
    wire N__25158;
    wire N__25155;
    wire N__25152;
    wire N__25147;
    wire N__25138;
    wire N__25135;
    wire N__25134;
    wire N__25133;
    wire N__25132;
    wire N__25129;
    wire N__25126;
    wire N__25123;
    wire N__25120;
    wire N__25117;
    wire N__25114;
    wire N__25111;
    wire N__25110;
    wire N__25109;
    wire N__25104;
    wire N__25099;
    wire N__25096;
    wire N__25093;
    wire N__25084;
    wire N__25081;
    wire N__25078;
    wire N__25075;
    wire N__25072;
    wire N__25069;
    wire N__25066;
    wire N__25063;
    wire N__25060;
    wire N__25057;
    wire N__25054;
    wire N__25051;
    wire N__25048;
    wire N__25045;
    wire N__25042;
    wire N__25039;
    wire N__25036;
    wire N__25033;
    wire N__25030;
    wire N__25027;
    wire N__25024;
    wire N__25021;
    wire N__25018;
    wire N__25015;
    wire N__25012;
    wire N__25009;
    wire N__25006;
    wire N__25003;
    wire N__25000;
    wire N__24997;
    wire N__24994;
    wire N__24991;
    wire N__24988;
    wire N__24985;
    wire N__24984;
    wire N__24981;
    wire N__24978;
    wire N__24973;
    wire N__24970;
    wire N__24967;
    wire N__24966;
    wire N__24963;
    wire N__24960;
    wire N__24955;
    wire N__24952;
    wire N__24949;
    wire N__24948;
    wire N__24945;
    wire N__24942;
    wire N__24937;
    wire N__24934;
    wire N__24931;
    wire N__24928;
    wire N__24927;
    wire N__24924;
    wire N__24921;
    wire N__24918;
    wire N__24913;
    wire N__24910;
    wire N__24907;
    wire N__24906;
    wire N__24903;
    wire N__24900;
    wire N__24895;
    wire N__24892;
    wire N__24889;
    wire N__24888;
    wire N__24885;
    wire N__24882;
    wire N__24877;
    wire N__24874;
    wire N__24871;
    wire N__24870;
    wire N__24867;
    wire N__24864;
    wire N__24859;
    wire N__24856;
    wire N__24853;
    wire N__24850;
    wire N__24847;
    wire N__24846;
    wire N__24843;
    wire N__24840;
    wire N__24835;
    wire N__24832;
    wire N__24829;
    wire N__24826;
    wire N__24823;
    wire N__24820;
    wire N__24817;
    wire N__24814;
    wire N__24811;
    wire N__24810;
    wire N__24807;
    wire N__24804;
    wire N__24799;
    wire N__24796;
    wire N__24793;
    wire N__24790;
    wire N__24787;
    wire N__24786;
    wire N__24783;
    wire N__24780;
    wire N__24775;
    wire N__24772;
    wire N__24769;
    wire N__24766;
    wire N__24763;
    wire N__24762;
    wire N__24759;
    wire N__24756;
    wire N__24751;
    wire N__24748;
    wire N__24745;
    wire N__24744;
    wire N__24741;
    wire N__24738;
    wire N__24735;
    wire N__24730;
    wire N__24727;
    wire N__24724;
    wire N__24723;
    wire N__24720;
    wire N__24717;
    wire N__24712;
    wire N__24709;
    wire N__24706;
    wire N__24705;
    wire N__24702;
    wire N__24699;
    wire N__24694;
    wire N__24691;
    wire N__24688;
    wire N__24687;
    wire N__24684;
    wire N__24681;
    wire N__24676;
    wire N__24673;
    wire N__24670;
    wire N__24669;
    wire N__24666;
    wire N__24663;
    wire N__24658;
    wire N__24655;
    wire N__24652;
    wire N__24649;
    wire N__24646;
    wire N__24645;
    wire N__24642;
    wire N__24639;
    wire N__24634;
    wire N__24631;
    wire N__24628;
    wire N__24625;
    wire N__24624;
    wire N__24621;
    wire N__24618;
    wire N__24617;
    wire N__24616;
    wire N__24615;
    wire N__24614;
    wire N__24609;
    wire N__24608;
    wire N__24605;
    wire N__24602;
    wire N__24601;
    wire N__24600;
    wire N__24597;
    wire N__24594;
    wire N__24593;
    wire N__24590;
    wire N__24581;
    wire N__24578;
    wire N__24575;
    wire N__24570;
    wire N__24563;
    wire N__24558;
    wire N__24555;
    wire N__24552;
    wire N__24549;
    wire N__24546;
    wire N__24543;
    wire N__24540;
    wire N__24535;
    wire N__24534;
    wire N__24531;
    wire N__24528;
    wire N__24525;
    wire N__24524;
    wire N__24519;
    wire N__24516;
    wire N__24511;
    wire N__24508;
    wire N__24505;
    wire N__24502;
    wire N__24501;
    wire N__24498;
    wire N__24495;
    wire N__24490;
    wire N__24487;
    wire N__24484;
    wire N__24481;
    wire N__24478;
    wire N__24477;
    wire N__24474;
    wire N__24471;
    wire N__24466;
    wire N__24463;
    wire N__24460;
    wire N__24459;
    wire N__24456;
    wire N__24453;
    wire N__24450;
    wire N__24447;
    wire N__24442;
    wire N__24439;
    wire N__24436;
    wire N__24435;
    wire N__24430;
    wire N__24427;
    wire N__24424;
    wire N__24423;
    wire N__24420;
    wire N__24417;
    wire N__24412;
    wire N__24409;
    wire N__24408;
    wire N__24405;
    wire N__24402;
    wire N__24397;
    wire N__24394;
    wire N__24391;
    wire N__24390;
    wire N__24385;
    wire N__24382;
    wire N__24379;
    wire N__24376;
    wire N__24375;
    wire N__24372;
    wire N__24369;
    wire N__24364;
    wire N__24361;
    wire N__24360;
    wire N__24357;
    wire N__24354;
    wire N__24351;
    wire N__24346;
    wire N__24343;
    wire N__24342;
    wire N__24339;
    wire N__24336;
    wire N__24333;
    wire N__24328;
    wire N__24325;
    wire N__24324;
    wire N__24321;
    wire N__24318;
    wire N__24315;
    wire N__24312;
    wire N__24309;
    wire N__24304;
    wire N__24301;
    wire N__24298;
    wire N__24297;
    wire N__24294;
    wire N__24291;
    wire N__24288;
    wire N__24285;
    wire N__24280;
    wire N__24277;
    wire N__24276;
    wire N__24271;
    wire N__24268;
    wire N__24265;
    wire N__24262;
    wire N__24261;
    wire N__24256;
    wire N__24253;
    wire N__24250;
    wire N__24247;
    wire N__24244;
    wire N__24241;
    wire N__24238;
    wire N__24235;
    wire N__24234;
    wire N__24229;
    wire N__24226;
    wire N__24223;
    wire N__24222;
    wire N__24219;
    wire N__24216;
    wire N__24211;
    wire N__24208;
    wire N__24207;
    wire N__24204;
    wire N__24201;
    wire N__24198;
    wire N__24195;
    wire N__24190;
    wire N__24187;
    wire N__24186;
    wire N__24183;
    wire N__24180;
    wire N__24177;
    wire N__24172;
    wire N__24169;
    wire N__24166;
    wire N__24165;
    wire N__24162;
    wire N__24159;
    wire N__24156;
    wire N__24151;
    wire N__24148;
    wire N__24147;
    wire N__24142;
    wire N__24139;
    wire N__24136;
    wire N__24135;
    wire N__24132;
    wire N__24131;
    wire N__24130;
    wire N__24127;
    wire N__24124;
    wire N__24121;
    wire N__24118;
    wire N__24115;
    wire N__24110;
    wire N__24107;
    wire N__24104;
    wire N__24101;
    wire N__24098;
    wire N__24095;
    wire N__24092;
    wire N__24085;
    wire N__24082;
    wire N__24079;
    wire N__24078;
    wire N__24077;
    wire N__24074;
    wire N__24071;
    wire N__24068;
    wire N__24061;
    wire N__24058;
    wire N__24055;
    wire N__24052;
    wire N__24049;
    wire N__24048;
    wire N__24047;
    wire N__24044;
    wire N__24041;
    wire N__24038;
    wire N__24031;
    wire N__24028;
    wire N__24025;
    wire N__24022;
    wire N__24019;
    wire N__24018;
    wire N__24017;
    wire N__24014;
    wire N__24011;
    wire N__24008;
    wire N__24001;
    wire N__23998;
    wire N__23995;
    wire N__23992;
    wire N__23989;
    wire N__23986;
    wire N__23985;
    wire N__23984;
    wire N__23981;
    wire N__23978;
    wire N__23975;
    wire N__23968;
    wire N__23965;
    wire N__23962;
    wire N__23959;
    wire N__23956;
    wire N__23955;
    wire N__23952;
    wire N__23949;
    wire N__23948;
    wire N__23943;
    wire N__23940;
    wire N__23935;
    wire N__23932;
    wire N__23929;
    wire N__23926;
    wire N__23923;
    wire N__23920;
    wire N__23919;
    wire N__23916;
    wire N__23913;
    wire N__23908;
    wire N__23905;
    wire N__23904;
    wire N__23899;
    wire N__23896;
    wire N__23893;
    wire N__23890;
    wire N__23887;
    wire N__23884;
    wire N__23881;
    wire N__23880;
    wire N__23877;
    wire N__23874;
    wire N__23873;
    wire N__23868;
    wire N__23865;
    wire N__23864;
    wire N__23859;
    wire N__23856;
    wire N__23853;
    wire N__23848;
    wire N__23845;
    wire N__23842;
    wire N__23839;
    wire N__23836;
    wire N__23833;
    wire N__23830;
    wire N__23827;
    wire N__23824;
    wire N__23821;
    wire N__23818;
    wire N__23815;
    wire N__23812;
    wire N__23809;
    wire N__23806;
    wire N__23803;
    wire N__23800;
    wire N__23797;
    wire N__23794;
    wire N__23791;
    wire N__23788;
    wire N__23785;
    wire N__23782;
    wire N__23779;
    wire N__23776;
    wire N__23773;
    wire N__23770;
    wire N__23767;
    wire N__23764;
    wire N__23761;
    wire N__23758;
    wire N__23755;
    wire N__23752;
    wire N__23751;
    wire N__23748;
    wire N__23745;
    wire N__23744;
    wire N__23739;
    wire N__23736;
    wire N__23731;
    wire N__23728;
    wire N__23725;
    wire N__23722;
    wire N__23721;
    wire N__23718;
    wire N__23715;
    wire N__23712;
    wire N__23707;
    wire N__23704;
    wire N__23701;
    wire N__23698;
    wire N__23697;
    wire N__23694;
    wire N__23691;
    wire N__23688;
    wire N__23683;
    wire N__23680;
    wire N__23677;
    wire N__23674;
    wire N__23671;
    wire N__23668;
    wire N__23665;
    wire N__23664;
    wire N__23661;
    wire N__23658;
    wire N__23653;
    wire N__23650;
    wire N__23647;
    wire N__23644;
    wire N__23641;
    wire N__23638;
    wire N__23635;
    wire N__23634;
    wire N__23631;
    wire N__23628;
    wire N__23625;
    wire N__23620;
    wire N__23617;
    wire N__23614;
    wire N__23611;
    wire N__23610;
    wire N__23607;
    wire N__23604;
    wire N__23601;
    wire N__23596;
    wire N__23593;
    wire N__23590;
    wire N__23587;
    wire N__23586;
    wire N__23583;
    wire N__23580;
    wire N__23577;
    wire N__23572;
    wire N__23569;
    wire N__23566;
    wire N__23563;
    wire N__23560;
    wire N__23557;
    wire N__23554;
    wire N__23553;
    wire N__23550;
    wire N__23547;
    wire N__23542;
    wire N__23539;
    wire N__23536;
    wire N__23533;
    wire N__23530;
    wire N__23527;
    wire N__23524;
    wire N__23521;
    wire N__23518;
    wire N__23517;
    wire N__23514;
    wire N__23511;
    wire N__23508;
    wire N__23503;
    wire N__23500;
    wire N__23497;
    wire N__23494;
    wire N__23493;
    wire N__23490;
    wire N__23487;
    wire N__23484;
    wire N__23479;
    wire N__23476;
    wire N__23473;
    wire N__23470;
    wire N__23467;
    wire N__23466;
    wire N__23463;
    wire N__23460;
    wire N__23457;
    wire N__23454;
    wire N__23449;
    wire N__23446;
    wire N__23443;
    wire N__23440;
    wire N__23439;
    wire N__23436;
    wire N__23433;
    wire N__23430;
    wire N__23425;
    wire N__23422;
    wire N__23419;
    wire N__23416;
    wire N__23413;
    wire N__23410;
    wire N__23407;
    wire N__23404;
    wire N__23401;
    wire N__23398;
    wire N__23395;
    wire N__23392;
    wire N__23389;
    wire N__23386;
    wire N__23383;
    wire N__23380;
    wire N__23377;
    wire N__23376;
    wire N__23375;
    wire N__23372;
    wire N__23369;
    wire N__23366;
    wire N__23363;
    wire N__23360;
    wire N__23353;
    wire N__23350;
    wire N__23349;
    wire N__23346;
    wire N__23343;
    wire N__23340;
    wire N__23335;
    wire N__23332;
    wire N__23329;
    wire N__23326;
    wire N__23325;
    wire N__23322;
    wire N__23319;
    wire N__23316;
    wire N__23313;
    wire N__23310;
    wire N__23305;
    wire N__23302;
    wire N__23299;
    wire N__23296;
    wire N__23293;
    wire N__23292;
    wire N__23289;
    wire N__23286;
    wire N__23283;
    wire N__23278;
    wire N__23275;
    wire N__23272;
    wire N__23269;
    wire N__23268;
    wire N__23265;
    wire N__23262;
    wire N__23257;
    wire N__23254;
    wire N__23251;
    wire N__23248;
    wire N__23245;
    wire N__23242;
    wire N__23239;
    wire N__23236;
    wire N__23233;
    wire N__23230;
    wire N__23227;
    wire N__23224;
    wire N__23221;
    wire N__23218;
    wire N__23215;
    wire N__23212;
    wire N__23209;
    wire N__23206;
    wire N__23203;
    wire N__23200;
    wire N__23197;
    wire N__23194;
    wire N__23191;
    wire N__23188;
    wire N__23185;
    wire N__23182;
    wire N__23179;
    wire N__23176;
    wire N__23173;
    wire N__23170;
    wire N__23167;
    wire N__23164;
    wire N__23161;
    wire N__23158;
    wire N__23155;
    wire N__23152;
    wire N__23149;
    wire N__23146;
    wire N__23143;
    wire N__23140;
    wire N__23137;
    wire N__23134;
    wire N__23131;
    wire N__23128;
    wire N__23125;
    wire N__23122;
    wire N__23119;
    wire N__23116;
    wire N__23113;
    wire N__23110;
    wire N__23107;
    wire N__23104;
    wire N__23101;
    wire N__23098;
    wire N__23095;
    wire N__23092;
    wire N__23089;
    wire N__23086;
    wire N__23083;
    wire N__23080;
    wire N__23077;
    wire N__23074;
    wire N__23071;
    wire N__23068;
    wire N__23065;
    wire N__23062;
    wire N__23059;
    wire N__23056;
    wire N__23053;
    wire N__23050;
    wire N__23047;
    wire N__23044;
    wire N__23041;
    wire N__23038;
    wire N__23035;
    wire N__23034;
    wire N__23033;
    wire N__23030;
    wire N__23027;
    wire N__23024;
    wire N__23017;
    wire N__23014;
    wire N__23011;
    wire N__23008;
    wire N__23005;
    wire N__23002;
    wire N__22999;
    wire N__22996;
    wire N__22993;
    wire N__22990;
    wire N__22987;
    wire N__22984;
    wire N__22981;
    wire N__22978;
    wire N__22975;
    wire N__22972;
    wire N__22969;
    wire N__22966;
    wire N__22963;
    wire N__22960;
    wire N__22957;
    wire N__22954;
    wire N__22951;
    wire N__22948;
    wire N__22945;
    wire N__22942;
    wire N__22939;
    wire N__22936;
    wire N__22933;
    wire N__22930;
    wire N__22927;
    wire N__22924;
    wire N__22921;
    wire N__22918;
    wire N__22915;
    wire N__22912;
    wire N__22909;
    wire N__22906;
    wire N__22903;
    wire N__22900;
    wire N__22897;
    wire N__22894;
    wire N__22891;
    wire N__22888;
    wire N__22885;
    wire N__22882;
    wire N__22879;
    wire N__22876;
    wire N__22873;
    wire N__22870;
    wire N__22867;
    wire N__22864;
    wire N__22861;
    wire N__22858;
    wire N__22855;
    wire N__22852;
    wire N__22849;
    wire N__22846;
    wire N__22843;
    wire N__22840;
    wire N__22837;
    wire N__22834;
    wire N__22831;
    wire N__22828;
    wire N__22825;
    wire N__22822;
    wire N__22821;
    wire N__22820;
    wire N__22817;
    wire N__22816;
    wire N__22815;
    wire N__22814;
    wire N__22813;
    wire N__22812;
    wire N__22807;
    wire N__22800;
    wire N__22797;
    wire N__22792;
    wire N__22789;
    wire N__22786;
    wire N__22781;
    wire N__22778;
    wire N__22775;
    wire N__22772;
    wire N__22769;
    wire N__22766;
    wire N__22763;
    wire N__22756;
    wire N__22753;
    wire N__22750;
    wire N__22747;
    wire N__22746;
    wire N__22745;
    wire N__22744;
    wire N__22743;
    wire N__22742;
    wire N__22735;
    wire N__22730;
    wire N__22727;
    wire N__22726;
    wire N__22723;
    wire N__22718;
    wire N__22715;
    wire N__22712;
    wire N__22707;
    wire N__22704;
    wire N__22701;
    wire N__22696;
    wire N__22693;
    wire N__22690;
    wire N__22687;
    wire N__22686;
    wire N__22685;
    wire N__22682;
    wire N__22679;
    wire N__22676;
    wire N__22675;
    wire N__22670;
    wire N__22667;
    wire N__22664;
    wire N__22657;
    wire N__22654;
    wire N__22651;
    wire N__22648;
    wire N__22645;
    wire N__22642;
    wire N__22639;
    wire N__22636;
    wire N__22633;
    wire N__22630;
    wire N__22629;
    wire N__22626;
    wire N__22625;
    wire N__22622;
    wire N__22619;
    wire N__22616;
    wire N__22613;
    wire N__22610;
    wire N__22603;
    wire N__22600;
    wire N__22597;
    wire N__22594;
    wire N__22591;
    wire N__22588;
    wire N__22587;
    wire N__22584;
    wire N__22581;
    wire N__22580;
    wire N__22575;
    wire N__22572;
    wire N__22569;
    wire N__22566;
    wire N__22563;
    wire N__22558;
    wire N__22557;
    wire N__22556;
    wire N__22553;
    wire N__22550;
    wire N__22547;
    wire N__22544;
    wire N__22537;
    wire N__22536;
    wire N__22533;
    wire N__22530;
    wire N__22527;
    wire N__22522;
    wire N__22519;
    wire N__22516;
    wire N__22513;
    wire N__22510;
    wire N__22507;
    wire N__22504;
    wire N__22501;
    wire N__22498;
    wire N__22495;
    wire N__22492;
    wire N__22491;
    wire N__22488;
    wire N__22485;
    wire N__22482;
    wire N__22479;
    wire N__22476;
    wire N__22471;
    wire N__22470;
    wire N__22469;
    wire N__22466;
    wire N__22463;
    wire N__22460;
    wire N__22453;
    wire N__22450;
    wire N__22447;
    wire N__22446;
    wire N__22445;
    wire N__22440;
    wire N__22437;
    wire N__22432;
    wire N__22431;
    wire N__22426;
    wire N__22423;
    wire N__22420;
    wire N__22417;
    wire N__22414;
    wire N__22411;
    wire N__22408;
    wire N__22405;
    wire N__22402;
    wire N__22399;
    wire N__22396;
    wire N__22393;
    wire N__22390;
    wire N__22387;
    wire N__22384;
    wire N__22381;
    wire N__22378;
    wire N__22375;
    wire N__22372;
    wire N__22369;
    wire N__22366;
    wire N__22363;
    wire N__22360;
    wire N__22357;
    wire N__22354;
    wire N__22351;
    wire N__22348;
    wire N__22345;
    wire N__22342;
    wire N__22339;
    wire N__22336;
    wire N__22333;
    wire N__22332;
    wire N__22329;
    wire N__22326;
    wire N__22321;
    wire N__22318;
    wire N__22317;
    wire N__22316;
    wire N__22313;
    wire N__22310;
    wire N__22307;
    wire N__22304;
    wire N__22299;
    wire N__22294;
    wire N__22291;
    wire N__22288;
    wire N__22285;
    wire N__22282;
    wire N__22279;
    wire N__22276;
    wire N__22273;
    wire N__22272;
    wire N__22269;
    wire N__22266;
    wire N__22261;
    wire N__22260;
    wire N__22259;
    wire N__22254;
    wire N__22251;
    wire N__22248;
    wire N__22245;
    wire N__22242;
    wire N__22239;
    wire N__22236;
    wire N__22233;
    wire N__22230;
    wire N__22227;
    wire N__22222;
    wire N__22219;
    wire N__22216;
    wire N__22213;
    wire N__22210;
    wire N__22207;
    wire N__22204;
    wire N__22201;
    wire N__22198;
    wire N__22197;
    wire N__22196;
    wire N__22193;
    wire N__22190;
    wire N__22187;
    wire N__22182;
    wire N__22177;
    wire N__22174;
    wire N__22171;
    wire N__22170;
    wire N__22169;
    wire N__22166;
    wire N__22163;
    wire N__22160;
    wire N__22155;
    wire N__22150;
    wire N__22147;
    wire N__22144;
    wire N__22141;
    wire N__22138;
    wire N__22135;
    wire N__22132;
    wire N__22129;
    wire N__22126;
    wire N__22125;
    wire N__22124;
    wire N__22121;
    wire N__22118;
    wire N__22115;
    wire N__22112;
    wire N__22109;
    wire N__22102;
    wire N__22099;
    wire N__22096;
    wire N__22093;
    wire N__22090;
    wire N__22087;
    wire N__22084;
    wire N__22081;
    wire N__22080;
    wire N__22079;
    wire N__22076;
    wire N__22073;
    wire N__22070;
    wire N__22067;
    wire N__22064;
    wire N__22057;
    wire N__22054;
    wire N__22051;
    wire N__22048;
    wire N__22045;
    wire N__22042;
    wire N__22041;
    wire N__22040;
    wire N__22037;
    wire N__22034;
    wire N__22031;
    wire N__22028;
    wire N__22021;
    wire N__22018;
    wire N__22015;
    wire N__22012;
    wire N__22009;
    wire N__22006;
    wire N__22003;
    wire N__22000;
    wire N__21997;
    wire N__21994;
    wire N__21991;
    wire N__21988;
    wire N__21987;
    wire N__21986;
    wire N__21985;
    wire N__21984;
    wire N__21983;
    wire N__21982;
    wire N__21981;
    wire N__21980;
    wire N__21979;
    wire N__21970;
    wire N__21961;
    wire N__21956;
    wire N__21951;
    wire N__21946;
    wire N__21943;
    wire N__21940;
    wire N__21937;
    wire N__21934;
    wire N__21931;
    wire N__21928;
    wire N__21925;
    wire N__21924;
    wire N__21923;
    wire N__21920;
    wire N__21917;
    wire N__21914;
    wire N__21911;
    wire N__21908;
    wire N__21901;
    wire N__21898;
    wire N__21895;
    wire N__21892;
    wire N__21889;
    wire N__21886;
    wire N__21885;
    wire N__21884;
    wire N__21881;
    wire N__21878;
    wire N__21875;
    wire N__21872;
    wire N__21869;
    wire N__21862;
    wire N__21859;
    wire N__21856;
    wire N__21853;
    wire N__21850;
    wire N__21847;
    wire N__21846;
    wire N__21845;
    wire N__21842;
    wire N__21839;
    wire N__21836;
    wire N__21831;
    wire N__21826;
    wire N__21823;
    wire N__21820;
    wire N__21817;
    wire N__21814;
    wire N__21811;
    wire N__21810;
    wire N__21809;
    wire N__21806;
    wire N__21803;
    wire N__21800;
    wire N__21795;
    wire N__21790;
    wire N__21787;
    wire N__21784;
    wire N__21781;
    wire N__21778;
    wire N__21775;
    wire N__21772;
    wire N__21769;
    wire N__21766;
    wire N__21765;
    wire N__21764;
    wire N__21761;
    wire N__21758;
    wire N__21755;
    wire N__21750;
    wire N__21745;
    wire N__21742;
    wire N__21739;
    wire N__21736;
    wire N__21733;
    wire N__21730;
    wire N__21727;
    wire N__21724;
    wire N__21721;
    wire N__21718;
    wire N__21715;
    wire N__21712;
    wire N__21709;
    wire N__21706;
    wire N__21703;
    wire N__21700;
    wire N__21697;
    wire N__21694;
    wire N__21691;
    wire N__21688;
    wire N__21685;
    wire N__21682;
    wire N__21679;
    wire N__21676;
    wire N__21673;
    wire N__21670;
    wire N__21667;
    wire N__21664;
    wire N__21661;
    wire N__21658;
    wire N__21655;
    wire N__21652;
    wire N__21649;
    wire N__21646;
    wire N__21643;
    wire N__21640;
    wire N__21637;
    wire N__21634;
    wire N__21631;
    wire N__21628;
    wire N__21627;
    wire N__21626;
    wire N__21625;
    wire N__21624;
    wire N__21621;
    wire N__21620;
    wire N__21617;
    wire N__21614;
    wire N__21613;
    wire N__21612;
    wire N__21611;
    wire N__21610;
    wire N__21609;
    wire N__21608;
    wire N__21607;
    wire N__21606;
    wire N__21605;
    wire N__21604;
    wire N__21603;
    wire N__21602;
    wire N__21601;
    wire N__21600;
    wire N__21599;
    wire N__21598;
    wire N__21597;
    wire N__21596;
    wire N__21595;
    wire N__21594;
    wire N__21589;
    wire N__21586;
    wire N__21583;
    wire N__21578;
    wire N__21569;
    wire N__21568;
    wire N__21551;
    wire N__21548;
    wire N__21533;
    wire N__21530;
    wire N__21521;
    wire N__21518;
    wire N__21515;
    wire N__21510;
    wire N__21509;
    wire N__21508;
    wire N__21507;
    wire N__21506;
    wire N__21505;
    wire N__21500;
    wire N__21497;
    wire N__21492;
    wire N__21487;
    wire N__21480;
    wire N__21469;
    wire N__21468;
    wire N__21467;
    wire N__21466;
    wire N__21465;
    wire N__21464;
    wire N__21463;
    wire N__21462;
    wire N__21461;
    wire N__21448;
    wire N__21445;
    wire N__21444;
    wire N__21439;
    wire N__21436;
    wire N__21431;
    wire N__21428;
    wire N__21423;
    wire N__21418;
    wire N__21417;
    wire N__21416;
    wire N__21415;
    wire N__21414;
    wire N__21413;
    wire N__21410;
    wire N__21407;
    wire N__21406;
    wire N__21405;
    wire N__21402;
    wire N__21399;
    wire N__21396;
    wire N__21395;
    wire N__21394;
    wire N__21389;
    wire N__21376;
    wire N__21371;
    wire N__21368;
    wire N__21363;
    wire N__21360;
    wire N__21357;
    wire N__21352;
    wire N__21349;
    wire N__21346;
    wire N__21343;
    wire N__21340;
    wire N__21337;
    wire N__21334;
    wire N__21331;
    wire N__21328;
    wire N__21325;
    wire N__21322;
    wire N__21319;
    wire N__21316;
    wire N__21313;
    wire N__21310;
    wire N__21307;
    wire N__21304;
    wire N__21303;
    wire N__21302;
    wire N__21299;
    wire N__21298;
    wire N__21297;
    wire N__21296;
    wire N__21295;
    wire N__21294;
    wire N__21293;
    wire N__21292;
    wire N__21291;
    wire N__21290;
    wire N__21287;
    wire N__21284;
    wire N__21281;
    wire N__21272;
    wire N__21263;
    wire N__21260;
    wire N__21253;
    wire N__21246;
    wire N__21243;
    wire N__21240;
    wire N__21235;
    wire N__21232;
    wire N__21229;
    wire N__21226;
    wire N__21223;
    wire N__21220;
    wire N__21217;
    wire N__21214;
    wire N__21211;
    wire N__21208;
    wire N__21205;
    wire N__21202;
    wire N__21199;
    wire N__21196;
    wire N__21193;
    wire N__21190;
    wire N__21187;
    wire N__21184;
    wire N__21181;
    wire N__21180;
    wire N__21179;
    wire N__21174;
    wire N__21171;
    wire N__21168;
    wire N__21163;
    wire N__21160;
    wire N__21157;
    wire N__21154;
    wire N__21151;
    wire N__21148;
    wire N__21145;
    wire N__21142;
    wire N__21139;
    wire N__21136;
    wire N__21133;
    wire N__21130;
    wire N__21127;
    wire N__21124;
    wire N__21121;
    wire N__21118;
    wire N__21115;
    wire N__21112;
    wire N__21109;
    wire N__21106;
    wire N__21103;
    wire N__21100;
    wire N__21097;
    wire N__21094;
    wire N__21091;
    wire N__21088;
    wire N__21085;
    wire N__21082;
    wire N__21079;
    wire N__21076;
    wire N__21073;
    wire N__21070;
    wire N__21067;
    wire N__21064;
    wire N__21061;
    wire N__21058;
    wire N__21055;
    wire N__21052;
    wire N__21049;
    wire N__21046;
    wire N__21043;
    wire N__21040;
    wire N__21037;
    wire N__21036;
    wire N__21035;
    wire N__21034;
    wire N__21033;
    wire N__21030;
    wire N__21027;
    wire N__21026;
    wire N__21023;
    wire N__21022;
    wire N__21019;
    wire N__21018;
    wire N__21015;
    wire N__21012;
    wire N__20999;
    wire N__20992;
    wire N__20989;
    wire N__20986;
    wire N__20983;
    wire N__20980;
    wire N__20977;
    wire N__20974;
    wire N__20971;
    wire N__20968;
    wire N__20965;
    wire N__20962;
    wire N__20959;
    wire N__20956;
    wire N__20953;
    wire N__20950;
    wire N__20947;
    wire N__20944;
    wire N__20941;
    wire N__20938;
    wire N__20935;
    wire N__20934;
    wire N__20933;
    wire N__20930;
    wire N__20927;
    wire N__20924;
    wire N__20919;
    wire N__20916;
    wire N__20911;
    wire N__20908;
    wire N__20905;
    wire N__20902;
    wire N__20901;
    wire N__20900;
    wire N__20897;
    wire N__20894;
    wire N__20891;
    wire N__20888;
    wire N__20883;
    wire N__20880;
    wire N__20875;
    wire N__20872;
    wire N__20869;
    wire N__20866;
    wire N__20863;
    wire N__20860;
    wire N__20857;
    wire N__20854;
    wire N__20851;
    wire N__20848;
    wire N__20845;
    wire N__20842;
    wire N__20839;
    wire N__20836;
    wire N__20833;
    wire N__20830;
    wire N__20827;
    wire N__20824;
    wire N__20821;
    wire N__20818;
    wire N__20815;
    wire N__20812;
    wire N__20809;
    wire N__20806;
    wire N__20803;
    wire N__20800;
    wire N__20797;
    wire N__20794;
    wire N__20791;
    wire N__20788;
    wire N__20785;
    wire N__20782;
    wire N__20779;
    wire N__20776;
    wire N__20773;
    wire N__20770;
    wire N__20767;
    wire N__20764;
    wire N__20761;
    wire N__20758;
    wire N__20755;
    wire N__20752;
    wire N__20749;
    wire N__20746;
    wire N__20743;
    wire N__20740;
    wire N__20737;
    wire N__20734;
    wire N__20731;
    wire N__20728;
    wire N__20725;
    wire N__20722;
    wire N__20719;
    wire N__20716;
    wire N__20713;
    wire N__20710;
    wire N__20707;
    wire N__20704;
    wire N__20701;
    wire N__20698;
    wire N__20695;
    wire N__20692;
    wire N__20689;
    wire N__20686;
    wire N__20683;
    wire N__20680;
    wire N__20677;
    wire N__20674;
    wire N__20671;
    wire N__20668;
    wire N__20665;
    wire N__20662;
    wire N__20659;
    wire N__20656;
    wire N__20653;
    wire N__20650;
    wire N__20647;
    wire N__20644;
    wire N__20641;
    wire N__20638;
    wire N__20635;
    wire N__20632;
    wire N__20631;
    wire N__20628;
    wire N__20625;
    wire N__20620;
    wire N__20619;
    wire N__20614;
    wire N__20611;
    wire N__20608;
    wire N__20605;
    wire N__20602;
    wire N__20599;
    wire N__20596;
    wire N__20593;
    wire N__20592;
    wire N__20589;
    wire N__20586;
    wire N__20581;
    wire N__20580;
    wire N__20577;
    wire N__20576;
    wire N__20573;
    wire N__20570;
    wire N__20567;
    wire N__20560;
    wire N__20557;
    wire N__20554;
    wire N__20551;
    wire N__20548;
    wire N__20545;
    wire N__20542;
    wire N__20539;
    wire N__20536;
    wire N__20533;
    wire N__20530;
    wire N__20527;
    wire N__20524;
    wire N__20521;
    wire N__20518;
    wire N__20515;
    wire N__20512;
    wire N__20509;
    wire N__20506;
    wire N__20503;
    wire N__20500;
    wire N__20497;
    wire N__20494;
    wire N__20491;
    wire N__20488;
    wire N__20485;
    wire N__20482;
    wire N__20479;
    wire N__20476;
    wire N__20473;
    wire N__20470;
    wire N__20467;
    wire N__20464;
    wire N__20461;
    wire N__20458;
    wire N__20455;
    wire N__20452;
    wire N__20449;
    wire N__20446;
    wire N__20443;
    wire N__20440;
    wire N__20437;
    wire N__20434;
    wire N__20431;
    wire N__20428;
    wire N__20425;
    wire N__20422;
    wire N__20419;
    wire N__20416;
    wire N__20413;
    wire N__20410;
    wire N__20407;
    wire N__20404;
    wire N__20401;
    wire N__20398;
    wire N__20395;
    wire N__20392;
    wire N__20389;
    wire N__20386;
    wire N__20383;
    wire N__20380;
    wire N__20377;
    wire N__20374;
    wire N__20373;
    wire N__20370;
    wire N__20367;
    wire N__20362;
    wire N__20359;
    wire N__20356;
    wire N__20353;
    wire N__20352;
    wire N__20349;
    wire N__20346;
    wire N__20341;
    wire N__20338;
    wire N__20337;
    wire N__20336;
    wire N__20333;
    wire N__20330;
    wire N__20327;
    wire N__20320;
    wire N__20317;
    wire N__20314;
    wire N__20311;
    wire N__20308;
    wire N__20307;
    wire N__20304;
    wire N__20301;
    wire N__20296;
    wire N__20293;
    wire N__20290;
    wire N__20289;
    wire N__20288;
    wire N__20285;
    wire N__20280;
    wire N__20275;
    wire N__20272;
    wire N__20271;
    wire N__20268;
    wire N__20265;
    wire N__20260;
    wire N__20259;
    wire N__20256;
    wire N__20253;
    wire N__20248;
    wire N__20247;
    wire N__20242;
    wire N__20239;
    wire N__20236;
    wire N__20233;
    wire N__20230;
    wire N__20229;
    wire N__20226;
    wire N__20223;
    wire N__20218;
    wire N__20217;
    wire N__20212;
    wire N__20209;
    wire N__20206;
    wire N__20203;
    wire N__20200;
    wire N__20197;
    wire N__20194;
    wire N__20191;
    wire N__20190;
    wire N__20189;
    wire N__20182;
    wire N__20179;
    wire N__20176;
    wire N__20173;
    wire N__20170;
    wire N__20167;
    wire N__20164;
    wire N__20161;
    wire N__20158;
    wire N__20155;
    wire N__20152;
    wire N__20151;
    wire N__20148;
    wire N__20145;
    wire N__20140;
    wire N__20139;
    wire N__20138;
    wire N__20135;
    wire N__20132;
    wire N__20129;
    wire N__20122;
    wire N__20119;
    wire N__20116;
    wire N__20113;
    wire N__20110;
    wire N__20107;
    wire N__20106;
    wire N__20103;
    wire N__20100;
    wire N__20095;
    wire N__20092;
    wire N__20089;
    wire N__20086;
    wire N__20083;
    wire N__20080;
    wire N__20079;
    wire N__20076;
    wire N__20073;
    wire N__20068;
    wire N__20065;
    wire N__20062;
    wire N__20059;
    wire N__20056;
    wire N__20053;
    wire N__20050;
    wire N__20049;
    wire N__20046;
    wire N__20043;
    wire N__20040;
    wire N__20035;
    wire N__20034;
    wire N__20031;
    wire N__20028;
    wire N__20025;
    wire N__20020;
    wire N__20019;
    wire N__20016;
    wire N__20013;
    wire N__20010;
    wire N__20005;
    wire N__20002;
    wire N__20001;
    wire N__20000;
    wire N__19995;
    wire N__19992;
    wire N__19987;
    wire N__19984;
    wire N__19983;
    wire N__19982;
    wire N__19979;
    wire N__19974;
    wire N__19971;
    wire N__19966;
    wire N__19965;
    wire N__19964;
    wire N__19961;
    wire N__19958;
    wire N__19955;
    wire N__19952;
    wire N__19945;
    wire N__19944;
    wire N__19943;
    wire N__19938;
    wire N__19935;
    wire N__19930;
    wire N__19927;
    wire N__19926;
    wire N__19925;
    wire N__19920;
    wire N__19917;
    wire N__19912;
    wire N__19909;
    wire N__19906;
    wire N__19903;
    wire N__19900;
    wire N__19897;
    wire N__19894;
    wire N__19891;
    wire N__19888;
    wire N__19885;
    wire N__19882;
    wire N__19879;
    wire N__19876;
    wire N__19873;
    wire N__19870;
    wire N__19867;
    wire N__19864;
    wire N__19861;
    wire N__19858;
    wire N__19855;
    wire N__19854;
    wire N__19851;
    wire N__19848;
    wire N__19843;
    wire N__19840;
    wire N__19837;
    wire N__19834;
    wire N__19831;
    wire N__19828;
    wire N__19825;
    wire N__19822;
    wire N__19819;
    wire N__19816;
    wire N__19813;
    wire N__19810;
    wire N__19807;
    wire N__19804;
    wire N__19801;
    wire N__19798;
    wire N__19795;
    wire N__19792;
    wire N__19789;
    wire N__19786;
    wire N__19783;
    wire N__19780;
    wire N__19777;
    wire N__19774;
    wire N__19771;
    wire N__19768;
    wire N__19765;
    wire N__19762;
    wire N__19759;
    wire N__19756;
    wire N__19753;
    wire N__19750;
    wire N__19747;
    wire N__19744;
    wire N__19741;
    wire N__19738;
    wire N__19735;
    wire N__19732;
    wire N__19729;
    wire N__19726;
    wire N__19723;
    wire N__19720;
    wire N__19717;
    wire N__19714;
    wire N__19711;
    wire N__19708;
    wire N__19705;
    wire N__19702;
    wire N__19699;
    wire N__19696;
    wire N__19693;
    wire N__19690;
    wire N__19687;
    wire N__19684;
    wire N__19681;
    wire N__19678;
    wire N__19675;
    wire N__19672;
    wire N__19669;
    wire N__19666;
    wire N__19663;
    wire N__19660;
    wire N__19657;
    wire N__19654;
    wire N__19651;
    wire N__19648;
    wire N__19645;
    wire N__19642;
    wire GNDG0;
    wire VCCG0;
    wire \pwm_generator_inst.O_0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_0 ;
    wire bfn_1_7_0_;
    wire \pwm_generator_inst.O_1 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_1 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_0 ;
    wire \pwm_generator_inst.O_2 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_2 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_1 ;
    wire \pwm_generator_inst.O_3 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_3 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_2 ;
    wire \pwm_generator_inst.O_4 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_4 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_3 ;
    wire \pwm_generator_inst.O_5 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_5 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_4 ;
    wire \pwm_generator_inst.O_6 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_6 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_5 ;
    wire \pwm_generator_inst.O_7 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_7 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_6 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_7 ;
    wire \pwm_generator_inst.O_8 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_8 ;
    wire bfn_1_8_0_;
    wire \pwm_generator_inst.O_9 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_9 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_8 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_9 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_10 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_11 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_12 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_13 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_14 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_15 ;
    wire bfn_1_9_0_;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_16 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_17 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_18 ;
    wire \pwm_generator_inst.un3_threshold_acc ;
    wire bfn_1_10_0_;
    wire \pwm_generator_inst.O_12 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_0 ;
    wire \pwm_generator_inst.O_13 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_1 ;
    wire \pwm_generator_inst.O_14 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_2 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_3 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_4 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_5 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_6 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_7 ;
    wire bfn_1_11_0_;
    wire \pwm_generator_inst.un3_threshold_acc_cry_8 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_9 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_10 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_11 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_12 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_13 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_14 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_15 ;
    wire bfn_1_12_0_;
    wire \pwm_generator_inst.un3_threshold_acc_cry_16 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_17 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_18 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_19 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_1_15 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_1_16 ;
    wire N_34_i_i;
    wire \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_ ;
    wire pwm_duty_input_0;
    wire pwm_duty_input_1;
    wire pwm_duty_input_2;
    wire pwm_duty_input_7;
    wire pwm_duty_input_5;
    wire pwm_duty_input_8;
    wire pwm_duty_input_9;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ;
    wire pwm_duty_input_6;
    wire \current_shift_inst.PI_CTRL.N_164 ;
    wire \current_shift_inst.PI_CTRL.N_164_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_120 ;
    wire \current_shift_inst.PI_CTRL.N_167 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_27 ;
    wire \current_shift_inst.PI_CTRL.N_168 ;
    wire \current_shift_inst.PI_CTRL.N_27_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_166 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_12 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_14 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_14_cascade_ ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_15 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_16 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_17 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_ ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_18 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_18_cascade_ ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_10 ;
    wire \pwm_generator_inst.O_10 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_10_cascade_ ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_13 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_0 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_15 ;
    wire \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4 ;
    wire bfn_2_11_0_;
    wire \pwm_generator_inst.un2_threshold_acc_1_16 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_1 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_17 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_2 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_18 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_3 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_19 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_4 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_20 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_5 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_21 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_6 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_22 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_7 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_7 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_23 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_8 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0 ;
    wire bfn_2_12_0_;
    wire \pwm_generator_inst.un2_threshold_acc_1_24 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_9 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_10 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_11 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_12 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_13 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_14 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_25 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_15 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO ;
    wire bfn_2_13_0_;
    wire rgb_drv_RNOZ0;
    wire \current_shift_inst.PI_CTRL.N_162 ;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ;
    wire pwm_duty_input_3;
    wire \pwm_generator_inst.un1_duty_inputlt3 ;
    wire pwm_duty_input_4;
    wire \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_31 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_0 ;
    wire bfn_3_8_0_;
    wire \pwm_generator_inst.un19_threshold_acc_axb_1 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_0 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_2 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_1 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_3 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_2 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_4 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_3 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_5 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_4 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_6 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_5 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_7 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_6 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_7 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_8 ;
    wire bfn_3_9_0_;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_8 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_8 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_4 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5 ;
    wire N_19_1;
    wire \pwm_generator_inst.N_16 ;
    wire \pwm_generator_inst.N_17 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_1 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_6 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_7 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_5 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_2 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_3 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_9 ;
    wire bfn_5_8_0_;
    wire \pwm_generator_inst.counter_cry_0 ;
    wire \pwm_generator_inst.counter_cry_1 ;
    wire \pwm_generator_inst.counter_cry_2 ;
    wire \pwm_generator_inst.counter_cry_3 ;
    wire \pwm_generator_inst.counter_cry_4 ;
    wire \pwm_generator_inst.counter_cry_5 ;
    wire \pwm_generator_inst.counter_cry_6 ;
    wire \pwm_generator_inst.counter_cry_7 ;
    wire bfn_5_9_0_;
    wire \pwm_generator_inst.counter_cry_8 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_0 ;
    wire \pwm_generator_inst.un1_counterlto9_2_cascade_ ;
    wire \pwm_generator_inst.un1_counter_0 ;
    wire \pwm_generator_inst.un1_counterlto2_0_cascade_ ;
    wire \pwm_generator_inst.un1_counterlt9 ;
    wire \pwm_generator_inst.thresholdZ0Z_0 ;
    wire \pwm_generator_inst.counterZ0Z_0 ;
    wire \pwm_generator_inst.counter_i_0 ;
    wire bfn_5_11_0_;
    wire \pwm_generator_inst.thresholdZ0Z_1 ;
    wire \pwm_generator_inst.counterZ0Z_1 ;
    wire \pwm_generator_inst.counter_i_1 ;
    wire \pwm_generator_inst.un14_counter_cry_0 ;
    wire \pwm_generator_inst.thresholdZ0Z_2 ;
    wire \pwm_generator_inst.counterZ0Z_2 ;
    wire \pwm_generator_inst.counter_i_2 ;
    wire \pwm_generator_inst.un14_counter_cry_1 ;
    wire \pwm_generator_inst.thresholdZ0Z_3 ;
    wire \pwm_generator_inst.counterZ0Z_3 ;
    wire \pwm_generator_inst.counter_i_3 ;
    wire \pwm_generator_inst.un14_counter_cry_2 ;
    wire \pwm_generator_inst.thresholdZ0Z_4 ;
    wire \pwm_generator_inst.counterZ0Z_4 ;
    wire \pwm_generator_inst.counter_i_4 ;
    wire \pwm_generator_inst.un14_counter_cry_3 ;
    wire \pwm_generator_inst.thresholdZ0Z_5 ;
    wire \pwm_generator_inst.counterZ0Z_5 ;
    wire \pwm_generator_inst.counter_i_5 ;
    wire \pwm_generator_inst.un14_counter_cry_4 ;
    wire \pwm_generator_inst.counterZ0Z_6 ;
    wire \pwm_generator_inst.thresholdZ0Z_6 ;
    wire \pwm_generator_inst.counter_i_6 ;
    wire \pwm_generator_inst.un14_counter_cry_5 ;
    wire \pwm_generator_inst.thresholdZ0Z_7 ;
    wire \pwm_generator_inst.counterZ0Z_7 ;
    wire \pwm_generator_inst.counter_i_7 ;
    wire \pwm_generator_inst.un14_counter_cry_6 ;
    wire \pwm_generator_inst.un14_counter_cry_7 ;
    wire \pwm_generator_inst.thresholdZ0Z_8 ;
    wire \pwm_generator_inst.counterZ0Z_8 ;
    wire \pwm_generator_inst.counter_i_8 ;
    wire bfn_5_12_0_;
    wire \pwm_generator_inst.thresholdZ0Z_9 ;
    wire \pwm_generator_inst.counterZ0Z_9 ;
    wire \pwm_generator_inst.counter_i_9 ;
    wire \pwm_generator_inst.un14_counter_cry_8 ;
    wire \pwm_generator_inst.un14_counter_cry_9 ;
    wire pwm_output_c;
    wire start_stop_c;
    wire \phase_controller_inst1.start_timer_tr_0_sqmuxa ;
    wire \phase_controller_inst1.state_RNI7NN7Z0Z_0 ;
    wire il_max_comp1_D2;
    wire il_min_comp2_c;
    wire il_min_comp2_D1;
    wire il_max_comp2_c;
    wire il_max_comp2_D1;
    wire \delay_measurement_inst.delay_hc_timer.N_302_i ;
    wire \phase_controller_inst2.start_timer_tr_0_sqmuxa ;
    wire \phase_controller_inst2.state_RNI9M3OZ0Z_0 ;
    wire \phase_controller_inst2.state_RNI9M3OZ0Z_0_cascade_ ;
    wire state_ns_i_a3_1;
    wire il_min_comp2_D2;
    wire \phase_controller_inst2.tr_time_passed ;
    wire \phase_controller_inst2.stateZ0Z_0 ;
    wire bfn_7_15_0_;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_4 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_7 ;
    wire bfn_7_16_0_;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_15 ;
    wire bfn_7_17_0_;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_inst1.stateZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa ;
    wire il_min_comp1_D2;
    wire \phase_controller_inst1.tr_time_passed ;
    wire \phase_controller_inst1.stateZ0Z_0 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0 ;
    wire \phase_controller_inst2.stateZ0Z_1 ;
    wire s4_phy_c;
    wire il_max_comp1_c;
    wire il_max_comp1_D1;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_53 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_118 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_7 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_3 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_6 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_5 ;
    wire \phase_controller_inst2.stoper_tr.time_passed_1_sqmuxa ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2 ;
    wire \phase_controller_inst2.stoper_tr.time_passed11_cascade_ ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNIF9HJZ0 ;
    wire \phase_controller_inst2.stoper_tr.time_passed11 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_axb_0 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_13 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_14 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_15 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_17 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_18 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_19 ;
    wire \phase_controller_inst1.start_timer_hc_0_sqmuxa ;
    wire \phase_controller_inst1.start_timer_hc_RNOZ0Z_0 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_1 ;
    wire bfn_8_17_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_9 ;
    wire bfn_8_18_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_17 ;
    wire bfn_8_19_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_19 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ;
    wire bfn_8_20_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7 ;
    wire bfn_8_21_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17 ;
    wire bfn_8_22_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19 ;
    wire \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa ;
    wire \phase_controller_inst1.hc_time_passed ;
    wire clk_12mhz;
    wire GB_BUFFER_clk_12mhz_THRU_CO;
    wire il_min_comp1_c;
    wire il_min_comp1_D1;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ;
    wire bfn_9_8_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto3 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto4 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ;
    wire bfn_9_9_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ;
    wire bfn_9_10_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ;
    wire bfn_9_11_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ;
    wire \current_shift_inst.PI_CTRL.un8_enablelto31 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_1 ;
    wire bfn_9_13_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_9 ;
    wire bfn_9_14_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_16 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_17 ;
    wire bfn_9_15_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_18 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_19 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ;
    wire \phase_controller_inst2.start_timer_hc_0_sqmuxa_cascade_ ;
    wire phase_controller_inst1_state_4;
    wire il_max_comp2_D2;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ;
    wire \phase_controller_inst1.start_timer_trZ0 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_inst1.stoper_tr.time_passed11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_0 ;
    wire bfn_9_22_0_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_1 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_8 ;
    wire bfn_9_23_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_9 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_16 ;
    wire bfn_9_24_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_17 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_inst2.stateZ0Z_3 ;
    wire s3_phy_c;
    wire \phase_controller_inst1.stateZ0Z_1 ;
    wire s2_phy_c;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_0 ;
    wire \delay_measurement_inst.hc_stateZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_26 ;
    wire \delay_measurement_inst.start_timer_hcZ0 ;
    wire \delay_measurement_inst.stop_timer_hcZ0 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3Z0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4Z0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.N_248 ;
    wire \phase_controller_inst1.stoper_tr.N_248_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.N_55 ;
    wire bfn_10_17_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_1 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_8 ;
    wire bfn_10_18_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_9 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_16 ;
    wire bfn_10_19_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_17 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_18 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_19 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_axb_0 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ1Z_6 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_0 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ;
    wire bfn_10_24_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9 ;
    wire bfn_10_25_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17 ;
    wire bfn_10_26_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19 ;
    wire delay_hc_input_c;
    wire delay_hc_d1;
    wire delay_hc_d2;
    wire \delay_measurement_inst.prev_hc_sigZ0 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_10 ;
    wire measured_delay_tr_7;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_21 ;
    wire measured_delay_tr_8;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_25 ;
    wire measured_delay_tr_5;
    wire measured_delay_tr_4;
    wire measured_delay_tr_9;
    wire measured_delay_tr_3;
    wire measured_delay_tr_2;
    wire measured_delay_tr_6;
    wire measured_delay_tr_1;
    wire measured_delay_tr_14;
    wire measured_delay_tr_12;
    wire measured_delay_tr_11;
    wire measured_delay_tr_13;
    wire measured_delay_tr_10;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6 ;
    wire measured_delay_tr_16;
    wire \phase_controller_inst2.stoper_hc.time_passed_1_sqmuxa ;
    wire \phase_controller_inst2.stateZ0Z_2 ;
    wire \phase_controller_inst2.hc_time_passed ;
    wire \phase_controller_inst2.start_timer_hc_RNO_0_0 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ;
    wire bfn_11_18_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_2 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_3 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_4 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_5 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_7 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_8 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_7 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_9 ;
    wire bfn_11_19_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_10 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_11 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_12 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_13 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_14 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_15 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_16 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_17 ;
    wire bfn_11_20_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_18 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_19 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ1Z_6 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.time_passed11 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_72 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_18_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_7 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_15 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ;
    wire \delay_measurement_inst.N_267 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3 ;
    wire \delay_measurement_inst.delay_tr_timer.N_287_4_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_290 ;
    wire \delay_measurement_inst.N_59 ;
    wire \delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10 ;
    wire \delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_5 ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_0_cascade_ ;
    wire \delay_measurement_inst.un3_elapsed_time_tr_0_i ;
    wire \delay_measurement_inst.un3_elapsed_time_tr_0_i_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_5 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6Z0Z_7 ;
    wire \delay_measurement_inst.N_299 ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_287_4 ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6 ;
    wire \delay_measurement_inst.N_265 ;
    wire \delay_measurement_inst.N_265_cascade_ ;
    wire \delay_measurement_inst.N_270 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19 ;
    wire measured_delay_tr_17;
    wire measured_delay_tr_18;
    wire \delay_measurement_inst.N_325 ;
    wire measured_delay_tr_19;
    wire \delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_fast_31 ;
    wire \current_shift_inst.un4_control_input1_1 ;
    wire \current_shift_inst.un4_control_input1_1_cascade_ ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0 ;
    wire \phase_controller_inst2.start_timer_hcZ0 ;
    wire \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.time_passed11 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIUO2PZ0 ;
    wire \phase_controller_inst2.start_timer_trZ0 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0 ;
    wire \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_11_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un2_startlt31 ;
    wire \delay_measurement_inst.delay_hc_timer.runningZ0 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto5Z0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlt9_0_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un1_startlt15 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto13Z0Z_1 ;
    wire \phase_controller_inst1.start_timer_hcZ0 ;
    wire \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto8Z0Z_0 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlt31_0 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ;
    wire measured_delay_hc_10;
    wire measured_delay_hc_31;
    wire measured_delay_hc_3;
    wire measured_delay_hc_12;
    wire measured_delay_hc_18;
    wire measured_delay_hc_17;
    wire measured_delay_hc_5;
    wire measured_delay_hc_11;
    wire measured_delay_hc_9;
    wire measured_delay_hc_14;
    wire measured_delay_hc_6;
    wire measured_delay_hc_13;
    wire measured_delay_hc_24;
    wire measured_delay_hc_25;
    wire measured_delay_hc_26;
    wire measured_delay_hc_23;
    wire state_3;
    wire s1_phy_c;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_11 ;
    wire \current_shift_inst.PI_CTRL.un1_enablelt3_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_71 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axb_0 ;
    wire bfn_13_10_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_0 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_7 ;
    wire bfn_13_11_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_8 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_11 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_12 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_13 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_14 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_15 ;
    wire bfn_13_12_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_16 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_17 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_18 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_19 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_20 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_21 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_22 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_23 ;
    wire bfn_13_13_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_24 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_25 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ;
    wire \current_shift_inst.un38_control_input_cry_0_s0_sf ;
    wire bfn_13_17_0_;
    wire \current_shift_inst.un38_control_input_cry_0_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ;
    wire \current_shift_inst.un38_control_input_cry_1_s0 ;
    wire \current_shift_inst.un38_control_input_cry_2_s0 ;
    wire \current_shift_inst.un38_control_input_cry_3_s0 ;
    wire \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_4_s0 ;
    wire \current_shift_inst.un38_control_input_cry_5_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8 ;
    wire \current_shift_inst.un38_control_input_cry_6_s0 ;
    wire \current_shift_inst.un38_control_input_cry_7_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9 ;
    wire \current_shift_inst.un38_control_input_0_s0_8 ;
    wire bfn_13_18_0_;
    wire \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10 ;
    wire \current_shift_inst.un38_control_input_0_s0_9 ;
    wire \current_shift_inst.un38_control_input_cry_8_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11 ;
    wire \current_shift_inst.un38_control_input_0_s0_10 ;
    wire \current_shift_inst.un38_control_input_cry_9_s0 ;
    wire \current_shift_inst.un38_control_input_cry_10_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_12 ;
    wire \current_shift_inst.un38_control_input_cry_11_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14 ;
    wire \current_shift_inst.un38_control_input_cry_12_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15 ;
    wire \current_shift_inst.un38_control_input_0_s0_14 ;
    wire \current_shift_inst.un38_control_input_cry_13_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16 ;
    wire \current_shift_inst.un38_control_input_0_s0_15 ;
    wire \current_shift_inst.un38_control_input_cry_14_s0 ;
    wire \current_shift_inst.un38_control_input_cry_15_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_16 ;
    wire bfn_13_19_0_;
    wire \current_shift_inst.un38_control_input_0_s0_17 ;
    wire \current_shift_inst.un38_control_input_cry_16_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_18 ;
    wire \current_shift_inst.un38_control_input_cry_17_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_19 ;
    wire \current_shift_inst.un38_control_input_cry_18_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_21 ;
    wire \current_shift_inst.un38_control_input_cry_20_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ;
    wire \current_shift_inst.un38_control_input_cry_21_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_23 ;
    wire \current_shift_inst.un38_control_input_cry_22_s0 ;
    wire \current_shift_inst.un38_control_input_cry_23_s0 ;
    wire bfn_13_20_0_;
    wire \current_shift_inst.un38_control_input_cry_24_s0 ;
    wire \current_shift_inst.un38_control_input_cry_25_s0 ;
    wire \current_shift_inst.un38_control_input_cry_26_s0 ;
    wire \current_shift_inst.un38_control_input_cry_27_s0 ;
    wire \current_shift_inst.un38_control_input_cry_28_s0 ;
    wire \current_shift_inst.un38_control_input_cry_29_s0 ;
    wire \current_shift_inst.un38_control_input_cry_30_s0 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlt3 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_6 ;
    wire measured_delay_hc_22;
    wire measured_delay_hc_7;
    wire measured_delay_hc_0;
    wire measured_delay_hc_20;
    wire measured_delay_hc_16;
    wire measured_delay_hc_1;
    wire measured_delay_hc_8;
    wire measured_delay_hc_21;
    wire measured_delay_hc_15;
    wire measured_delay_hc_4;
    wire measured_delay_hc_2;
    wire measured_delay_hc_19;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto5_2_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclt31_0_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_7 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt13_0 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt19 ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt8 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt13_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt19_0_cascade_ ;
    wire \current_shift_inst.start_timer_sZ0Z1 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_2 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_3 ;
    wire \current_shift_inst.stop_timer_sZ0Z1 ;
    wire \current_shift_inst.timer_s1.N_180_i ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_0 ;
    wire bfn_14_7_0_;
    wire \current_shift_inst.PI_CTRL.prop_term_1_1 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_1 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_2 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_2 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_3 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_3 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_4 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_5 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_6 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_7 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_8 ;
    wire bfn_14_8_0_;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_9 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_10 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_11 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ;
    wire bfn_14_9_0_;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23 ;
    wire bfn_14_10_0_;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_31 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15 ;
    wire measured_delay_tr_15;
    wire \phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23 ;
    wire \current_shift_inst.control_inputZ0Z_0 ;
    wire bfn_14_15_0_;
    wire \current_shift_inst.control_inputZ0Z_1 ;
    wire \current_shift_inst.control_input_1_cry_0 ;
    wire \current_shift_inst.control_input_1_axb_2 ;
    wire \current_shift_inst.control_inputZ0Z_2 ;
    wire \current_shift_inst.control_input_1_cry_1 ;
    wire \current_shift_inst.control_input_1_axb_3 ;
    wire \current_shift_inst.control_inputZ0Z_3 ;
    wire \current_shift_inst.control_input_1_cry_2 ;
    wire \current_shift_inst.control_input_1_axb_4 ;
    wire \current_shift_inst.control_inputZ0Z_4 ;
    wire \current_shift_inst.control_input_1_cry_3 ;
    wire \current_shift_inst.control_inputZ0Z_5 ;
    wire \current_shift_inst.control_input_1_cry_4 ;
    wire \current_shift_inst.control_input_1_axb_6 ;
    wire \current_shift_inst.control_inputZ0Z_6 ;
    wire \current_shift_inst.control_input_1_cry_5 ;
    wire \current_shift_inst.control_inputZ0Z_7 ;
    wire \current_shift_inst.control_input_1_cry_6 ;
    wire \current_shift_inst.control_input_1_cry_7 ;
    wire \current_shift_inst.control_input_1_axb_8 ;
    wire \current_shift_inst.control_inputZ0Z_8 ;
    wire bfn_14_16_0_;
    wire \current_shift_inst.control_input_1_axb_9 ;
    wire \current_shift_inst.control_inputZ0Z_9 ;
    wire \current_shift_inst.control_input_1_cry_8 ;
    wire \current_shift_inst.control_input_1_axb_10 ;
    wire \current_shift_inst.control_inputZ0Z_10 ;
    wire \current_shift_inst.control_input_1_cry_9 ;
    wire \current_shift_inst.control_input_1_axb_11 ;
    wire \current_shift_inst.control_inputZ0Z_11 ;
    wire \current_shift_inst.control_input_1_cry_10 ;
    wire \current_shift_inst.control_input_1_axb_12 ;
    wire \current_shift_inst.control_inputZ0Z_12 ;
    wire \current_shift_inst.control_input_1_cry_11 ;
    wire \current_shift_inst.control_input_1_axb_13 ;
    wire \current_shift_inst.control_inputZ0Z_13 ;
    wire \current_shift_inst.control_input_1_cry_12 ;
    wire \current_shift_inst.control_input_1_axb_14 ;
    wire \current_shift_inst.control_inputZ0Z_14 ;
    wire \current_shift_inst.control_input_1_cry_13 ;
    wire \current_shift_inst.control_input_1_axb_15 ;
    wire \current_shift_inst.control_inputZ0Z_15 ;
    wire \current_shift_inst.control_input_1_cry_14 ;
    wire \current_shift_inst.control_input_1_cry_15 ;
    wire \current_shift_inst.control_inputZ0Z_16 ;
    wire bfn_14_17_0_;
    wire \current_shift_inst.control_input_1_axb_17 ;
    wire \current_shift_inst.control_inputZ0Z_17 ;
    wire \current_shift_inst.control_input_1_cry_16 ;
    wire \current_shift_inst.control_inputZ0Z_18 ;
    wire \current_shift_inst.control_input_1_cry_17 ;
    wire \current_shift_inst.control_inputZ0Z_19 ;
    wire \current_shift_inst.control_input_1_cry_18 ;
    wire \current_shift_inst.control_inputZ0Z_20 ;
    wire \current_shift_inst.control_input_1_cry_19 ;
    wire \current_shift_inst.control_inputZ0Z_21 ;
    wire \current_shift_inst.control_input_1_cry_20 ;
    wire \current_shift_inst.control_inputZ0Z_22 ;
    wire \current_shift_inst.control_input_1_cry_21 ;
    wire \current_shift_inst.control_inputZ0Z_23 ;
    wire \current_shift_inst.control_input_1_cry_22 ;
    wire \current_shift_inst.control_input_1_cry_23 ;
    wire \current_shift_inst.control_inputZ0Z_24 ;
    wire bfn_14_18_0_;
    wire \current_shift_inst.control_input_1_axb_25 ;
    wire \current_shift_inst.control_input_1_cry_24 ;
    wire \current_shift_inst.control_inputZ0Z_25 ;
    wire \current_shift_inst.un38_control_input_0_s0_28 ;
    wire \current_shift_inst.control_input_1_axb_22 ;
    wire \current_shift_inst.N_1355_i ;
    wire \current_shift_inst.un38_control_input_0_s0_6 ;
    wire \current_shift_inst.control_input_1_axb_0 ;
    wire \current_shift_inst.un38_control_input_0_s0_22 ;
    wire \current_shift_inst.control_input_1_axb_16 ;
    wire \current_shift_inst.un38_control_input_0_s0_29 ;
    wire \current_shift_inst.control_input_1_axb_23 ;
    wire \current_shift_inst.un38_control_input_0_s0_7 ;
    wire \current_shift_inst.control_input_1_axb_1 ;
    wire \current_shift_inst.un38_control_input_0_s0_27 ;
    wire \current_shift_inst.control_input_1_axb_21 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19 ;
    wire \current_shift_inst.un38_control_input_0_s0_24 ;
    wire \current_shift_inst.control_input_1_axb_18 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ;
    wire \current_shift_inst.un38_control_input_0_s0_26 ;
    wire \current_shift_inst.control_input_1_axb_20 ;
    wire \current_shift_inst.un38_control_input_0_s0_25 ;
    wire \current_shift_inst.control_input_1_axb_19 ;
    wire \current_shift_inst.un38_control_input_0_s0_30 ;
    wire \current_shift_inst.control_input_1_axb_24 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ;
    wire bfn_14_21_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_7 ;
    wire bfn_14_22_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_15 ;
    wire bfn_14_23_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_23 ;
    wire bfn_14_24_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.running_i ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.N_303_i ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_10 ;
    wire \delay_measurement_inst.elapsed_time_hc_3 ;
    wire bfn_14_26_0_;
    wire \delay_measurement_inst.elapsed_time_hc_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.elapsed_time_hc_5 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_hc_reg3lto6 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.elapsed_time_hc_7 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.elapsed_time_hc_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_hc_reg3lto9 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.elapsed_time_hc_10 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ;
    wire \delay_measurement_inst.elapsed_time_hc_11 ;
    wire bfn_14_27_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.elapsed_time_hc_12 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.elapsed_time_hc_13 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_hc_reg3lto14 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_hc_reg3lto15 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ;
    wire bfn_14_28_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ;
    wire bfn_14_29_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ;
    wire delay_tr_input_c;
    wire delay_tr_d1;
    wire red_c_i;
    wire \current_shift_inst.PI_CTRL.prop_term_1_13 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_13 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_6 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_6 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_5 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_5 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_4 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_4 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_8 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_8 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_7 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_7 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_9 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_9 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_10 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_10 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_12 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_12 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_11 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_11 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_22 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_22 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_19 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_19 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_15 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_15 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_16 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_16 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_23 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_23 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_20 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_20 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO ;
    wire \delay_measurement_inst.elapsed_time_tr_3 ;
    wire bfn_15_11_0_;
    wire \delay_measurement_inst.elapsed_time_tr_4 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.elapsed_time_tr_5 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_tr_reg3lto6 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.elapsed_time_tr_7 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.elapsed_time_tr_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_tr_reg3lto9 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.elapsed_time_tr_10 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.elapsed_time_tr_11 ;
    wire bfn_15_12_0_;
    wire \delay_measurement_inst.elapsed_time_tr_12 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.elapsed_time_tr_13 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_tr_reg3lto14 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_tr_reg3lto15 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.elapsed_time_tr_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.elapsed_time_tr_17 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.elapsed_time_tr_18 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.elapsed_time_tr_19 ;
    wire bfn_15_13_0_;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ;
    wire bfn_15_14_0_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.elapsed_time_tr_31 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_31 ;
    wire bfn_15_15_0_;
    wire \current_shift_inst.un10_control_input_cry_0 ;
    wire \current_shift_inst.un10_control_input_cry_1 ;
    wire \current_shift_inst.un10_control_input_cry_2 ;
    wire \current_shift_inst.un10_control_input_cry_3 ;
    wire \current_shift_inst.un10_control_input_cry_4 ;
    wire \current_shift_inst.un10_control_input_cry_5 ;
    wire \current_shift_inst.un10_control_input_cry_6 ;
    wire \current_shift_inst.un10_control_input_cry_7 ;
    wire bfn_15_16_0_;
    wire \current_shift_inst.un10_control_input_cry_8 ;
    wire \current_shift_inst.un10_control_input_cry_9 ;
    wire \current_shift_inst.un10_control_input_cry_10 ;
    wire \current_shift_inst.un10_control_input_cry_11 ;
    wire \current_shift_inst.un10_control_input_cry_12 ;
    wire \current_shift_inst.un10_control_input_cry_13 ;
    wire \current_shift_inst.un10_control_input_cry_14 ;
    wire \current_shift_inst.un10_control_input_cry_15 ;
    wire bfn_15_17_0_;
    wire \current_shift_inst.un10_control_input_cry_16 ;
    wire \current_shift_inst.un10_control_input_cry_17 ;
    wire \current_shift_inst.un10_control_input_cry_18 ;
    wire \current_shift_inst.un10_control_input_cry_19 ;
    wire \current_shift_inst.un10_control_input_cry_20 ;
    wire \current_shift_inst.un10_control_input_cry_21 ;
    wire \current_shift_inst.un10_control_input_cry_22 ;
    wire \current_shift_inst.un10_control_input_cry_23 ;
    wire bfn_15_18_0_;
    wire \current_shift_inst.un10_control_input_cry_24 ;
    wire \current_shift_inst.un10_control_input_cry_25 ;
    wire \current_shift_inst.un10_control_input_cry_26 ;
    wire \current_shift_inst.un10_control_input_cry_27 ;
    wire \current_shift_inst.un10_control_input_cry_28 ;
    wire CONSTANT_ONE_NET;
    wire \current_shift_inst.un10_control_input_cry_29 ;
    wire \current_shift_inst.un10_control_input_cry_30 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ;
    wire \current_shift_inst.un38_control_input_5_0 ;
    wire bfn_15_19_0_;
    wire \current_shift_inst.un38_control_input_cry_0_s1 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1 ;
    wire \current_shift_inst.un38_control_input_cry_3_s1 ;
    wire \current_shift_inst.un38_control_input_cry_4_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_6 ;
    wire \current_shift_inst.un38_control_input_cry_5_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_7 ;
    wire \current_shift_inst.un38_control_input_cry_6_s1 ;
    wire \current_shift_inst.un38_control_input_cry_7_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_8 ;
    wire bfn_15_20_0_;
    wire \current_shift_inst.un38_control_input_0_s1_9 ;
    wire \current_shift_inst.un38_control_input_cry_8_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_10 ;
    wire \current_shift_inst.un38_control_input_cry_9_s1 ;
    wire \current_shift_inst.un38_control_input_cry_10_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_12 ;
    wire \current_shift_inst.un38_control_input_cry_11_s1 ;
    wire \current_shift_inst.un38_control_input_cry_12_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_14 ;
    wire \current_shift_inst.un38_control_input_cry_13_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_15 ;
    wire \current_shift_inst.un38_control_input_cry_14_s1 ;
    wire \current_shift_inst.un38_control_input_cry_15_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_16 ;
    wire bfn_15_21_0_;
    wire \current_shift_inst.un38_control_input_0_s1_17 ;
    wire \current_shift_inst.un38_control_input_cry_16_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_18 ;
    wire \current_shift_inst.un38_control_input_cry_17_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_19 ;
    wire \current_shift_inst.un38_control_input_cry_18_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_21 ;
    wire \current_shift_inst.un38_control_input_cry_20_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_22 ;
    wire \current_shift_inst.un38_control_input_cry_21_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_23 ;
    wire \current_shift_inst.un38_control_input_cry_22_s1 ;
    wire \current_shift_inst.un38_control_input_cry_23_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_24 ;
    wire bfn_15_22_0_;
    wire \current_shift_inst.un38_control_input_0_s1_25 ;
    wire \current_shift_inst.un38_control_input_cry_24_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_26 ;
    wire \current_shift_inst.un38_control_input_cry_25_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_27 ;
    wire \current_shift_inst.un38_control_input_cry_26_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_28 ;
    wire \current_shift_inst.un38_control_input_cry_27_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_29 ;
    wire \current_shift_inst.un38_control_input_cry_28_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_30 ;
    wire \current_shift_inst.un38_control_input_cry_29_s1 ;
    wire \current_shift_inst.un38_control_input_cry_30_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_31 ;
    wire \delay_measurement_inst.elapsed_time_hc_18 ;
    wire \delay_measurement_inst.elapsed_time_hc_17 ;
    wire \delay_measurement_inst.elapsed_time_hc_16 ;
    wire \delay_measurement_inst.elapsed_time_hc_19 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ;
    wire \delay_measurement_inst.elapsed_time_hc_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.elapsed_time_hc_2 ;
    wire \delay_measurement_inst.delay_hc_timer.N_302_i_g ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_3_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto30Z0Z_1 ;
    wire \delay_measurement_inst.delay_tr_timer.N_304_i ;
    wire \delay_measurement_inst.tr_stateZ0Z_0 ;
    wire delay_tr_d2;
    wire \delay_measurement_inst.prev_tr_sigZ0 ;
    wire \delay_measurement_inst.start_timer_trZ0 ;
    wire \delay_measurement_inst.stop_timer_trZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.runningZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_i_26 ;
    wire bfn_16_8_0_;
    wire \current_shift_inst.PI_CTRL.error_control_RNI4Q3UZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_0 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.error_control_RNI8V4UZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_0 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIC46UZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIG97UZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_3 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIKE8UZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIOJ9UZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_5 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIA1B41Z0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_5 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIL0S01Z0Z_11 ;
    wire bfn_16_9_0_;
    wire \current_shift_inst.PI_CTRL.error_control_RNIP5T01Z0Z_12 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNITAU01Z0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_8 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNICE9PZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_11 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIGJAPZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_13 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_14 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIS2EPZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ;
    wire bfn_16_10_0_;
    wire \current_shift_inst.PI_CTRL.error_control_RNIENGPZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_17 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_16 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIDGBQZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_17 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIHLCQZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_18 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_21 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_20 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIKD7JZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_21 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_22 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIMG8JZ0 ;
    wire bfn_16_11_0_;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIOJ9JZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_23 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNIQMAJZ0 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_24 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNISPBJZ0 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_25 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNILB5KZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_26 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_29 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_30 ;
    wire bfn_16_12_0_;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_20 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_i_0_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_19 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_24 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_24 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNICIEQZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_19 ;
    wire \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ;
    wire \current_shift_inst.un38_control_input_5_1 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_2 ;
    wire \current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10 ;
    wire \current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13 ;
    wire \current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ;
    wire \current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14 ;
    wire \current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11 ;
    wire \current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNID8O11_12 ;
    wire \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJO221_20 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI25021_19 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ;
    wire \current_shift_inst.un4_control_input_0_31 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_26 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_28 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISST11_17 ;
    wire measured_delay_hc_29;
    wire measured_delay_hc_30;
    wire measured_delay_hc_27;
    wire \delay_measurement_inst.un1_elapsed_time_hc ;
    wire \delay_measurement_inst.delay_hc_reg3 ;
    wire measured_delay_hc_28;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_18 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_18 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIOTCPZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_25 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIGNFQZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_25 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_21 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_21 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNI9BAQZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_12 ;
    wire bfn_17_11_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ;
    wire bfn_17_12_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ;
    wire bfn_17_13_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ;
    wire bfn_17_14_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.running_i ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_tr_timer.N_305_i ;
    wire \current_shift_inst.un4_control_input_1_axb_1 ;
    wire \current_shift_inst.un4_control_input1_2 ;
    wire bfn_17_15_0_;
    wire \current_shift_inst.un4_control_input_1_cry_1 ;
    wire \current_shift_inst.un4_control_input1_4 ;
    wire \current_shift_inst.un4_control_input_1_cry_2 ;
    wire \current_shift_inst.un4_control_input_1_cry_3 ;
    wire \current_shift_inst.un4_control_input1_6 ;
    wire \current_shift_inst.un4_control_input_1_cry_4 ;
    wire \current_shift_inst.un4_control_input_1_cry_5 ;
    wire \current_shift_inst.un4_control_input_1_cry_6 ;
    wire \current_shift_inst.un4_control_input1_9 ;
    wire \current_shift_inst.un4_control_input_1_cry_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_8 ;
    wire \current_shift_inst.un4_control_input1_10 ;
    wire bfn_17_16_0_;
    wire \current_shift_inst.un4_control_input1_11 ;
    wire \current_shift_inst.un4_control_input_1_cry_9 ;
    wire \current_shift_inst.un4_control_input_1_cry_10 ;
    wire \current_shift_inst.un4_control_input1_13 ;
    wire \current_shift_inst.un4_control_input_1_cry_11 ;
    wire \current_shift_inst.un4_control_input1_14 ;
    wire \current_shift_inst.un4_control_input_1_cry_12 ;
    wire \current_shift_inst.un4_control_input1_15 ;
    wire \current_shift_inst.un4_control_input_1_cry_13 ;
    wire \current_shift_inst.un4_control_input1_16 ;
    wire \current_shift_inst.un4_control_input_1_cry_14 ;
    wire \current_shift_inst.un4_control_input_1_cry_15 ;
    wire \current_shift_inst.un4_control_input_1_cry_16 ;
    wire bfn_17_17_0_;
    wire \current_shift_inst.un4_control_input_1_cry_17 ;
    wire \current_shift_inst.un4_control_input1_20 ;
    wire \current_shift_inst.un4_control_input_1_cry_18 ;
    wire \current_shift_inst.un4_control_input1_21 ;
    wire \current_shift_inst.un4_control_input_1_cry_19 ;
    wire \current_shift_inst.un4_control_input1_22 ;
    wire \current_shift_inst.un4_control_input_1_cry_20 ;
    wire \current_shift_inst.un4_control_input1_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_21 ;
    wire \current_shift_inst.un4_control_input_1_cry_22 ;
    wire \current_shift_inst.un4_control_input1_25 ;
    wire \current_shift_inst.un4_control_input_1_cry_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_24 ;
    wire bfn_17_18_0_;
    wire \current_shift_inst.un4_control_input1_27 ;
    wire \current_shift_inst.un4_control_input_1_cry_25 ;
    wire \current_shift_inst.un4_control_input_1_cry_26 ;
    wire \current_shift_inst.un4_control_input1_29 ;
    wire \current_shift_inst.un4_control_input_1_cry_27 ;
    wire \current_shift_inst.un4_control_input1_30 ;
    wire \current_shift_inst.un4_control_input_1_cry_28 ;
    wire \current_shift_inst.un4_control_input1_31 ;
    wire \current_shift_inst.un4_control_input1_31_THRU_CO ;
    wire \current_shift_inst.un4_control_input1_31_THRU_CO_cascade_ ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_axb_18 ;
    wire \current_shift_inst.un4_control_input1_24 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ;
    wire \current_shift_inst.un4_control_input_1_axb_21 ;
    wire \current_shift_inst.un4_control_input_1_axb_22 ;
    wire \current_shift_inst.un4_control_input_1_axb_17 ;
    wire \current_shift_inst.un4_control_input_1_axb_25 ;
    wire \current_shift_inst.un4_control_input_1_axb_20 ;
    wire \current_shift_inst.un4_control_input1_18 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18 ;
    wire \current_shift_inst.un4_control_input_1_axb_19 ;
    wire \current_shift_inst.un4_control_input_1_axb_24 ;
    wire \current_shift_inst.un4_control_input1_28 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ;
    wire \current_shift_inst.un4_control_input_1_axb_26 ;
    wire \current_shift_inst.un4_control_input_1_axb_28 ;
    wire \current_shift_inst.un4_control_input1_26 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ;
    wire \current_shift_inst.un4_control_input_1_axb_29 ;
    wire \current_shift_inst.timer_s1.runningZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_17 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_17 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIKOBPZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_10 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_7 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_13 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_26 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_14 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_14 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNI898PZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ;
    wire \current_shift_inst.PI_CTRL.N_74 ;
    wire \current_shift_inst.PI_CTRL.N_75 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_31 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_26 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_24 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_28 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_23 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.elapsed_time_tr_2 ;
    wire \current_shift_inst.un4_control_input_1_axb_27 ;
    wire \current_shift_inst.un4_control_input1_5 ;
    wire \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7 ;
    wire \current_shift_inst.un4_control_input1_17 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17 ;
    wire \current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_axb_31_s0 ;
    wire \current_shift_inst.un4_control_input1_19 ;
    wire \current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ;
    wire \current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_1 ;
    wire \current_shift_inst.un4_control_input_1_axb_8 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31_rep1 ;
    wire \current_shift_inst.un4_control_input1_3 ;
    wire \current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_12 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12 ;
    wire \current_shift_inst.un4_control_input1_7 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7 ;
    wire \current_shift_inst.un38_control_input_0_s0_11 ;
    wire \current_shift_inst.un38_control_input_0_s1_11 ;
    wire \current_shift_inst.control_input_1_axb_5 ;
    wire \current_shift_inst.un38_control_input_0_s0_13 ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ;
    wire \current_shift_inst.un38_control_input_0_s1_13 ;
    wire \current_shift_inst.control_input_1_axb_7 ;
    wire \current_shift_inst.un4_control_input_1_axb_3 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31 ;
    wire \current_shift_inst.un38_control_input_5_2 ;
    wire \current_shift_inst.un4_control_input1_8 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8 ;
    wire \current_shift_inst.un4_control_input_1_axb_15 ;
    wire \current_shift_inst.un4_control_input_1_axb_7 ;
    wire \current_shift_inst.un4_control_input_1_axb_2 ;
    wire \current_shift_inst.un4_control_input_1_axb_6 ;
    wire \current_shift_inst.un4_control_input_1_axb_4 ;
    wire \current_shift_inst.un4_control_input_1_axb_5 ;
    wire \current_shift_inst.un4_control_input_1_axb_11 ;
    wire \current_shift_inst.un4_control_input_1_axb_13 ;
    wire \current_shift_inst.un4_control_input_1_axb_9 ;
    wire \current_shift_inst.un4_control_input_1_axb_14 ;
    wire \current_shift_inst.un4_control_input_1_axb_16 ;
    wire \current_shift_inst.un4_control_input_1_axb_23 ;
    wire \current_shift_inst.un4_control_input_1_axb_10 ;
    wire \current_shift_inst.un4_control_input_1_axb_12 ;
    wire \current_shift_inst.elapsed_time_ns_s1_3 ;
    wire bfn_18_18_0_;
    wire \current_shift_inst.elapsed_time_ns_s1_4 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ;
    wire \current_shift_inst.elapsed_time_ns_s1_5 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ;
    wire \current_shift_inst.elapsed_time_ns_s1_6 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ;
    wire \current_shift_inst.elapsed_time_ns_s1_7 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ;
    wire \current_shift_inst.elapsed_time_ns_s1_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ;
    wire \current_shift_inst.elapsed_time_ns_s1_9 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ;
    wire \current_shift_inst.elapsed_time_ns_s1_10 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ;
    wire \current_shift_inst.elapsed_time_ns_s1_11 ;
    wire bfn_18_19_0_;
    wire \current_shift_inst.elapsed_time_ns_s1_12 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ;
    wire \current_shift_inst.elapsed_time_ns_s1_13 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ;
    wire \current_shift_inst.elapsed_time_ns_s1_14 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ;
    wire \current_shift_inst.elapsed_time_ns_s1_15 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ;
    wire \current_shift_inst.elapsed_time_ns_s1_16 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ;
    wire \current_shift_inst.elapsed_time_ns_s1_17 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ;
    wire \current_shift_inst.elapsed_time_ns_s1_18 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ;
    wire \current_shift_inst.elapsed_time_ns_s1_19 ;
    wire bfn_18_20_0_;
    wire \current_shift_inst.elapsed_time_ns_s1_20 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ;
    wire \current_shift_inst.elapsed_time_ns_s1_21 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ;
    wire \current_shift_inst.elapsed_time_ns_s1_22 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ;
    wire \current_shift_inst.elapsed_time_ns_s1_23 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ;
    wire \current_shift_inst.elapsed_time_ns_s1_24 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ;
    wire \current_shift_inst.elapsed_time_ns_s1_25 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ;
    wire \current_shift_inst.elapsed_time_ns_s1_26 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ;
    wire \current_shift_inst.elapsed_time_ns_s1_27 ;
    wire bfn_18_21_0_;
    wire \current_shift_inst.elapsed_time_ns_s1_28 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ;
    wire \current_shift_inst.elapsed_time_ns_s1_29 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ;
    wire \current_shift_inst.elapsed_time_ns_s1_30 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ;
    wire \current_shift_inst.timer_s1.N_180_i_g ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ;
    wire \current_shift_inst.timer_s1.counterZ0Z_0 ;
    wire bfn_18_22_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_1 ;
    wire \current_shift_inst.timer_s1.counter_cry_0 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_2 ;
    wire \current_shift_inst.timer_s1.counter_cry_1 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_3 ;
    wire \current_shift_inst.timer_s1.counter_cry_2 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_4 ;
    wire \current_shift_inst.timer_s1.counter_cry_3 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_5 ;
    wire \current_shift_inst.timer_s1.counter_cry_4 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_5 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_7 ;
    wire \current_shift_inst.timer_s1.counter_cry_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_7 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_8 ;
    wire bfn_18_23_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_9 ;
    wire \current_shift_inst.timer_s1.counter_cry_8 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_10 ;
    wire \current_shift_inst.timer_s1.counter_cry_9 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_11 ;
    wire \current_shift_inst.timer_s1.counter_cry_10 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_12 ;
    wire \current_shift_inst.timer_s1.counter_cry_11 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_13 ;
    wire \current_shift_inst.timer_s1.counter_cry_12 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_13 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_15 ;
    wire \current_shift_inst.timer_s1.counter_cry_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_15 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_16 ;
    wire bfn_18_24_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_17 ;
    wire \current_shift_inst.timer_s1.counter_cry_16 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_18 ;
    wire \current_shift_inst.timer_s1.counter_cry_17 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_19 ;
    wire \current_shift_inst.timer_s1.counter_cry_18 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_20 ;
    wire \current_shift_inst.timer_s1.counter_cry_19 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_21 ;
    wire \current_shift_inst.timer_s1.counter_cry_20 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_21 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_23 ;
    wire \current_shift_inst.timer_s1.counter_cry_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_23 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_24 ;
    wire bfn_18_25_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_25 ;
    wire \current_shift_inst.timer_s1.counter_cry_24 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_26 ;
    wire \current_shift_inst.timer_s1.counter_cry_25 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_27 ;
    wire \current_shift_inst.timer_s1.counter_cry_26 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_28 ;
    wire \current_shift_inst.timer_s1.counter_cry_27 ;
    wire \current_shift_inst.timer_s1.running_i ;
    wire \current_shift_inst.timer_s1.counter_cry_28 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_29 ;
    wire \current_shift_inst.timer_s1.N_181_i_g ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ;
    wire \delay_measurement_inst.elapsed_time_tr_1 ;
    wire _gnd_net_;
    wire clk_100mhz_0;
    wire \delay_measurement_inst.delay_tr_timer.N_304_i_g ;
    wire red_c_g;

    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .TEST_MODE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FILTER_RANGE=3'b001;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVR=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVQ=3'b011;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVF=7'b1000010;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__23836),
            .RESETB(N__36395),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(clk_100mhz_0));
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__38398),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__38388),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15}),
            .ADDSUBBOT(),
            .A({dangling_wire_16,N__21505,N__21508,N__21506,N__21509,N__21507,N__19943,N__19966,N__20000,N__19925,N__19987,N__20902,N__20933,N__20020,N__20035,N__20050}),
            .C({dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31,dangling_wire_32}),
            .B({dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,N__38394,N__38391,dangling_wire_40,dangling_wire_41,dangling_wire_42,N__38389,N__38393,N__38390,N__38392}),
            .OHOLDTOP(),
            .O({dangling_wire_43,dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,dangling_wire_48,\pwm_generator_inst.un2_threshold_acc_1_25 ,\pwm_generator_inst.un2_threshold_acc_1_24 ,\pwm_generator_inst.un2_threshold_acc_1_23 ,\pwm_generator_inst.un2_threshold_acc_1_22 ,\pwm_generator_inst.un2_threshold_acc_1_21 ,\pwm_generator_inst.un2_threshold_acc_1_20 ,\pwm_generator_inst.un2_threshold_acc_1_19 ,\pwm_generator_inst.un2_threshold_acc_1_18 ,\pwm_generator_inst.un2_threshold_acc_1_17 ,\pwm_generator_inst.un2_threshold_acc_1_16 ,\pwm_generator_inst.un2_threshold_acc_1_15 ,\pwm_generator_inst.O_14 ,\pwm_generator_inst.O_13 ,\pwm_generator_inst.O_12 ,\pwm_generator_inst.un3_threshold_acc ,\pwm_generator_inst.O_10 ,\pwm_generator_inst.O_9 ,\pwm_generator_inst.O_8 ,\pwm_generator_inst.O_7 ,\pwm_generator_inst.O_6 ,\pwm_generator_inst.O_5 ,\pwm_generator_inst.O_4 ,\pwm_generator_inst.O_3 ,\pwm_generator_inst.O_2 ,\pwm_generator_inst.O_1 ,\pwm_generator_inst.O_0 }));
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__38279),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__38362),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64}),
            .ADDSUBBOT(),
            .A({dangling_wire_65,N__21608,N__21600,N__21606,N__21599,N__21607,N__21598,N__21609,N__21595,N__21602,N__21594,N__21603,N__21596,N__21604,N__21597,N__21605}),
            .C({dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73,dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81}),
            .B({dangling_wire_82,dangling_wire_83,dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,N__38368,N__38365,dangling_wire_89,dangling_wire_90,dangling_wire_91,N__38363,N__38367,N__38364,N__38366}),
            .OHOLDTOP(),
            .O({dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,\pwm_generator_inst.un2_threshold_acc_2_1_16 ,\pwm_generator_inst.un2_threshold_acc_2_1_15 ,\pwm_generator_inst.un2_threshold_acc_2_14 ,\pwm_generator_inst.un2_threshold_acc_2_13 ,\pwm_generator_inst.un2_threshold_acc_2_12 ,\pwm_generator_inst.un2_threshold_acc_2_11 ,\pwm_generator_inst.un2_threshold_acc_2_10 ,\pwm_generator_inst.un2_threshold_acc_2_9 ,\pwm_generator_inst.un2_threshold_acc_2_8 ,\pwm_generator_inst.un2_threshold_acc_2_7 ,\pwm_generator_inst.un2_threshold_acc_2_6 ,\pwm_generator_inst.un2_threshold_acc_2_5 ,\pwm_generator_inst.un2_threshold_acc_2_4 ,\pwm_generator_inst.un2_threshold_acc_2_3 ,\pwm_generator_inst.un2_threshold_acc_2_2 ,\pwm_generator_inst.un2_threshold_acc_2_1 ,\pwm_generator_inst.un2_threshold_acc_2_0 }));
    PRE_IO_GBUF reset_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__50759),
            .GLOBALBUFFEROUTPUT(red_c_g));
    IO_PAD reset_ibuf_gb_io_iopad (
            .OE(N__50761),
            .DIN(N__50760),
            .DOUT(N__50759),
            .PACKAGEPIN(reset));
    defparam reset_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam reset_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO reset_ibuf_gb_io_preio (
            .PADOEN(N__50761),
            .PADOUT(N__50760),
            .PADIN(N__50759),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_output_obuf_iopad (
            .OE(N__50750),
            .DIN(N__50749),
            .DOUT(N__50748),
            .PACKAGEPIN(pwm_output));
    defparam pwm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam pwm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO pwm_output_obuf_preio (
            .PADOEN(N__50750),
            .PADOUT(N__50749),
            .PADIN(N__50748),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__22012),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp1_ibuf_iopad (
            .OE(N__50741),
            .DIN(N__50740),
            .DOUT(N__50739),
            .PACKAGEPIN(il_max_comp1));
    defparam il_max_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp1_ibuf_preio (
            .PADOEN(N__50741),
            .PADOUT(N__50740),
            .PADIN(N__50739),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s2_phy_obuf_iopad (
            .OE(N__50732),
            .DIN(N__50731),
            .DOUT(N__50730),
            .PACKAGEPIN(s2_phy));
    defparam s2_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s2_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s2_phy_obuf_preio (
            .PADOEN(N__50732),
            .PADOUT(N__50731),
            .PADIN(N__50730),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__26020),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_hc_input_ibuf_iopad (
            .OE(N__50723),
            .DIN(N__50722),
            .DOUT(N__50721),
            .PACKAGEPIN(delay_hc_input));
    defparam delay_hc_input_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam delay_hc_input_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_hc_input_ibuf_preio (
            .PADOEN(N__50723),
            .PADOUT(N__50722),
            .PADIN(N__50721),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_hc_input_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_tr_input_ibuf_iopad (
            .OE(N__50714),
            .DIN(N__50713),
            .DOUT(N__50712),
            .PACKAGEPIN(delay_tr_input));
    defparam delay_tr_input_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam delay_tr_input_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_tr_input_ibuf_preio (
            .PADOEN(N__50714),
            .PADOUT(N__50713),
            .PADIN(N__50712),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_tr_input_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp2_ibuf_iopad (
            .OE(N__50705),
            .DIN(N__50704),
            .DOUT(N__50703),
            .PACKAGEPIN(il_min_comp2));
    defparam il_min_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp2_ibuf_preio (
            .PADOEN(N__50705),
            .PADOUT(N__50704),
            .PADIN(N__50703),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s1_phy_obuf_iopad (
            .OE(N__50696),
            .DIN(N__50695),
            .DOUT(N__50694),
            .PACKAGEPIN(s1_phy));
    defparam s1_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s1_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s1_phy_obuf_preio (
            .PADOEN(N__50696),
            .PADOUT(N__50695),
            .PADIN(N__50694),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__32089),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s4_phy_obuf_iopad (
            .OE(N__50687),
            .DIN(N__50686),
            .DOUT(N__50685),
            .PACKAGEPIN(s4_phy));
    defparam s4_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s4_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s4_phy_obuf_preio (
            .PADOEN(N__50687),
            .PADOUT(N__50686),
            .PADIN(N__50685),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__22657),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp1_ibuf_iopad (
            .OE(N__50678),
            .DIN(N__50677),
            .DOUT(N__50676),
            .PACKAGEPIN(il_min_comp1));
    defparam il_min_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp1_ibuf_preio (
            .PADOEN(N__50678),
            .PADOUT(N__50677),
            .PADIN(N__50676),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s3_phy_obuf_iopad (
            .OE(N__50669),
            .DIN(N__50668),
            .DOUT(N__50667),
            .PACKAGEPIN(s3_phy));
    defparam s3_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s3_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s3_phy_obuf_preio (
            .PADOEN(N__50669),
            .PADOUT(N__50668),
            .PADIN(N__50667),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__26071),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD start_stop_ibuf_iopad (
            .OE(N__50660),
            .DIN(N__50659),
            .DOUT(N__50658),
            .PACKAGEPIN(start_stop));
    defparam start_stop_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam start_stop_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO start_stop_ibuf_preio (
            .PADOEN(N__50660),
            .PADOUT(N__50659),
            .PADIN(N__50658),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(start_stop_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp2_ibuf_iopad (
            .OE(N__50651),
            .DIN(N__50650),
            .DOUT(N__50649),
            .PACKAGEPIN(il_max_comp2));
    defparam il_max_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp2_ibuf_preio (
            .PADOEN(N__50651),
            .PADOUT(N__50650),
            .PADIN(N__50649),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__11973 (
            .O(N__50632),
            .I(N__50628));
    InMux I__11972 (
            .O(N__50631),
            .I(N__50625));
    LocalMux I__11971 (
            .O(N__50628),
            .I(N__50619));
    LocalMux I__11970 (
            .O(N__50625),
            .I(N__50619));
    InMux I__11969 (
            .O(N__50624),
            .I(N__50616));
    Span4Mux_v I__11968 (
            .O(N__50619),
            .I(N__50613));
    LocalMux I__11967 (
            .O(N__50616),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    Odrv4 I__11966 (
            .O(N__50613),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    InMux I__11965 (
            .O(N__50608),
            .I(\current_shift_inst.timer_s1.counter_cry_24 ));
    CascadeMux I__11964 (
            .O(N__50605),
            .I(N__50601));
    CascadeMux I__11963 (
            .O(N__50604),
            .I(N__50598));
    InMux I__11962 (
            .O(N__50601),
            .I(N__50592));
    InMux I__11961 (
            .O(N__50598),
            .I(N__50592));
    InMux I__11960 (
            .O(N__50597),
            .I(N__50589));
    LocalMux I__11959 (
            .O(N__50592),
            .I(N__50586));
    LocalMux I__11958 (
            .O(N__50589),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    Odrv12 I__11957 (
            .O(N__50586),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    InMux I__11956 (
            .O(N__50581),
            .I(\current_shift_inst.timer_s1.counter_cry_25 ));
    CascadeMux I__11955 (
            .O(N__50578),
            .I(N__50574));
    CascadeMux I__11954 (
            .O(N__50577),
            .I(N__50571));
    InMux I__11953 (
            .O(N__50574),
            .I(N__50565));
    InMux I__11952 (
            .O(N__50571),
            .I(N__50565));
    InMux I__11951 (
            .O(N__50570),
            .I(N__50562));
    LocalMux I__11950 (
            .O(N__50565),
            .I(N__50559));
    LocalMux I__11949 (
            .O(N__50562),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    Odrv12 I__11948 (
            .O(N__50559),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    InMux I__11947 (
            .O(N__50554),
            .I(\current_shift_inst.timer_s1.counter_cry_26 ));
    InMux I__11946 (
            .O(N__50551),
            .I(N__50547));
    InMux I__11945 (
            .O(N__50550),
            .I(N__50544));
    LocalMux I__11944 (
            .O(N__50547),
            .I(N__50541));
    LocalMux I__11943 (
            .O(N__50544),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    Odrv12 I__11942 (
            .O(N__50541),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    InMux I__11941 (
            .O(N__50536),
            .I(\current_shift_inst.timer_s1.counter_cry_27 ));
    InMux I__11940 (
            .O(N__50533),
            .I(N__50499));
    InMux I__11939 (
            .O(N__50532),
            .I(N__50499));
    InMux I__11938 (
            .O(N__50531),
            .I(N__50490));
    InMux I__11937 (
            .O(N__50530),
            .I(N__50490));
    InMux I__11936 (
            .O(N__50529),
            .I(N__50490));
    InMux I__11935 (
            .O(N__50528),
            .I(N__50490));
    InMux I__11934 (
            .O(N__50527),
            .I(N__50481));
    InMux I__11933 (
            .O(N__50526),
            .I(N__50481));
    InMux I__11932 (
            .O(N__50525),
            .I(N__50481));
    InMux I__11931 (
            .O(N__50524),
            .I(N__50481));
    InMux I__11930 (
            .O(N__50523),
            .I(N__50472));
    InMux I__11929 (
            .O(N__50522),
            .I(N__50472));
    InMux I__11928 (
            .O(N__50521),
            .I(N__50472));
    InMux I__11927 (
            .O(N__50520),
            .I(N__50472));
    InMux I__11926 (
            .O(N__50519),
            .I(N__50463));
    InMux I__11925 (
            .O(N__50518),
            .I(N__50463));
    InMux I__11924 (
            .O(N__50517),
            .I(N__50463));
    InMux I__11923 (
            .O(N__50516),
            .I(N__50463));
    InMux I__11922 (
            .O(N__50515),
            .I(N__50454));
    InMux I__11921 (
            .O(N__50514),
            .I(N__50454));
    InMux I__11920 (
            .O(N__50513),
            .I(N__50454));
    InMux I__11919 (
            .O(N__50512),
            .I(N__50454));
    InMux I__11918 (
            .O(N__50511),
            .I(N__50445));
    InMux I__11917 (
            .O(N__50510),
            .I(N__50445));
    InMux I__11916 (
            .O(N__50509),
            .I(N__50445));
    InMux I__11915 (
            .O(N__50508),
            .I(N__50445));
    InMux I__11914 (
            .O(N__50507),
            .I(N__50436));
    InMux I__11913 (
            .O(N__50506),
            .I(N__50436));
    InMux I__11912 (
            .O(N__50505),
            .I(N__50436));
    InMux I__11911 (
            .O(N__50504),
            .I(N__50436));
    LocalMux I__11910 (
            .O(N__50499),
            .I(N__50427));
    LocalMux I__11909 (
            .O(N__50490),
            .I(N__50427));
    LocalMux I__11908 (
            .O(N__50481),
            .I(N__50427));
    LocalMux I__11907 (
            .O(N__50472),
            .I(N__50427));
    LocalMux I__11906 (
            .O(N__50463),
            .I(N__50418));
    LocalMux I__11905 (
            .O(N__50454),
            .I(N__50418));
    LocalMux I__11904 (
            .O(N__50445),
            .I(N__50418));
    LocalMux I__11903 (
            .O(N__50436),
            .I(N__50418));
    Span4Mux_v I__11902 (
            .O(N__50427),
            .I(N__50413));
    Span4Mux_v I__11901 (
            .O(N__50418),
            .I(N__50413));
    Odrv4 I__11900 (
            .O(N__50413),
            .I(\current_shift_inst.timer_s1.running_i ));
    InMux I__11899 (
            .O(N__50410),
            .I(\current_shift_inst.timer_s1.counter_cry_28 ));
    InMux I__11898 (
            .O(N__50407),
            .I(N__50404));
    LocalMux I__11897 (
            .O(N__50404),
            .I(N__50400));
    InMux I__11896 (
            .O(N__50403),
            .I(N__50397));
    Span4Mux_h I__11895 (
            .O(N__50400),
            .I(N__50394));
    LocalMux I__11894 (
            .O(N__50397),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    Odrv4 I__11893 (
            .O(N__50394),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    CEMux I__11892 (
            .O(N__50389),
            .I(N__50386));
    LocalMux I__11891 (
            .O(N__50386),
            .I(N__50380));
    CEMux I__11890 (
            .O(N__50385),
            .I(N__50377));
    CEMux I__11889 (
            .O(N__50384),
            .I(N__50374));
    CEMux I__11888 (
            .O(N__50383),
            .I(N__50371));
    Span4Mux_v I__11887 (
            .O(N__50380),
            .I(N__50368));
    LocalMux I__11886 (
            .O(N__50377),
            .I(N__50365));
    LocalMux I__11885 (
            .O(N__50374),
            .I(N__50362));
    LocalMux I__11884 (
            .O(N__50371),
            .I(N__50359));
    Span4Mux_h I__11883 (
            .O(N__50368),
            .I(N__50354));
    Span4Mux_v I__11882 (
            .O(N__50365),
            .I(N__50354));
    Span4Mux_h I__11881 (
            .O(N__50362),
            .I(N__50351));
    Span4Mux_h I__11880 (
            .O(N__50359),
            .I(N__50348));
    Span4Mux_h I__11879 (
            .O(N__50354),
            .I(N__50345));
    Span4Mux_h I__11878 (
            .O(N__50351),
            .I(N__50342));
    Span4Mux_h I__11877 (
            .O(N__50348),
            .I(N__50339));
    Odrv4 I__11876 (
            .O(N__50345),
            .I(\current_shift_inst.timer_s1.N_181_i_g ));
    Odrv4 I__11875 (
            .O(N__50342),
            .I(\current_shift_inst.timer_s1.N_181_i_g ));
    Odrv4 I__11874 (
            .O(N__50339),
            .I(\current_shift_inst.timer_s1.N_181_i_g ));
    InMux I__11873 (
            .O(N__50332),
            .I(N__50329));
    LocalMux I__11872 (
            .O(N__50329),
            .I(N__50325));
    InMux I__11871 (
            .O(N__50328),
            .I(N__50322));
    Span4Mux_h I__11870 (
            .O(N__50325),
            .I(N__50318));
    LocalMux I__11869 (
            .O(N__50322),
            .I(N__50315));
    InMux I__11868 (
            .O(N__50321),
            .I(N__50312));
    Odrv4 I__11867 (
            .O(N__50318),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    Odrv4 I__11866 (
            .O(N__50315),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__11865 (
            .O(N__50312),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    InMux I__11864 (
            .O(N__50305),
            .I(N__50301));
    CascadeMux I__11863 (
            .O(N__50304),
            .I(N__50298));
    LocalMux I__11862 (
            .O(N__50301),
            .I(N__50295));
    InMux I__11861 (
            .O(N__50298),
            .I(N__50292));
    Span4Mux_v I__11860 (
            .O(N__50295),
            .I(N__50287));
    LocalMux I__11859 (
            .O(N__50292),
            .I(N__50287));
    Span4Mux_h I__11858 (
            .O(N__50287),
            .I(N__50284));
    Span4Mux_h I__11857 (
            .O(N__50284),
            .I(N__50281));
    Odrv4 I__11856 (
            .O(N__50281),
            .I(\delay_measurement_inst.elapsed_time_tr_1 ));
    ClkMux I__11855 (
            .O(N__50278),
            .I(N__49819));
    ClkMux I__11854 (
            .O(N__50277),
            .I(N__49819));
    ClkMux I__11853 (
            .O(N__50276),
            .I(N__49819));
    ClkMux I__11852 (
            .O(N__50275),
            .I(N__49819));
    ClkMux I__11851 (
            .O(N__50274),
            .I(N__49819));
    ClkMux I__11850 (
            .O(N__50273),
            .I(N__49819));
    ClkMux I__11849 (
            .O(N__50272),
            .I(N__49819));
    ClkMux I__11848 (
            .O(N__50271),
            .I(N__49819));
    ClkMux I__11847 (
            .O(N__50270),
            .I(N__49819));
    ClkMux I__11846 (
            .O(N__50269),
            .I(N__49819));
    ClkMux I__11845 (
            .O(N__50268),
            .I(N__49819));
    ClkMux I__11844 (
            .O(N__50267),
            .I(N__49819));
    ClkMux I__11843 (
            .O(N__50266),
            .I(N__49819));
    ClkMux I__11842 (
            .O(N__50265),
            .I(N__49819));
    ClkMux I__11841 (
            .O(N__50264),
            .I(N__49819));
    ClkMux I__11840 (
            .O(N__50263),
            .I(N__49819));
    ClkMux I__11839 (
            .O(N__50262),
            .I(N__49819));
    ClkMux I__11838 (
            .O(N__50261),
            .I(N__49819));
    ClkMux I__11837 (
            .O(N__50260),
            .I(N__49819));
    ClkMux I__11836 (
            .O(N__50259),
            .I(N__49819));
    ClkMux I__11835 (
            .O(N__50258),
            .I(N__49819));
    ClkMux I__11834 (
            .O(N__50257),
            .I(N__49819));
    ClkMux I__11833 (
            .O(N__50256),
            .I(N__49819));
    ClkMux I__11832 (
            .O(N__50255),
            .I(N__49819));
    ClkMux I__11831 (
            .O(N__50254),
            .I(N__49819));
    ClkMux I__11830 (
            .O(N__50253),
            .I(N__49819));
    ClkMux I__11829 (
            .O(N__50252),
            .I(N__49819));
    ClkMux I__11828 (
            .O(N__50251),
            .I(N__49819));
    ClkMux I__11827 (
            .O(N__50250),
            .I(N__49819));
    ClkMux I__11826 (
            .O(N__50249),
            .I(N__49819));
    ClkMux I__11825 (
            .O(N__50248),
            .I(N__49819));
    ClkMux I__11824 (
            .O(N__50247),
            .I(N__49819));
    ClkMux I__11823 (
            .O(N__50246),
            .I(N__49819));
    ClkMux I__11822 (
            .O(N__50245),
            .I(N__49819));
    ClkMux I__11821 (
            .O(N__50244),
            .I(N__49819));
    ClkMux I__11820 (
            .O(N__50243),
            .I(N__49819));
    ClkMux I__11819 (
            .O(N__50242),
            .I(N__49819));
    ClkMux I__11818 (
            .O(N__50241),
            .I(N__49819));
    ClkMux I__11817 (
            .O(N__50240),
            .I(N__49819));
    ClkMux I__11816 (
            .O(N__50239),
            .I(N__49819));
    ClkMux I__11815 (
            .O(N__50238),
            .I(N__49819));
    ClkMux I__11814 (
            .O(N__50237),
            .I(N__49819));
    ClkMux I__11813 (
            .O(N__50236),
            .I(N__49819));
    ClkMux I__11812 (
            .O(N__50235),
            .I(N__49819));
    ClkMux I__11811 (
            .O(N__50234),
            .I(N__49819));
    ClkMux I__11810 (
            .O(N__50233),
            .I(N__49819));
    ClkMux I__11809 (
            .O(N__50232),
            .I(N__49819));
    ClkMux I__11808 (
            .O(N__50231),
            .I(N__49819));
    ClkMux I__11807 (
            .O(N__50230),
            .I(N__49819));
    ClkMux I__11806 (
            .O(N__50229),
            .I(N__49819));
    ClkMux I__11805 (
            .O(N__50228),
            .I(N__49819));
    ClkMux I__11804 (
            .O(N__50227),
            .I(N__49819));
    ClkMux I__11803 (
            .O(N__50226),
            .I(N__49819));
    ClkMux I__11802 (
            .O(N__50225),
            .I(N__49819));
    ClkMux I__11801 (
            .O(N__50224),
            .I(N__49819));
    ClkMux I__11800 (
            .O(N__50223),
            .I(N__49819));
    ClkMux I__11799 (
            .O(N__50222),
            .I(N__49819));
    ClkMux I__11798 (
            .O(N__50221),
            .I(N__49819));
    ClkMux I__11797 (
            .O(N__50220),
            .I(N__49819));
    ClkMux I__11796 (
            .O(N__50219),
            .I(N__49819));
    ClkMux I__11795 (
            .O(N__50218),
            .I(N__49819));
    ClkMux I__11794 (
            .O(N__50217),
            .I(N__49819));
    ClkMux I__11793 (
            .O(N__50216),
            .I(N__49819));
    ClkMux I__11792 (
            .O(N__50215),
            .I(N__49819));
    ClkMux I__11791 (
            .O(N__50214),
            .I(N__49819));
    ClkMux I__11790 (
            .O(N__50213),
            .I(N__49819));
    ClkMux I__11789 (
            .O(N__50212),
            .I(N__49819));
    ClkMux I__11788 (
            .O(N__50211),
            .I(N__49819));
    ClkMux I__11787 (
            .O(N__50210),
            .I(N__49819));
    ClkMux I__11786 (
            .O(N__50209),
            .I(N__49819));
    ClkMux I__11785 (
            .O(N__50208),
            .I(N__49819));
    ClkMux I__11784 (
            .O(N__50207),
            .I(N__49819));
    ClkMux I__11783 (
            .O(N__50206),
            .I(N__49819));
    ClkMux I__11782 (
            .O(N__50205),
            .I(N__49819));
    ClkMux I__11781 (
            .O(N__50204),
            .I(N__49819));
    ClkMux I__11780 (
            .O(N__50203),
            .I(N__49819));
    ClkMux I__11779 (
            .O(N__50202),
            .I(N__49819));
    ClkMux I__11778 (
            .O(N__50201),
            .I(N__49819));
    ClkMux I__11777 (
            .O(N__50200),
            .I(N__49819));
    ClkMux I__11776 (
            .O(N__50199),
            .I(N__49819));
    ClkMux I__11775 (
            .O(N__50198),
            .I(N__49819));
    ClkMux I__11774 (
            .O(N__50197),
            .I(N__49819));
    ClkMux I__11773 (
            .O(N__50196),
            .I(N__49819));
    ClkMux I__11772 (
            .O(N__50195),
            .I(N__49819));
    ClkMux I__11771 (
            .O(N__50194),
            .I(N__49819));
    ClkMux I__11770 (
            .O(N__50193),
            .I(N__49819));
    ClkMux I__11769 (
            .O(N__50192),
            .I(N__49819));
    ClkMux I__11768 (
            .O(N__50191),
            .I(N__49819));
    ClkMux I__11767 (
            .O(N__50190),
            .I(N__49819));
    ClkMux I__11766 (
            .O(N__50189),
            .I(N__49819));
    ClkMux I__11765 (
            .O(N__50188),
            .I(N__49819));
    ClkMux I__11764 (
            .O(N__50187),
            .I(N__49819));
    ClkMux I__11763 (
            .O(N__50186),
            .I(N__49819));
    ClkMux I__11762 (
            .O(N__50185),
            .I(N__49819));
    ClkMux I__11761 (
            .O(N__50184),
            .I(N__49819));
    ClkMux I__11760 (
            .O(N__50183),
            .I(N__49819));
    ClkMux I__11759 (
            .O(N__50182),
            .I(N__49819));
    ClkMux I__11758 (
            .O(N__50181),
            .I(N__49819));
    ClkMux I__11757 (
            .O(N__50180),
            .I(N__49819));
    ClkMux I__11756 (
            .O(N__50179),
            .I(N__49819));
    ClkMux I__11755 (
            .O(N__50178),
            .I(N__49819));
    ClkMux I__11754 (
            .O(N__50177),
            .I(N__49819));
    ClkMux I__11753 (
            .O(N__50176),
            .I(N__49819));
    ClkMux I__11752 (
            .O(N__50175),
            .I(N__49819));
    ClkMux I__11751 (
            .O(N__50174),
            .I(N__49819));
    ClkMux I__11750 (
            .O(N__50173),
            .I(N__49819));
    ClkMux I__11749 (
            .O(N__50172),
            .I(N__49819));
    ClkMux I__11748 (
            .O(N__50171),
            .I(N__49819));
    ClkMux I__11747 (
            .O(N__50170),
            .I(N__49819));
    ClkMux I__11746 (
            .O(N__50169),
            .I(N__49819));
    ClkMux I__11745 (
            .O(N__50168),
            .I(N__49819));
    ClkMux I__11744 (
            .O(N__50167),
            .I(N__49819));
    ClkMux I__11743 (
            .O(N__50166),
            .I(N__49819));
    ClkMux I__11742 (
            .O(N__50165),
            .I(N__49819));
    ClkMux I__11741 (
            .O(N__50164),
            .I(N__49819));
    ClkMux I__11740 (
            .O(N__50163),
            .I(N__49819));
    ClkMux I__11739 (
            .O(N__50162),
            .I(N__49819));
    ClkMux I__11738 (
            .O(N__50161),
            .I(N__49819));
    ClkMux I__11737 (
            .O(N__50160),
            .I(N__49819));
    ClkMux I__11736 (
            .O(N__50159),
            .I(N__49819));
    ClkMux I__11735 (
            .O(N__50158),
            .I(N__49819));
    ClkMux I__11734 (
            .O(N__50157),
            .I(N__49819));
    ClkMux I__11733 (
            .O(N__50156),
            .I(N__49819));
    ClkMux I__11732 (
            .O(N__50155),
            .I(N__49819));
    ClkMux I__11731 (
            .O(N__50154),
            .I(N__49819));
    ClkMux I__11730 (
            .O(N__50153),
            .I(N__49819));
    ClkMux I__11729 (
            .O(N__50152),
            .I(N__49819));
    ClkMux I__11728 (
            .O(N__50151),
            .I(N__49819));
    ClkMux I__11727 (
            .O(N__50150),
            .I(N__49819));
    ClkMux I__11726 (
            .O(N__50149),
            .I(N__49819));
    ClkMux I__11725 (
            .O(N__50148),
            .I(N__49819));
    ClkMux I__11724 (
            .O(N__50147),
            .I(N__49819));
    ClkMux I__11723 (
            .O(N__50146),
            .I(N__49819));
    ClkMux I__11722 (
            .O(N__50145),
            .I(N__49819));
    ClkMux I__11721 (
            .O(N__50144),
            .I(N__49819));
    ClkMux I__11720 (
            .O(N__50143),
            .I(N__49819));
    ClkMux I__11719 (
            .O(N__50142),
            .I(N__49819));
    ClkMux I__11718 (
            .O(N__50141),
            .I(N__49819));
    ClkMux I__11717 (
            .O(N__50140),
            .I(N__49819));
    ClkMux I__11716 (
            .O(N__50139),
            .I(N__49819));
    ClkMux I__11715 (
            .O(N__50138),
            .I(N__49819));
    ClkMux I__11714 (
            .O(N__50137),
            .I(N__49819));
    ClkMux I__11713 (
            .O(N__50136),
            .I(N__49819));
    ClkMux I__11712 (
            .O(N__50135),
            .I(N__49819));
    ClkMux I__11711 (
            .O(N__50134),
            .I(N__49819));
    ClkMux I__11710 (
            .O(N__50133),
            .I(N__49819));
    ClkMux I__11709 (
            .O(N__50132),
            .I(N__49819));
    ClkMux I__11708 (
            .O(N__50131),
            .I(N__49819));
    ClkMux I__11707 (
            .O(N__50130),
            .I(N__49819));
    ClkMux I__11706 (
            .O(N__50129),
            .I(N__49819));
    ClkMux I__11705 (
            .O(N__50128),
            .I(N__49819));
    ClkMux I__11704 (
            .O(N__50127),
            .I(N__49819));
    ClkMux I__11703 (
            .O(N__50126),
            .I(N__49819));
    GlobalMux I__11702 (
            .O(N__49819),
            .I(clk_100mhz_0));
    CEMux I__11701 (
            .O(N__49816),
            .I(N__49798));
    CEMux I__11700 (
            .O(N__49815),
            .I(N__49798));
    CEMux I__11699 (
            .O(N__49814),
            .I(N__49798));
    CEMux I__11698 (
            .O(N__49813),
            .I(N__49798));
    CEMux I__11697 (
            .O(N__49812),
            .I(N__49798));
    CEMux I__11696 (
            .O(N__49811),
            .I(N__49798));
    GlobalMux I__11695 (
            .O(N__49798),
            .I(N__49795));
    gio2CtrlBuf I__11694 (
            .O(N__49795),
            .I(\delay_measurement_inst.delay_tr_timer.N_304_i_g ));
    CascadeMux I__11693 (
            .O(N__49792),
            .I(N__49783));
    CascadeMux I__11692 (
            .O(N__49791),
            .I(N__49780));
    InMux I__11691 (
            .O(N__49790),
            .I(N__49777));
    InMux I__11690 (
            .O(N__49789),
            .I(N__49774));
    InMux I__11689 (
            .O(N__49788),
            .I(N__49771));
    InMux I__11688 (
            .O(N__49787),
            .I(N__49768));
    InMux I__11687 (
            .O(N__49786),
            .I(N__49765));
    InMux I__11686 (
            .O(N__49783),
            .I(N__49762));
    InMux I__11685 (
            .O(N__49780),
            .I(N__49759));
    LocalMux I__11684 (
            .O(N__49777),
            .I(N__49756));
    LocalMux I__11683 (
            .O(N__49774),
            .I(N__49753));
    LocalMux I__11682 (
            .O(N__49771),
            .I(N__49750));
    LocalMux I__11681 (
            .O(N__49768),
            .I(N__49747));
    LocalMux I__11680 (
            .O(N__49765),
            .I(N__49657));
    LocalMux I__11679 (
            .O(N__49762),
            .I(N__49633));
    LocalMux I__11678 (
            .O(N__49759),
            .I(N__49604));
    Glb2LocalMux I__11677 (
            .O(N__49756),
            .I(N__49318));
    Glb2LocalMux I__11676 (
            .O(N__49753),
            .I(N__49318));
    Glb2LocalMux I__11675 (
            .O(N__49750),
            .I(N__49318));
    Glb2LocalMux I__11674 (
            .O(N__49747),
            .I(N__49318));
    SRMux I__11673 (
            .O(N__49746),
            .I(N__49318));
    SRMux I__11672 (
            .O(N__49745),
            .I(N__49318));
    SRMux I__11671 (
            .O(N__49744),
            .I(N__49318));
    SRMux I__11670 (
            .O(N__49743),
            .I(N__49318));
    SRMux I__11669 (
            .O(N__49742),
            .I(N__49318));
    SRMux I__11668 (
            .O(N__49741),
            .I(N__49318));
    SRMux I__11667 (
            .O(N__49740),
            .I(N__49318));
    SRMux I__11666 (
            .O(N__49739),
            .I(N__49318));
    SRMux I__11665 (
            .O(N__49738),
            .I(N__49318));
    SRMux I__11664 (
            .O(N__49737),
            .I(N__49318));
    SRMux I__11663 (
            .O(N__49736),
            .I(N__49318));
    SRMux I__11662 (
            .O(N__49735),
            .I(N__49318));
    SRMux I__11661 (
            .O(N__49734),
            .I(N__49318));
    SRMux I__11660 (
            .O(N__49733),
            .I(N__49318));
    SRMux I__11659 (
            .O(N__49732),
            .I(N__49318));
    SRMux I__11658 (
            .O(N__49731),
            .I(N__49318));
    SRMux I__11657 (
            .O(N__49730),
            .I(N__49318));
    SRMux I__11656 (
            .O(N__49729),
            .I(N__49318));
    SRMux I__11655 (
            .O(N__49728),
            .I(N__49318));
    SRMux I__11654 (
            .O(N__49727),
            .I(N__49318));
    SRMux I__11653 (
            .O(N__49726),
            .I(N__49318));
    SRMux I__11652 (
            .O(N__49725),
            .I(N__49318));
    SRMux I__11651 (
            .O(N__49724),
            .I(N__49318));
    SRMux I__11650 (
            .O(N__49723),
            .I(N__49318));
    SRMux I__11649 (
            .O(N__49722),
            .I(N__49318));
    SRMux I__11648 (
            .O(N__49721),
            .I(N__49318));
    SRMux I__11647 (
            .O(N__49720),
            .I(N__49318));
    SRMux I__11646 (
            .O(N__49719),
            .I(N__49318));
    SRMux I__11645 (
            .O(N__49718),
            .I(N__49318));
    SRMux I__11644 (
            .O(N__49717),
            .I(N__49318));
    SRMux I__11643 (
            .O(N__49716),
            .I(N__49318));
    SRMux I__11642 (
            .O(N__49715),
            .I(N__49318));
    SRMux I__11641 (
            .O(N__49714),
            .I(N__49318));
    SRMux I__11640 (
            .O(N__49713),
            .I(N__49318));
    SRMux I__11639 (
            .O(N__49712),
            .I(N__49318));
    SRMux I__11638 (
            .O(N__49711),
            .I(N__49318));
    SRMux I__11637 (
            .O(N__49710),
            .I(N__49318));
    SRMux I__11636 (
            .O(N__49709),
            .I(N__49318));
    SRMux I__11635 (
            .O(N__49708),
            .I(N__49318));
    SRMux I__11634 (
            .O(N__49707),
            .I(N__49318));
    SRMux I__11633 (
            .O(N__49706),
            .I(N__49318));
    SRMux I__11632 (
            .O(N__49705),
            .I(N__49318));
    SRMux I__11631 (
            .O(N__49704),
            .I(N__49318));
    SRMux I__11630 (
            .O(N__49703),
            .I(N__49318));
    SRMux I__11629 (
            .O(N__49702),
            .I(N__49318));
    SRMux I__11628 (
            .O(N__49701),
            .I(N__49318));
    SRMux I__11627 (
            .O(N__49700),
            .I(N__49318));
    SRMux I__11626 (
            .O(N__49699),
            .I(N__49318));
    SRMux I__11625 (
            .O(N__49698),
            .I(N__49318));
    SRMux I__11624 (
            .O(N__49697),
            .I(N__49318));
    SRMux I__11623 (
            .O(N__49696),
            .I(N__49318));
    SRMux I__11622 (
            .O(N__49695),
            .I(N__49318));
    SRMux I__11621 (
            .O(N__49694),
            .I(N__49318));
    SRMux I__11620 (
            .O(N__49693),
            .I(N__49318));
    SRMux I__11619 (
            .O(N__49692),
            .I(N__49318));
    SRMux I__11618 (
            .O(N__49691),
            .I(N__49318));
    SRMux I__11617 (
            .O(N__49690),
            .I(N__49318));
    SRMux I__11616 (
            .O(N__49689),
            .I(N__49318));
    SRMux I__11615 (
            .O(N__49688),
            .I(N__49318));
    SRMux I__11614 (
            .O(N__49687),
            .I(N__49318));
    SRMux I__11613 (
            .O(N__49686),
            .I(N__49318));
    SRMux I__11612 (
            .O(N__49685),
            .I(N__49318));
    SRMux I__11611 (
            .O(N__49684),
            .I(N__49318));
    SRMux I__11610 (
            .O(N__49683),
            .I(N__49318));
    SRMux I__11609 (
            .O(N__49682),
            .I(N__49318));
    SRMux I__11608 (
            .O(N__49681),
            .I(N__49318));
    SRMux I__11607 (
            .O(N__49680),
            .I(N__49318));
    SRMux I__11606 (
            .O(N__49679),
            .I(N__49318));
    SRMux I__11605 (
            .O(N__49678),
            .I(N__49318));
    SRMux I__11604 (
            .O(N__49677),
            .I(N__49318));
    SRMux I__11603 (
            .O(N__49676),
            .I(N__49318));
    SRMux I__11602 (
            .O(N__49675),
            .I(N__49318));
    SRMux I__11601 (
            .O(N__49674),
            .I(N__49318));
    SRMux I__11600 (
            .O(N__49673),
            .I(N__49318));
    SRMux I__11599 (
            .O(N__49672),
            .I(N__49318));
    SRMux I__11598 (
            .O(N__49671),
            .I(N__49318));
    SRMux I__11597 (
            .O(N__49670),
            .I(N__49318));
    SRMux I__11596 (
            .O(N__49669),
            .I(N__49318));
    SRMux I__11595 (
            .O(N__49668),
            .I(N__49318));
    SRMux I__11594 (
            .O(N__49667),
            .I(N__49318));
    SRMux I__11593 (
            .O(N__49666),
            .I(N__49318));
    SRMux I__11592 (
            .O(N__49665),
            .I(N__49318));
    SRMux I__11591 (
            .O(N__49664),
            .I(N__49318));
    SRMux I__11590 (
            .O(N__49663),
            .I(N__49318));
    SRMux I__11589 (
            .O(N__49662),
            .I(N__49318));
    SRMux I__11588 (
            .O(N__49661),
            .I(N__49318));
    SRMux I__11587 (
            .O(N__49660),
            .I(N__49318));
    Glb2LocalMux I__11586 (
            .O(N__49657),
            .I(N__49318));
    SRMux I__11585 (
            .O(N__49656),
            .I(N__49318));
    SRMux I__11584 (
            .O(N__49655),
            .I(N__49318));
    SRMux I__11583 (
            .O(N__49654),
            .I(N__49318));
    SRMux I__11582 (
            .O(N__49653),
            .I(N__49318));
    SRMux I__11581 (
            .O(N__49652),
            .I(N__49318));
    SRMux I__11580 (
            .O(N__49651),
            .I(N__49318));
    SRMux I__11579 (
            .O(N__49650),
            .I(N__49318));
    SRMux I__11578 (
            .O(N__49649),
            .I(N__49318));
    SRMux I__11577 (
            .O(N__49648),
            .I(N__49318));
    SRMux I__11576 (
            .O(N__49647),
            .I(N__49318));
    SRMux I__11575 (
            .O(N__49646),
            .I(N__49318));
    SRMux I__11574 (
            .O(N__49645),
            .I(N__49318));
    SRMux I__11573 (
            .O(N__49644),
            .I(N__49318));
    SRMux I__11572 (
            .O(N__49643),
            .I(N__49318));
    SRMux I__11571 (
            .O(N__49642),
            .I(N__49318));
    SRMux I__11570 (
            .O(N__49641),
            .I(N__49318));
    SRMux I__11569 (
            .O(N__49640),
            .I(N__49318));
    SRMux I__11568 (
            .O(N__49639),
            .I(N__49318));
    SRMux I__11567 (
            .O(N__49638),
            .I(N__49318));
    SRMux I__11566 (
            .O(N__49637),
            .I(N__49318));
    SRMux I__11565 (
            .O(N__49636),
            .I(N__49318));
    Glb2LocalMux I__11564 (
            .O(N__49633),
            .I(N__49318));
    SRMux I__11563 (
            .O(N__49632),
            .I(N__49318));
    SRMux I__11562 (
            .O(N__49631),
            .I(N__49318));
    SRMux I__11561 (
            .O(N__49630),
            .I(N__49318));
    SRMux I__11560 (
            .O(N__49629),
            .I(N__49318));
    SRMux I__11559 (
            .O(N__49628),
            .I(N__49318));
    SRMux I__11558 (
            .O(N__49627),
            .I(N__49318));
    SRMux I__11557 (
            .O(N__49626),
            .I(N__49318));
    SRMux I__11556 (
            .O(N__49625),
            .I(N__49318));
    SRMux I__11555 (
            .O(N__49624),
            .I(N__49318));
    SRMux I__11554 (
            .O(N__49623),
            .I(N__49318));
    SRMux I__11553 (
            .O(N__49622),
            .I(N__49318));
    SRMux I__11552 (
            .O(N__49621),
            .I(N__49318));
    SRMux I__11551 (
            .O(N__49620),
            .I(N__49318));
    SRMux I__11550 (
            .O(N__49619),
            .I(N__49318));
    SRMux I__11549 (
            .O(N__49618),
            .I(N__49318));
    SRMux I__11548 (
            .O(N__49617),
            .I(N__49318));
    SRMux I__11547 (
            .O(N__49616),
            .I(N__49318));
    SRMux I__11546 (
            .O(N__49615),
            .I(N__49318));
    SRMux I__11545 (
            .O(N__49614),
            .I(N__49318));
    SRMux I__11544 (
            .O(N__49613),
            .I(N__49318));
    SRMux I__11543 (
            .O(N__49612),
            .I(N__49318));
    SRMux I__11542 (
            .O(N__49611),
            .I(N__49318));
    SRMux I__11541 (
            .O(N__49610),
            .I(N__49318));
    SRMux I__11540 (
            .O(N__49609),
            .I(N__49318));
    SRMux I__11539 (
            .O(N__49608),
            .I(N__49318));
    SRMux I__11538 (
            .O(N__49607),
            .I(N__49318));
    Glb2LocalMux I__11537 (
            .O(N__49604),
            .I(N__49318));
    SRMux I__11536 (
            .O(N__49603),
            .I(N__49318));
    GlobalMux I__11535 (
            .O(N__49318),
            .I(N__49315));
    gio2CtrlBuf I__11534 (
            .O(N__49315),
            .I(red_c_g));
    InMux I__11533 (
            .O(N__49312),
            .I(N__49308));
    InMux I__11532 (
            .O(N__49311),
            .I(N__49305));
    LocalMux I__11531 (
            .O(N__49308),
            .I(N__49299));
    LocalMux I__11530 (
            .O(N__49305),
            .I(N__49299));
    InMux I__11529 (
            .O(N__49304),
            .I(N__49296));
    Span4Mux_v I__11528 (
            .O(N__49299),
            .I(N__49293));
    LocalMux I__11527 (
            .O(N__49296),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    Odrv4 I__11526 (
            .O(N__49293),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    InMux I__11525 (
            .O(N__49288),
            .I(bfn_18_24_0_));
    CascadeMux I__11524 (
            .O(N__49285),
            .I(N__49281));
    InMux I__11523 (
            .O(N__49284),
            .I(N__49278));
    InMux I__11522 (
            .O(N__49281),
            .I(N__49275));
    LocalMux I__11521 (
            .O(N__49278),
            .I(N__49269));
    LocalMux I__11520 (
            .O(N__49275),
            .I(N__49269));
    InMux I__11519 (
            .O(N__49274),
            .I(N__49266));
    Span4Mux_v I__11518 (
            .O(N__49269),
            .I(N__49263));
    LocalMux I__11517 (
            .O(N__49266),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    Odrv4 I__11516 (
            .O(N__49263),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    InMux I__11515 (
            .O(N__49258),
            .I(\current_shift_inst.timer_s1.counter_cry_16 ));
    CascadeMux I__11514 (
            .O(N__49255),
            .I(N__49251));
    CascadeMux I__11513 (
            .O(N__49254),
            .I(N__49248));
    InMux I__11512 (
            .O(N__49251),
            .I(N__49243));
    InMux I__11511 (
            .O(N__49248),
            .I(N__49243));
    LocalMux I__11510 (
            .O(N__49243),
            .I(N__49239));
    InMux I__11509 (
            .O(N__49242),
            .I(N__49236));
    Span4Mux_h I__11508 (
            .O(N__49239),
            .I(N__49233));
    LocalMux I__11507 (
            .O(N__49236),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    Odrv4 I__11506 (
            .O(N__49233),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    InMux I__11505 (
            .O(N__49228),
            .I(\current_shift_inst.timer_s1.counter_cry_17 ));
    CascadeMux I__11504 (
            .O(N__49225),
            .I(N__49221));
    CascadeMux I__11503 (
            .O(N__49224),
            .I(N__49218));
    InMux I__11502 (
            .O(N__49221),
            .I(N__49213));
    InMux I__11501 (
            .O(N__49218),
            .I(N__49213));
    LocalMux I__11500 (
            .O(N__49213),
            .I(N__49209));
    InMux I__11499 (
            .O(N__49212),
            .I(N__49206));
    Span4Mux_h I__11498 (
            .O(N__49209),
            .I(N__49203));
    LocalMux I__11497 (
            .O(N__49206),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    Odrv4 I__11496 (
            .O(N__49203),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    InMux I__11495 (
            .O(N__49198),
            .I(\current_shift_inst.timer_s1.counter_cry_18 ));
    InMux I__11494 (
            .O(N__49195),
            .I(N__49189));
    InMux I__11493 (
            .O(N__49194),
            .I(N__49189));
    LocalMux I__11492 (
            .O(N__49189),
            .I(N__49185));
    InMux I__11491 (
            .O(N__49188),
            .I(N__49182));
    Span4Mux_h I__11490 (
            .O(N__49185),
            .I(N__49179));
    LocalMux I__11489 (
            .O(N__49182),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    Odrv4 I__11488 (
            .O(N__49179),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    InMux I__11487 (
            .O(N__49174),
            .I(\current_shift_inst.timer_s1.counter_cry_19 ));
    InMux I__11486 (
            .O(N__49171),
            .I(N__49165));
    InMux I__11485 (
            .O(N__49170),
            .I(N__49165));
    LocalMux I__11484 (
            .O(N__49165),
            .I(N__49161));
    InMux I__11483 (
            .O(N__49164),
            .I(N__49158));
    Span4Mux_h I__11482 (
            .O(N__49161),
            .I(N__49155));
    LocalMux I__11481 (
            .O(N__49158),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    Odrv4 I__11480 (
            .O(N__49155),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    InMux I__11479 (
            .O(N__49150),
            .I(\current_shift_inst.timer_s1.counter_cry_20 ));
    CascadeMux I__11478 (
            .O(N__49147),
            .I(N__49143));
    CascadeMux I__11477 (
            .O(N__49146),
            .I(N__49140));
    InMux I__11476 (
            .O(N__49143),
            .I(N__49134));
    InMux I__11475 (
            .O(N__49140),
            .I(N__49134));
    InMux I__11474 (
            .O(N__49139),
            .I(N__49131));
    LocalMux I__11473 (
            .O(N__49134),
            .I(N__49128));
    LocalMux I__11472 (
            .O(N__49131),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    Odrv12 I__11471 (
            .O(N__49128),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    InMux I__11470 (
            .O(N__49123),
            .I(\current_shift_inst.timer_s1.counter_cry_21 ));
    CascadeMux I__11469 (
            .O(N__49120),
            .I(N__49116));
    CascadeMux I__11468 (
            .O(N__49119),
            .I(N__49113));
    InMux I__11467 (
            .O(N__49116),
            .I(N__49107));
    InMux I__11466 (
            .O(N__49113),
            .I(N__49107));
    InMux I__11465 (
            .O(N__49112),
            .I(N__49104));
    LocalMux I__11464 (
            .O(N__49107),
            .I(N__49101));
    LocalMux I__11463 (
            .O(N__49104),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    Odrv12 I__11462 (
            .O(N__49101),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    InMux I__11461 (
            .O(N__49096),
            .I(\current_shift_inst.timer_s1.counter_cry_22 ));
    InMux I__11460 (
            .O(N__49093),
            .I(N__49089));
    InMux I__11459 (
            .O(N__49092),
            .I(N__49086));
    LocalMux I__11458 (
            .O(N__49089),
            .I(N__49080));
    LocalMux I__11457 (
            .O(N__49086),
            .I(N__49080));
    InMux I__11456 (
            .O(N__49085),
            .I(N__49077));
    Span4Mux_v I__11455 (
            .O(N__49080),
            .I(N__49074));
    LocalMux I__11454 (
            .O(N__49077),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    Odrv4 I__11453 (
            .O(N__49074),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    InMux I__11452 (
            .O(N__49069),
            .I(bfn_18_25_0_));
    CascadeMux I__11451 (
            .O(N__49066),
            .I(N__49062));
    InMux I__11450 (
            .O(N__49065),
            .I(N__49058));
    InMux I__11449 (
            .O(N__49062),
            .I(N__49055));
    InMux I__11448 (
            .O(N__49061),
            .I(N__49052));
    LocalMux I__11447 (
            .O(N__49058),
            .I(N__49047));
    LocalMux I__11446 (
            .O(N__49055),
            .I(N__49047));
    LocalMux I__11445 (
            .O(N__49052),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    Odrv12 I__11444 (
            .O(N__49047),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    InMux I__11443 (
            .O(N__49042),
            .I(bfn_18_23_0_));
    InMux I__11442 (
            .O(N__49039),
            .I(N__49034));
    InMux I__11441 (
            .O(N__49038),
            .I(N__49031));
    InMux I__11440 (
            .O(N__49037),
            .I(N__49028));
    LocalMux I__11439 (
            .O(N__49034),
            .I(N__49023));
    LocalMux I__11438 (
            .O(N__49031),
            .I(N__49023));
    LocalMux I__11437 (
            .O(N__49028),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    Odrv12 I__11436 (
            .O(N__49023),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    InMux I__11435 (
            .O(N__49018),
            .I(\current_shift_inst.timer_s1.counter_cry_8 ));
    CascadeMux I__11434 (
            .O(N__49015),
            .I(N__49011));
    CascadeMux I__11433 (
            .O(N__49014),
            .I(N__49008));
    InMux I__11432 (
            .O(N__49011),
            .I(N__49002));
    InMux I__11431 (
            .O(N__49008),
            .I(N__49002));
    InMux I__11430 (
            .O(N__49007),
            .I(N__48999));
    LocalMux I__11429 (
            .O(N__49002),
            .I(N__48996));
    LocalMux I__11428 (
            .O(N__48999),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    Odrv12 I__11427 (
            .O(N__48996),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    InMux I__11426 (
            .O(N__48991),
            .I(\current_shift_inst.timer_s1.counter_cry_9 ));
    CascadeMux I__11425 (
            .O(N__48988),
            .I(N__48984));
    CascadeMux I__11424 (
            .O(N__48987),
            .I(N__48981));
    InMux I__11423 (
            .O(N__48984),
            .I(N__48975));
    InMux I__11422 (
            .O(N__48981),
            .I(N__48975));
    InMux I__11421 (
            .O(N__48980),
            .I(N__48972));
    LocalMux I__11420 (
            .O(N__48975),
            .I(N__48969));
    LocalMux I__11419 (
            .O(N__48972),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    Odrv12 I__11418 (
            .O(N__48969),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    InMux I__11417 (
            .O(N__48964),
            .I(\current_shift_inst.timer_s1.counter_cry_10 ));
    InMux I__11416 (
            .O(N__48961),
            .I(N__48955));
    InMux I__11415 (
            .O(N__48960),
            .I(N__48955));
    LocalMux I__11414 (
            .O(N__48955),
            .I(N__48951));
    InMux I__11413 (
            .O(N__48954),
            .I(N__48948));
    Span4Mux_h I__11412 (
            .O(N__48951),
            .I(N__48945));
    LocalMux I__11411 (
            .O(N__48948),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    Odrv4 I__11410 (
            .O(N__48945),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    InMux I__11409 (
            .O(N__48940),
            .I(\current_shift_inst.timer_s1.counter_cry_11 ));
    CascadeMux I__11408 (
            .O(N__48937),
            .I(N__48934));
    InMux I__11407 (
            .O(N__48934),
            .I(N__48930));
    InMux I__11406 (
            .O(N__48933),
            .I(N__48927));
    LocalMux I__11405 (
            .O(N__48930),
            .I(N__48921));
    LocalMux I__11404 (
            .O(N__48927),
            .I(N__48921));
    InMux I__11403 (
            .O(N__48926),
            .I(N__48918));
    Span4Mux_h I__11402 (
            .O(N__48921),
            .I(N__48915));
    LocalMux I__11401 (
            .O(N__48918),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    Odrv4 I__11400 (
            .O(N__48915),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    InMux I__11399 (
            .O(N__48910),
            .I(\current_shift_inst.timer_s1.counter_cry_12 ));
    CascadeMux I__11398 (
            .O(N__48907),
            .I(N__48903));
    CascadeMux I__11397 (
            .O(N__48906),
            .I(N__48900));
    InMux I__11396 (
            .O(N__48903),
            .I(N__48895));
    InMux I__11395 (
            .O(N__48900),
            .I(N__48895));
    LocalMux I__11394 (
            .O(N__48895),
            .I(N__48891));
    InMux I__11393 (
            .O(N__48894),
            .I(N__48888));
    Span4Mux_v I__11392 (
            .O(N__48891),
            .I(N__48885));
    LocalMux I__11391 (
            .O(N__48888),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    Odrv4 I__11390 (
            .O(N__48885),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    InMux I__11389 (
            .O(N__48880),
            .I(\current_shift_inst.timer_s1.counter_cry_13 ));
    InMux I__11388 (
            .O(N__48877),
            .I(N__48870));
    InMux I__11387 (
            .O(N__48876),
            .I(N__48870));
    InMux I__11386 (
            .O(N__48875),
            .I(N__48867));
    LocalMux I__11385 (
            .O(N__48870),
            .I(N__48864));
    LocalMux I__11384 (
            .O(N__48867),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    Odrv12 I__11383 (
            .O(N__48864),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    InMux I__11382 (
            .O(N__48859),
            .I(\current_shift_inst.timer_s1.counter_cry_14 ));
    InMux I__11381 (
            .O(N__48856),
            .I(N__48853));
    LocalMux I__11380 (
            .O(N__48853),
            .I(N__48849));
    InMux I__11379 (
            .O(N__48852),
            .I(N__48846));
    Span4Mux_h I__11378 (
            .O(N__48849),
            .I(N__48842));
    LocalMux I__11377 (
            .O(N__48846),
            .I(N__48839));
    InMux I__11376 (
            .O(N__48845),
            .I(N__48836));
    Span4Mux_v I__11375 (
            .O(N__48842),
            .I(N__48833));
    Span4Mux_h I__11374 (
            .O(N__48839),
            .I(N__48830));
    LocalMux I__11373 (
            .O(N__48836),
            .I(N__48827));
    Span4Mux_h I__11372 (
            .O(N__48833),
            .I(N__48824));
    Span4Mux_h I__11371 (
            .O(N__48830),
            .I(N__48819));
    Span4Mux_v I__11370 (
            .O(N__48827),
            .I(N__48819));
    Odrv4 I__11369 (
            .O(N__48824),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    Odrv4 I__11368 (
            .O(N__48819),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    InMux I__11367 (
            .O(N__48814),
            .I(N__48811));
    LocalMux I__11366 (
            .O(N__48811),
            .I(N__48807));
    CascadeMux I__11365 (
            .O(N__48810),
            .I(N__48804));
    Span4Mux_h I__11364 (
            .O(N__48807),
            .I(N__48801));
    InMux I__11363 (
            .O(N__48804),
            .I(N__48798));
    Span4Mux_v I__11362 (
            .O(N__48801),
            .I(N__48792));
    LocalMux I__11361 (
            .O(N__48798),
            .I(N__48792));
    InMux I__11360 (
            .O(N__48797),
            .I(N__48789));
    Span4Mux_h I__11359 (
            .O(N__48792),
            .I(N__48786));
    LocalMux I__11358 (
            .O(N__48789),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    Odrv4 I__11357 (
            .O(N__48786),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    InMux I__11356 (
            .O(N__48781),
            .I(bfn_18_22_0_));
    InMux I__11355 (
            .O(N__48778),
            .I(N__48775));
    LocalMux I__11354 (
            .O(N__48775),
            .I(N__48771));
    CascadeMux I__11353 (
            .O(N__48774),
            .I(N__48768));
    Span4Mux_h I__11352 (
            .O(N__48771),
            .I(N__48765));
    InMux I__11351 (
            .O(N__48768),
            .I(N__48761));
    Span4Mux_v I__11350 (
            .O(N__48765),
            .I(N__48758));
    InMux I__11349 (
            .O(N__48764),
            .I(N__48755));
    LocalMux I__11348 (
            .O(N__48761),
            .I(N__48752));
    Odrv4 I__11347 (
            .O(N__48758),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    LocalMux I__11346 (
            .O(N__48755),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    Odrv12 I__11345 (
            .O(N__48752),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    InMux I__11344 (
            .O(N__48745),
            .I(\current_shift_inst.timer_s1.counter_cry_0 ));
    InMux I__11343 (
            .O(N__48742),
            .I(N__48736));
    InMux I__11342 (
            .O(N__48741),
            .I(N__48736));
    LocalMux I__11341 (
            .O(N__48736),
            .I(N__48732));
    InMux I__11340 (
            .O(N__48735),
            .I(N__48729));
    Span4Mux_h I__11339 (
            .O(N__48732),
            .I(N__48726));
    LocalMux I__11338 (
            .O(N__48729),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    Odrv4 I__11337 (
            .O(N__48726),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    InMux I__11336 (
            .O(N__48721),
            .I(\current_shift_inst.timer_s1.counter_cry_1 ));
    InMux I__11335 (
            .O(N__48718),
            .I(N__48711));
    InMux I__11334 (
            .O(N__48717),
            .I(N__48711));
    InMux I__11333 (
            .O(N__48716),
            .I(N__48708));
    LocalMux I__11332 (
            .O(N__48711),
            .I(N__48705));
    LocalMux I__11331 (
            .O(N__48708),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    Odrv12 I__11330 (
            .O(N__48705),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    InMux I__11329 (
            .O(N__48700),
            .I(\current_shift_inst.timer_s1.counter_cry_2 ));
    CascadeMux I__11328 (
            .O(N__48697),
            .I(N__48693));
    CascadeMux I__11327 (
            .O(N__48696),
            .I(N__48690));
    InMux I__11326 (
            .O(N__48693),
            .I(N__48684));
    InMux I__11325 (
            .O(N__48690),
            .I(N__48684));
    InMux I__11324 (
            .O(N__48689),
            .I(N__48681));
    LocalMux I__11323 (
            .O(N__48684),
            .I(N__48678));
    LocalMux I__11322 (
            .O(N__48681),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    Odrv12 I__11321 (
            .O(N__48678),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    InMux I__11320 (
            .O(N__48673),
            .I(\current_shift_inst.timer_s1.counter_cry_3 ));
    CascadeMux I__11319 (
            .O(N__48670),
            .I(N__48667));
    InMux I__11318 (
            .O(N__48667),
            .I(N__48663));
    InMux I__11317 (
            .O(N__48666),
            .I(N__48659));
    LocalMux I__11316 (
            .O(N__48663),
            .I(N__48656));
    InMux I__11315 (
            .O(N__48662),
            .I(N__48653));
    LocalMux I__11314 (
            .O(N__48659),
            .I(N__48650));
    Span4Mux_h I__11313 (
            .O(N__48656),
            .I(N__48647));
    LocalMux I__11312 (
            .O(N__48653),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    Odrv12 I__11311 (
            .O(N__48650),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    Odrv4 I__11310 (
            .O(N__48647),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    InMux I__11309 (
            .O(N__48640),
            .I(\current_shift_inst.timer_s1.counter_cry_4 ));
    InMux I__11308 (
            .O(N__48637),
            .I(N__48630));
    InMux I__11307 (
            .O(N__48636),
            .I(N__48630));
    InMux I__11306 (
            .O(N__48635),
            .I(N__48627));
    LocalMux I__11305 (
            .O(N__48630),
            .I(N__48624));
    LocalMux I__11304 (
            .O(N__48627),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    Odrv12 I__11303 (
            .O(N__48624),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    InMux I__11302 (
            .O(N__48619),
            .I(\current_shift_inst.timer_s1.counter_cry_5 ));
    CascadeMux I__11301 (
            .O(N__48616),
            .I(N__48612));
    CascadeMux I__11300 (
            .O(N__48615),
            .I(N__48609));
    InMux I__11299 (
            .O(N__48612),
            .I(N__48604));
    InMux I__11298 (
            .O(N__48609),
            .I(N__48604));
    LocalMux I__11297 (
            .O(N__48604),
            .I(N__48600));
    InMux I__11296 (
            .O(N__48603),
            .I(N__48597));
    Span4Mux_v I__11295 (
            .O(N__48600),
            .I(N__48594));
    LocalMux I__11294 (
            .O(N__48597),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    Odrv4 I__11293 (
            .O(N__48594),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    InMux I__11292 (
            .O(N__48589),
            .I(\current_shift_inst.timer_s1.counter_cry_6 ));
    CascadeMux I__11291 (
            .O(N__48586),
            .I(N__48583));
    InMux I__11290 (
            .O(N__48583),
            .I(N__48580));
    LocalMux I__11289 (
            .O(N__48580),
            .I(N__48575));
    InMux I__11288 (
            .O(N__48579),
            .I(N__48572));
    InMux I__11287 (
            .O(N__48578),
            .I(N__48569));
    Span4Mux_v I__11286 (
            .O(N__48575),
            .I(N__48566));
    LocalMux I__11285 (
            .O(N__48572),
            .I(N__48563));
    LocalMux I__11284 (
            .O(N__48569),
            .I(N__48560));
    Span4Mux_h I__11283 (
            .O(N__48566),
            .I(N__48556));
    Span4Mux_v I__11282 (
            .O(N__48563),
            .I(N__48551));
    Span4Mux_v I__11281 (
            .O(N__48560),
            .I(N__48551));
    InMux I__11280 (
            .O(N__48559),
            .I(N__48548));
    Odrv4 I__11279 (
            .O(N__48556),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    Odrv4 I__11278 (
            .O(N__48551),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    LocalMux I__11277 (
            .O(N__48548),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    InMux I__11276 (
            .O(N__48541),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ));
    InMux I__11275 (
            .O(N__48538),
            .I(N__48534));
    InMux I__11274 (
            .O(N__48537),
            .I(N__48531));
    LocalMux I__11273 (
            .O(N__48534),
            .I(N__48524));
    LocalMux I__11272 (
            .O(N__48531),
            .I(N__48524));
    InMux I__11271 (
            .O(N__48530),
            .I(N__48521));
    InMux I__11270 (
            .O(N__48529),
            .I(N__48518));
    Span4Mux_v I__11269 (
            .O(N__48524),
            .I(N__48515));
    LocalMux I__11268 (
            .O(N__48521),
            .I(N__48512));
    LocalMux I__11267 (
            .O(N__48518),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    Odrv4 I__11266 (
            .O(N__48515),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    Odrv4 I__11265 (
            .O(N__48512),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    InMux I__11264 (
            .O(N__48505),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ));
    CascadeMux I__11263 (
            .O(N__48502),
            .I(N__48499));
    InMux I__11262 (
            .O(N__48499),
            .I(N__48492));
    InMux I__11261 (
            .O(N__48498),
            .I(N__48492));
    InMux I__11260 (
            .O(N__48497),
            .I(N__48489));
    LocalMux I__11259 (
            .O(N__48492),
            .I(N__48486));
    LocalMux I__11258 (
            .O(N__48489),
            .I(N__48482));
    Span4Mux_h I__11257 (
            .O(N__48486),
            .I(N__48479));
    InMux I__11256 (
            .O(N__48485),
            .I(N__48476));
    Odrv12 I__11255 (
            .O(N__48482),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    Odrv4 I__11254 (
            .O(N__48479),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    LocalMux I__11253 (
            .O(N__48476),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    InMux I__11252 (
            .O(N__48469),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ));
    InMux I__11251 (
            .O(N__48466),
            .I(N__48462));
    InMux I__11250 (
            .O(N__48465),
            .I(N__48459));
    LocalMux I__11249 (
            .O(N__48462),
            .I(N__48456));
    LocalMux I__11248 (
            .O(N__48459),
            .I(N__48452));
    Span4Mux_h I__11247 (
            .O(N__48456),
            .I(N__48448));
    InMux I__11246 (
            .O(N__48455),
            .I(N__48445));
    Span4Mux_h I__11245 (
            .O(N__48452),
            .I(N__48442));
    InMux I__11244 (
            .O(N__48451),
            .I(N__48439));
    Odrv4 I__11243 (
            .O(N__48448),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    LocalMux I__11242 (
            .O(N__48445),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    Odrv4 I__11241 (
            .O(N__48442),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    LocalMux I__11240 (
            .O(N__48439),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    InMux I__11239 (
            .O(N__48430),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ));
    InMux I__11238 (
            .O(N__48427),
            .I(N__48423));
    InMux I__11237 (
            .O(N__48426),
            .I(N__48420));
    LocalMux I__11236 (
            .O(N__48423),
            .I(N__48416));
    LocalMux I__11235 (
            .O(N__48420),
            .I(N__48413));
    InMux I__11234 (
            .O(N__48419),
            .I(N__48410));
    Span4Mux_v I__11233 (
            .O(N__48416),
            .I(N__48407));
    Span4Mux_h I__11232 (
            .O(N__48413),
            .I(N__48404));
    LocalMux I__11231 (
            .O(N__48410),
            .I(N__48400));
    Span4Mux_h I__11230 (
            .O(N__48407),
            .I(N__48395));
    Span4Mux_v I__11229 (
            .O(N__48404),
            .I(N__48395));
    InMux I__11228 (
            .O(N__48403),
            .I(N__48392));
    Odrv4 I__11227 (
            .O(N__48400),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    Odrv4 I__11226 (
            .O(N__48395),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    LocalMux I__11225 (
            .O(N__48392),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    InMux I__11224 (
            .O(N__48385),
            .I(bfn_18_21_0_));
    InMux I__11223 (
            .O(N__48382),
            .I(N__48378));
    InMux I__11222 (
            .O(N__48381),
            .I(N__48375));
    LocalMux I__11221 (
            .O(N__48378),
            .I(N__48370));
    LocalMux I__11220 (
            .O(N__48375),
            .I(N__48367));
    InMux I__11219 (
            .O(N__48374),
            .I(N__48364));
    InMux I__11218 (
            .O(N__48373),
            .I(N__48361));
    Span4Mux_h I__11217 (
            .O(N__48370),
            .I(N__48356));
    Span4Mux_h I__11216 (
            .O(N__48367),
            .I(N__48356));
    LocalMux I__11215 (
            .O(N__48364),
            .I(N__48353));
    LocalMux I__11214 (
            .O(N__48361),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    Odrv4 I__11213 (
            .O(N__48356),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    Odrv12 I__11212 (
            .O(N__48353),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    InMux I__11211 (
            .O(N__48346),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ));
    InMux I__11210 (
            .O(N__48343),
            .I(N__48338));
    InMux I__11209 (
            .O(N__48342),
            .I(N__48333));
    InMux I__11208 (
            .O(N__48341),
            .I(N__48333));
    LocalMux I__11207 (
            .O(N__48338),
            .I(N__48330));
    LocalMux I__11206 (
            .O(N__48333),
            .I(N__48327));
    Span4Mux_h I__11205 (
            .O(N__48330),
            .I(N__48323));
    Span4Mux_v I__11204 (
            .O(N__48327),
            .I(N__48320));
    InMux I__11203 (
            .O(N__48326),
            .I(N__48317));
    Odrv4 I__11202 (
            .O(N__48323),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    Odrv4 I__11201 (
            .O(N__48320),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    LocalMux I__11200 (
            .O(N__48317),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    InMux I__11199 (
            .O(N__48310),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ));
    InMux I__11198 (
            .O(N__48307),
            .I(N__48304));
    LocalMux I__11197 (
            .O(N__48304),
            .I(N__48299));
    InMux I__11196 (
            .O(N__48303),
            .I(N__48296));
    InMux I__11195 (
            .O(N__48302),
            .I(N__48293));
    Span4Mux_v I__11194 (
            .O(N__48299),
            .I(N__48288));
    LocalMux I__11193 (
            .O(N__48296),
            .I(N__48288));
    LocalMux I__11192 (
            .O(N__48293),
            .I(N__48285));
    Span4Mux_h I__11191 (
            .O(N__48288),
            .I(N__48279));
    Span4Mux_v I__11190 (
            .O(N__48285),
            .I(N__48279));
    InMux I__11189 (
            .O(N__48284),
            .I(N__48276));
    Odrv4 I__11188 (
            .O(N__48279),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    LocalMux I__11187 (
            .O(N__48276),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    InMux I__11186 (
            .O(N__48271),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ));
    CEMux I__11185 (
            .O(N__48268),
            .I(N__48244));
    CEMux I__11184 (
            .O(N__48267),
            .I(N__48244));
    CEMux I__11183 (
            .O(N__48266),
            .I(N__48244));
    CEMux I__11182 (
            .O(N__48265),
            .I(N__48244));
    CEMux I__11181 (
            .O(N__48264),
            .I(N__48244));
    CEMux I__11180 (
            .O(N__48263),
            .I(N__48244));
    CEMux I__11179 (
            .O(N__48262),
            .I(N__48244));
    CEMux I__11178 (
            .O(N__48261),
            .I(N__48244));
    GlobalMux I__11177 (
            .O(N__48244),
            .I(N__48241));
    gio2CtrlBuf I__11176 (
            .O(N__48241),
            .I(\current_shift_inst.timer_s1.N_180_i_g ));
    InMux I__11175 (
            .O(N__48238),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ));
    InMux I__11174 (
            .O(N__48235),
            .I(N__48230));
    InMux I__11173 (
            .O(N__48234),
            .I(N__48227));
    InMux I__11172 (
            .O(N__48233),
            .I(N__48224));
    LocalMux I__11171 (
            .O(N__48230),
            .I(N__48221));
    LocalMux I__11170 (
            .O(N__48227),
            .I(N__48217));
    LocalMux I__11169 (
            .O(N__48224),
            .I(N__48214));
    Span4Mux_v I__11168 (
            .O(N__48221),
            .I(N__48211));
    InMux I__11167 (
            .O(N__48220),
            .I(N__48208));
    Span4Mux_v I__11166 (
            .O(N__48217),
            .I(N__48203));
    Span4Mux_v I__11165 (
            .O(N__48214),
            .I(N__48203));
    Span4Mux_h I__11164 (
            .O(N__48211),
            .I(N__48198));
    LocalMux I__11163 (
            .O(N__48208),
            .I(N__48198));
    Odrv4 I__11162 (
            .O(N__48203),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    Odrv4 I__11161 (
            .O(N__48198),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    InMux I__11160 (
            .O(N__48193),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ));
    InMux I__11159 (
            .O(N__48190),
            .I(N__48185));
    InMux I__11158 (
            .O(N__48189),
            .I(N__48182));
    InMux I__11157 (
            .O(N__48188),
            .I(N__48179));
    LocalMux I__11156 (
            .O(N__48185),
            .I(N__48176));
    LocalMux I__11155 (
            .O(N__48182),
            .I(N__48172));
    LocalMux I__11154 (
            .O(N__48179),
            .I(N__48169));
    Span4Mux_v I__11153 (
            .O(N__48176),
            .I(N__48166));
    InMux I__11152 (
            .O(N__48175),
            .I(N__48163));
    Span4Mux_v I__11151 (
            .O(N__48172),
            .I(N__48158));
    Span4Mux_v I__11150 (
            .O(N__48169),
            .I(N__48158));
    Span4Mux_h I__11149 (
            .O(N__48166),
            .I(N__48153));
    LocalMux I__11148 (
            .O(N__48163),
            .I(N__48153));
    Odrv4 I__11147 (
            .O(N__48158),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    Odrv4 I__11146 (
            .O(N__48153),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    InMux I__11145 (
            .O(N__48148),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ));
    InMux I__11144 (
            .O(N__48145),
            .I(N__48140));
    InMux I__11143 (
            .O(N__48144),
            .I(N__48137));
    InMux I__11142 (
            .O(N__48143),
            .I(N__48134));
    LocalMux I__11141 (
            .O(N__48140),
            .I(N__48130));
    LocalMux I__11140 (
            .O(N__48137),
            .I(N__48127));
    LocalMux I__11139 (
            .O(N__48134),
            .I(N__48124));
    InMux I__11138 (
            .O(N__48133),
            .I(N__48121));
    Span4Mux_h I__11137 (
            .O(N__48130),
            .I(N__48118));
    Span4Mux_h I__11136 (
            .O(N__48127),
            .I(N__48115));
    Span4Mux_v I__11135 (
            .O(N__48124),
            .I(N__48110));
    LocalMux I__11134 (
            .O(N__48121),
            .I(N__48110));
    Odrv4 I__11133 (
            .O(N__48118),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    Odrv4 I__11132 (
            .O(N__48115),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    Odrv4 I__11131 (
            .O(N__48110),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    InMux I__11130 (
            .O(N__48103),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ));
    InMux I__11129 (
            .O(N__48100),
            .I(N__48096));
    InMux I__11128 (
            .O(N__48099),
            .I(N__48093));
    LocalMux I__11127 (
            .O(N__48096),
            .I(N__48090));
    LocalMux I__11126 (
            .O(N__48093),
            .I(N__48087));
    Span4Mux_h I__11125 (
            .O(N__48090),
            .I(N__48082));
    Span4Mux_h I__11124 (
            .O(N__48087),
            .I(N__48079));
    InMux I__11123 (
            .O(N__48086),
            .I(N__48074));
    InMux I__11122 (
            .O(N__48085),
            .I(N__48074));
    Odrv4 I__11121 (
            .O(N__48082),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    Odrv4 I__11120 (
            .O(N__48079),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    LocalMux I__11119 (
            .O(N__48074),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    InMux I__11118 (
            .O(N__48067),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__11117 (
            .O(N__48064),
            .I(N__48061));
    InMux I__11116 (
            .O(N__48061),
            .I(N__48058));
    LocalMux I__11115 (
            .O(N__48058),
            .I(N__48053));
    InMux I__11114 (
            .O(N__48057),
            .I(N__48050));
    InMux I__11113 (
            .O(N__48056),
            .I(N__48046));
    Span4Mux_v I__11112 (
            .O(N__48053),
            .I(N__48043));
    LocalMux I__11111 (
            .O(N__48050),
            .I(N__48040));
    InMux I__11110 (
            .O(N__48049),
            .I(N__48037));
    LocalMux I__11109 (
            .O(N__48046),
            .I(N__48034));
    Span4Mux_h I__11108 (
            .O(N__48043),
            .I(N__48027));
    Span4Mux_v I__11107 (
            .O(N__48040),
            .I(N__48027));
    LocalMux I__11106 (
            .O(N__48037),
            .I(N__48027));
    Odrv4 I__11105 (
            .O(N__48034),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    Odrv4 I__11104 (
            .O(N__48027),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    InMux I__11103 (
            .O(N__48022),
            .I(bfn_18_20_0_));
    InMux I__11102 (
            .O(N__48019),
            .I(N__48012));
    InMux I__11101 (
            .O(N__48018),
            .I(N__48012));
    InMux I__11100 (
            .O(N__48017),
            .I(N__48009));
    LocalMux I__11099 (
            .O(N__48012),
            .I(N__48006));
    LocalMux I__11098 (
            .O(N__48009),
            .I(N__48002));
    Span4Mux_h I__11097 (
            .O(N__48006),
            .I(N__47999));
    InMux I__11096 (
            .O(N__48005),
            .I(N__47996));
    Odrv4 I__11095 (
            .O(N__48002),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    Odrv4 I__11094 (
            .O(N__47999),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    LocalMux I__11093 (
            .O(N__47996),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    InMux I__11092 (
            .O(N__47989),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ));
    CascadeMux I__11091 (
            .O(N__47986),
            .I(N__47982));
    InMux I__11090 (
            .O(N__47985),
            .I(N__47978));
    InMux I__11089 (
            .O(N__47982),
            .I(N__47973));
    InMux I__11088 (
            .O(N__47981),
            .I(N__47973));
    LocalMux I__11087 (
            .O(N__47978),
            .I(N__47968));
    LocalMux I__11086 (
            .O(N__47973),
            .I(N__47968));
    Span4Mux_v I__11085 (
            .O(N__47968),
            .I(N__47964));
    InMux I__11084 (
            .O(N__47967),
            .I(N__47961));
    Odrv4 I__11083 (
            .O(N__47964),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    LocalMux I__11082 (
            .O(N__47961),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    InMux I__11081 (
            .O(N__47956),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ));
    CascadeMux I__11080 (
            .O(N__47953),
            .I(N__47949));
    InMux I__11079 (
            .O(N__47952),
            .I(N__47945));
    InMux I__11078 (
            .O(N__47949),
            .I(N__47942));
    InMux I__11077 (
            .O(N__47948),
            .I(N__47939));
    LocalMux I__11076 (
            .O(N__47945),
            .I(N__47936));
    LocalMux I__11075 (
            .O(N__47942),
            .I(N__47933));
    LocalMux I__11074 (
            .O(N__47939),
            .I(N__47930));
    Span4Mux_v I__11073 (
            .O(N__47936),
            .I(N__47927));
    Span4Mux_h I__11072 (
            .O(N__47933),
            .I(N__47923));
    Span4Mux_v I__11071 (
            .O(N__47930),
            .I(N__47918));
    Span4Mux_h I__11070 (
            .O(N__47927),
            .I(N__47918));
    InMux I__11069 (
            .O(N__47926),
            .I(N__47915));
    Odrv4 I__11068 (
            .O(N__47923),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    Odrv4 I__11067 (
            .O(N__47918),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    LocalMux I__11066 (
            .O(N__47915),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    InMux I__11065 (
            .O(N__47908),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ));
    InMux I__11064 (
            .O(N__47905),
            .I(N__47902));
    LocalMux I__11063 (
            .O(N__47902),
            .I(N__47897));
    InMux I__11062 (
            .O(N__47901),
            .I(N__47894));
    InMux I__11061 (
            .O(N__47900),
            .I(N__47890));
    Span4Mux_v I__11060 (
            .O(N__47897),
            .I(N__47885));
    LocalMux I__11059 (
            .O(N__47894),
            .I(N__47885));
    InMux I__11058 (
            .O(N__47893),
            .I(N__47882));
    LocalMux I__11057 (
            .O(N__47890),
            .I(N__47879));
    Span4Mux_h I__11056 (
            .O(N__47885),
            .I(N__47876));
    LocalMux I__11055 (
            .O(N__47882),
            .I(N__47873));
    Odrv4 I__11054 (
            .O(N__47879),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    Odrv4 I__11053 (
            .O(N__47876),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    Odrv4 I__11052 (
            .O(N__47873),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    InMux I__11051 (
            .O(N__47866),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ));
    InMux I__11050 (
            .O(N__47863),
            .I(N__47855));
    InMux I__11049 (
            .O(N__47862),
            .I(N__47855));
    InMux I__11048 (
            .O(N__47861),
            .I(N__47852));
    InMux I__11047 (
            .O(N__47860),
            .I(N__47849));
    LocalMux I__11046 (
            .O(N__47855),
            .I(N__47846));
    LocalMux I__11045 (
            .O(N__47852),
            .I(N__47841));
    LocalMux I__11044 (
            .O(N__47849),
            .I(N__47841));
    Odrv12 I__11043 (
            .O(N__47846),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    Odrv4 I__11042 (
            .O(N__47841),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    InMux I__11041 (
            .O(N__47836),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ));
    InMux I__11040 (
            .O(N__47833),
            .I(N__47830));
    LocalMux I__11039 (
            .O(N__47830),
            .I(N__47826));
    InMux I__11038 (
            .O(N__47829),
            .I(N__47823));
    Span4Mux_v I__11037 (
            .O(N__47826),
            .I(N__47816));
    LocalMux I__11036 (
            .O(N__47823),
            .I(N__47816));
    InMux I__11035 (
            .O(N__47822),
            .I(N__47811));
    InMux I__11034 (
            .O(N__47821),
            .I(N__47811));
    Span4Mux_h I__11033 (
            .O(N__47816),
            .I(N__47806));
    LocalMux I__11032 (
            .O(N__47811),
            .I(N__47806));
    Odrv4 I__11031 (
            .O(N__47806),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    InMux I__11030 (
            .O(N__47803),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ));
    InMux I__11029 (
            .O(N__47800),
            .I(N__47797));
    LocalMux I__11028 (
            .O(N__47797),
            .I(N__47792));
    InMux I__11027 (
            .O(N__47796),
            .I(N__47789));
    InMux I__11026 (
            .O(N__47795),
            .I(N__47786));
    Span4Mux_v I__11025 (
            .O(N__47792),
            .I(N__47780));
    LocalMux I__11024 (
            .O(N__47789),
            .I(N__47780));
    LocalMux I__11023 (
            .O(N__47786),
            .I(N__47777));
    InMux I__11022 (
            .O(N__47785),
            .I(N__47774));
    Span4Mux_h I__11021 (
            .O(N__47780),
            .I(N__47771));
    Span4Mux_h I__11020 (
            .O(N__47777),
            .I(N__47768));
    LocalMux I__11019 (
            .O(N__47774),
            .I(N__47765));
    Odrv4 I__11018 (
            .O(N__47771),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    Odrv4 I__11017 (
            .O(N__47768),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    Odrv12 I__11016 (
            .O(N__47765),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    InMux I__11015 (
            .O(N__47758),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ));
    InMux I__11014 (
            .O(N__47755),
            .I(N__47752));
    LocalMux I__11013 (
            .O(N__47752),
            .I(N__47747));
    InMux I__11012 (
            .O(N__47751),
            .I(N__47744));
    InMux I__11011 (
            .O(N__47750),
            .I(N__47741));
    Span4Mux_h I__11010 (
            .O(N__47747),
            .I(N__47736));
    LocalMux I__11009 (
            .O(N__47744),
            .I(N__47736));
    LocalMux I__11008 (
            .O(N__47741),
            .I(N__47733));
    Span4Mux_h I__11007 (
            .O(N__47736),
            .I(N__47729));
    Span4Mux_h I__11006 (
            .O(N__47733),
            .I(N__47726));
    InMux I__11005 (
            .O(N__47732),
            .I(N__47723));
    Odrv4 I__11004 (
            .O(N__47729),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    Odrv4 I__11003 (
            .O(N__47726),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    LocalMux I__11002 (
            .O(N__47723),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    InMux I__11001 (
            .O(N__47716),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ));
    InMux I__11000 (
            .O(N__47713),
            .I(N__47710));
    LocalMux I__10999 (
            .O(N__47710),
            .I(N__47705));
    InMux I__10998 (
            .O(N__47709),
            .I(N__47702));
    InMux I__10997 (
            .O(N__47708),
            .I(N__47698));
    Span4Mux_h I__10996 (
            .O(N__47705),
            .I(N__47693));
    LocalMux I__10995 (
            .O(N__47702),
            .I(N__47693));
    InMux I__10994 (
            .O(N__47701),
            .I(N__47690));
    LocalMux I__10993 (
            .O(N__47698),
            .I(N__47687));
    Span4Mux_h I__10992 (
            .O(N__47693),
            .I(N__47682));
    LocalMux I__10991 (
            .O(N__47690),
            .I(N__47682));
    Odrv4 I__10990 (
            .O(N__47687),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    Odrv4 I__10989 (
            .O(N__47682),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    InMux I__10988 (
            .O(N__47677),
            .I(bfn_18_19_0_));
    InMux I__10987 (
            .O(N__47674),
            .I(N__47669));
    InMux I__10986 (
            .O(N__47673),
            .I(N__47666));
    InMux I__10985 (
            .O(N__47672),
            .I(N__47662));
    LocalMux I__10984 (
            .O(N__47669),
            .I(N__47659));
    LocalMux I__10983 (
            .O(N__47666),
            .I(N__47656));
    InMux I__10982 (
            .O(N__47665),
            .I(N__47653));
    LocalMux I__10981 (
            .O(N__47662),
            .I(N__47650));
    Span4Mux_v I__10980 (
            .O(N__47659),
            .I(N__47643));
    Span4Mux_h I__10979 (
            .O(N__47656),
            .I(N__47643));
    LocalMux I__10978 (
            .O(N__47653),
            .I(N__47643));
    Odrv4 I__10977 (
            .O(N__47650),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    Odrv4 I__10976 (
            .O(N__47643),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    InMux I__10975 (
            .O(N__47638),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__10974 (
            .O(N__47635),
            .I(N__47632));
    InMux I__10973 (
            .O(N__47632),
            .I(N__47627));
    InMux I__10972 (
            .O(N__47631),
            .I(N__47624));
    InMux I__10971 (
            .O(N__47630),
            .I(N__47621));
    LocalMux I__10970 (
            .O(N__47627),
            .I(N__47617));
    LocalMux I__10969 (
            .O(N__47624),
            .I(N__47614));
    LocalMux I__10968 (
            .O(N__47621),
            .I(N__47611));
    InMux I__10967 (
            .O(N__47620),
            .I(N__47608));
    Span4Mux_h I__10966 (
            .O(N__47617),
            .I(N__47603));
    Span4Mux_v I__10965 (
            .O(N__47614),
            .I(N__47603));
    Span4Mux_h I__10964 (
            .O(N__47611),
            .I(N__47598));
    LocalMux I__10963 (
            .O(N__47608),
            .I(N__47598));
    Odrv4 I__10962 (
            .O(N__47603),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    Odrv4 I__10961 (
            .O(N__47598),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    InMux I__10960 (
            .O(N__47593),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ));
    InMux I__10959 (
            .O(N__47590),
            .I(N__47587));
    LocalMux I__10958 (
            .O(N__47587),
            .I(N__47582));
    InMux I__10957 (
            .O(N__47586),
            .I(N__47579));
    InMux I__10956 (
            .O(N__47585),
            .I(N__47575));
    Span4Mux_v I__10955 (
            .O(N__47582),
            .I(N__47570));
    LocalMux I__10954 (
            .O(N__47579),
            .I(N__47570));
    InMux I__10953 (
            .O(N__47578),
            .I(N__47567));
    LocalMux I__10952 (
            .O(N__47575),
            .I(N__47564));
    Span4Mux_h I__10951 (
            .O(N__47570),
            .I(N__47559));
    LocalMux I__10950 (
            .O(N__47567),
            .I(N__47559));
    Odrv4 I__10949 (
            .O(N__47564),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    Odrv4 I__10948 (
            .O(N__47559),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    InMux I__10947 (
            .O(N__47554),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ));
    InMux I__10946 (
            .O(N__47551),
            .I(N__47548));
    LocalMux I__10945 (
            .O(N__47548),
            .I(\current_shift_inst.un4_control_input_1_axb_14 ));
    InMux I__10944 (
            .O(N__47545),
            .I(N__47542));
    LocalMux I__10943 (
            .O(N__47542),
            .I(\current_shift_inst.un4_control_input_1_axb_16 ));
    InMux I__10942 (
            .O(N__47539),
            .I(N__47536));
    LocalMux I__10941 (
            .O(N__47536),
            .I(\current_shift_inst.un4_control_input_1_axb_23 ));
    InMux I__10940 (
            .O(N__47533),
            .I(N__47530));
    LocalMux I__10939 (
            .O(N__47530),
            .I(\current_shift_inst.un4_control_input_1_axb_10 ));
    InMux I__10938 (
            .O(N__47527),
            .I(N__47524));
    LocalMux I__10937 (
            .O(N__47524),
            .I(\current_shift_inst.un4_control_input_1_axb_12 ));
    CascadeMux I__10936 (
            .O(N__47521),
            .I(N__47518));
    InMux I__10935 (
            .O(N__47518),
            .I(N__47512));
    InMux I__10934 (
            .O(N__47517),
            .I(N__47512));
    LocalMux I__10933 (
            .O(N__47512),
            .I(N__47509));
    Span4Mux_v I__10932 (
            .O(N__47509),
            .I(N__47504));
    InMux I__10931 (
            .O(N__47508),
            .I(N__47501));
    InMux I__10930 (
            .O(N__47507),
            .I(N__47498));
    Span4Mux_h I__10929 (
            .O(N__47504),
            .I(N__47495));
    LocalMux I__10928 (
            .O(N__47501),
            .I(N__47492));
    LocalMux I__10927 (
            .O(N__47498),
            .I(N__47489));
    Odrv4 I__10926 (
            .O(N__47495),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    Odrv4 I__10925 (
            .O(N__47492),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    Odrv4 I__10924 (
            .O(N__47489),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    CascadeMux I__10923 (
            .O(N__47482),
            .I(N__47479));
    InMux I__10922 (
            .O(N__47479),
            .I(N__47470));
    InMux I__10921 (
            .O(N__47478),
            .I(N__47470));
    InMux I__10920 (
            .O(N__47477),
            .I(N__47470));
    LocalMux I__10919 (
            .O(N__47470),
            .I(N__47466));
    InMux I__10918 (
            .O(N__47469),
            .I(N__47463));
    Span4Mux_h I__10917 (
            .O(N__47466),
            .I(N__47460));
    LocalMux I__10916 (
            .O(N__47463),
            .I(N__47457));
    Odrv4 I__10915 (
            .O(N__47460),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    Odrv4 I__10914 (
            .O(N__47457),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    InMux I__10913 (
            .O(N__47452),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ));
    InMux I__10912 (
            .O(N__47449),
            .I(N__47444));
    InMux I__10911 (
            .O(N__47448),
            .I(N__47441));
    InMux I__10910 (
            .O(N__47447),
            .I(N__47438));
    LocalMux I__10909 (
            .O(N__47444),
            .I(N__47434));
    LocalMux I__10908 (
            .O(N__47441),
            .I(N__47431));
    LocalMux I__10907 (
            .O(N__47438),
            .I(N__47428));
    InMux I__10906 (
            .O(N__47437),
            .I(N__47425));
    Span4Mux_h I__10905 (
            .O(N__47434),
            .I(N__47422));
    Span4Mux_v I__10904 (
            .O(N__47431),
            .I(N__47415));
    Span4Mux_h I__10903 (
            .O(N__47428),
            .I(N__47415));
    LocalMux I__10902 (
            .O(N__47425),
            .I(N__47415));
    Odrv4 I__10901 (
            .O(N__47422),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    Odrv4 I__10900 (
            .O(N__47415),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    InMux I__10899 (
            .O(N__47410),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ));
    InMux I__10898 (
            .O(N__47407),
            .I(N__47404));
    LocalMux I__10897 (
            .O(N__47404),
            .I(N__47401));
    Span4Mux_h I__10896 (
            .O(N__47401),
            .I(N__47396));
    InMux I__10895 (
            .O(N__47400),
            .I(N__47393));
    InMux I__10894 (
            .O(N__47399),
            .I(N__47390));
    Odrv4 I__10893 (
            .O(N__47396),
            .I(\current_shift_inst.un4_control_input1_8 ));
    LocalMux I__10892 (
            .O(N__47393),
            .I(\current_shift_inst.un4_control_input1_8 ));
    LocalMux I__10891 (
            .O(N__47390),
            .I(\current_shift_inst.un4_control_input1_8 ));
    InMux I__10890 (
            .O(N__47383),
            .I(N__47380));
    LocalMux I__10889 (
            .O(N__47380),
            .I(N__47377));
    Span4Mux_v I__10888 (
            .O(N__47377),
            .I(N__47374));
    Odrv4 I__10887 (
            .O(N__47374),
            .I(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_8 ));
    CascadeMux I__10886 (
            .O(N__47371),
            .I(N__47368));
    InMux I__10885 (
            .O(N__47368),
            .I(N__47365));
    LocalMux I__10884 (
            .O(N__47365),
            .I(\current_shift_inst.un4_control_input_1_axb_15 ));
    InMux I__10883 (
            .O(N__47362),
            .I(N__47359));
    LocalMux I__10882 (
            .O(N__47359),
            .I(\current_shift_inst.un4_control_input_1_axb_7 ));
    InMux I__10881 (
            .O(N__47356),
            .I(N__47353));
    LocalMux I__10880 (
            .O(N__47353),
            .I(\current_shift_inst.un4_control_input_1_axb_2 ));
    InMux I__10879 (
            .O(N__47350),
            .I(N__47347));
    LocalMux I__10878 (
            .O(N__47347),
            .I(\current_shift_inst.un4_control_input_1_axb_6 ));
    InMux I__10877 (
            .O(N__47344),
            .I(N__47341));
    LocalMux I__10876 (
            .O(N__47341),
            .I(\current_shift_inst.un4_control_input_1_axb_4 ));
    InMux I__10875 (
            .O(N__47338),
            .I(N__47335));
    LocalMux I__10874 (
            .O(N__47335),
            .I(\current_shift_inst.un4_control_input_1_axb_5 ));
    InMux I__10873 (
            .O(N__47332),
            .I(N__47329));
    LocalMux I__10872 (
            .O(N__47329),
            .I(\current_shift_inst.un4_control_input_1_axb_11 ));
    InMux I__10871 (
            .O(N__47326),
            .I(N__47323));
    LocalMux I__10870 (
            .O(N__47323),
            .I(\current_shift_inst.un4_control_input_1_axb_13 ));
    InMux I__10869 (
            .O(N__47320),
            .I(N__47317));
    LocalMux I__10868 (
            .O(N__47317),
            .I(\current_shift_inst.un4_control_input_1_axb_9 ));
    InMux I__10867 (
            .O(N__47314),
            .I(N__47308));
    InMux I__10866 (
            .O(N__47313),
            .I(N__47308));
    LocalMux I__10865 (
            .O(N__47308),
            .I(N__47305));
    Span4Mux_h I__10864 (
            .O(N__47305),
            .I(N__47302));
    Span4Mux_h I__10863 (
            .O(N__47302),
            .I(N__47297));
    InMux I__10862 (
            .O(N__47301),
            .I(N__47292));
    InMux I__10861 (
            .O(N__47300),
            .I(N__47292));
    Odrv4 I__10860 (
            .O(N__47297),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    LocalMux I__10859 (
            .O(N__47292),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    InMux I__10858 (
            .O(N__47287),
            .I(N__47284));
    LocalMux I__10857 (
            .O(N__47284),
            .I(\current_shift_inst.un4_control_input_1_axb_8 ));
    InMux I__10856 (
            .O(N__47281),
            .I(N__47254));
    InMux I__10855 (
            .O(N__47280),
            .I(N__47254));
    InMux I__10854 (
            .O(N__47279),
            .I(N__47254));
    InMux I__10853 (
            .O(N__47278),
            .I(N__47254));
    InMux I__10852 (
            .O(N__47277),
            .I(N__47254));
    InMux I__10851 (
            .O(N__47276),
            .I(N__47251));
    InMux I__10850 (
            .O(N__47275),
            .I(N__47246));
    InMux I__10849 (
            .O(N__47274),
            .I(N__47246));
    InMux I__10848 (
            .O(N__47273),
            .I(N__47241));
    InMux I__10847 (
            .O(N__47272),
            .I(N__47241));
    InMux I__10846 (
            .O(N__47271),
            .I(N__47234));
    InMux I__10845 (
            .O(N__47270),
            .I(N__47234));
    InMux I__10844 (
            .O(N__47269),
            .I(N__47234));
    InMux I__10843 (
            .O(N__47268),
            .I(N__47227));
    InMux I__10842 (
            .O(N__47267),
            .I(N__47227));
    InMux I__10841 (
            .O(N__47266),
            .I(N__47227));
    InMux I__10840 (
            .O(N__47265),
            .I(N__47220));
    LocalMux I__10839 (
            .O(N__47254),
            .I(N__47216));
    LocalMux I__10838 (
            .O(N__47251),
            .I(N__47212));
    LocalMux I__10837 (
            .O(N__47246),
            .I(N__47203));
    LocalMux I__10836 (
            .O(N__47241),
            .I(N__47203));
    LocalMux I__10835 (
            .O(N__47234),
            .I(N__47203));
    LocalMux I__10834 (
            .O(N__47227),
            .I(N__47203));
    InMux I__10833 (
            .O(N__47226),
            .I(N__47198));
    InMux I__10832 (
            .O(N__47225),
            .I(N__47198));
    InMux I__10831 (
            .O(N__47224),
            .I(N__47193));
    InMux I__10830 (
            .O(N__47223),
            .I(N__47193));
    LocalMux I__10829 (
            .O(N__47220),
            .I(N__47189));
    InMux I__10828 (
            .O(N__47219),
            .I(N__47185));
    Span4Mux_h I__10827 (
            .O(N__47216),
            .I(N__47182));
    InMux I__10826 (
            .O(N__47215),
            .I(N__47179));
    Span4Mux_v I__10825 (
            .O(N__47212),
            .I(N__47170));
    Span4Mux_v I__10824 (
            .O(N__47203),
            .I(N__47170));
    LocalMux I__10823 (
            .O(N__47198),
            .I(N__47170));
    LocalMux I__10822 (
            .O(N__47193),
            .I(N__47170));
    InMux I__10821 (
            .O(N__47192),
            .I(N__47167));
    Span4Mux_h I__10820 (
            .O(N__47189),
            .I(N__47164));
    InMux I__10819 (
            .O(N__47188),
            .I(N__47161));
    LocalMux I__10818 (
            .O(N__47185),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__10817 (
            .O(N__47182),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__10816 (
            .O(N__47179),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__10815 (
            .O(N__47170),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__10814 (
            .O(N__47167),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__10813 (
            .O(N__47164),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__10812 (
            .O(N__47161),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    InMux I__10811 (
            .O(N__47146),
            .I(N__47140));
    InMux I__10810 (
            .O(N__47145),
            .I(N__47140));
    LocalMux I__10809 (
            .O(N__47140),
            .I(N__47137));
    Span12Mux_v I__10808 (
            .O(N__47137),
            .I(N__47133));
    InMux I__10807 (
            .O(N__47136),
            .I(N__47130));
    Odrv12 I__10806 (
            .O(N__47133),
            .I(\current_shift_inst.un4_control_input1_3 ));
    LocalMux I__10805 (
            .O(N__47130),
            .I(\current_shift_inst.un4_control_input1_3 ));
    InMux I__10804 (
            .O(N__47125),
            .I(N__47122));
    LocalMux I__10803 (
            .O(N__47122),
            .I(N__47119));
    Odrv4 I__10802 (
            .O(N__47119),
            .I(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ));
    InMux I__10801 (
            .O(N__47116),
            .I(N__47113));
    LocalMux I__10800 (
            .O(N__47113),
            .I(N__47108));
    InMux I__10799 (
            .O(N__47112),
            .I(N__47105));
    InMux I__10798 (
            .O(N__47111),
            .I(N__47102));
    Odrv4 I__10797 (
            .O(N__47108),
            .I(\current_shift_inst.un4_control_input1_12 ));
    LocalMux I__10796 (
            .O(N__47105),
            .I(\current_shift_inst.un4_control_input1_12 ));
    LocalMux I__10795 (
            .O(N__47102),
            .I(\current_shift_inst.un4_control_input1_12 ));
    InMux I__10794 (
            .O(N__47095),
            .I(N__47092));
    LocalMux I__10793 (
            .O(N__47092),
            .I(N__47089));
    Span4Mux_h I__10792 (
            .O(N__47089),
            .I(N__47086));
    Span4Mux_h I__10791 (
            .O(N__47086),
            .I(N__47083));
    Odrv4 I__10790 (
            .O(N__47083),
            .I(\current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12 ));
    InMux I__10789 (
            .O(N__47080),
            .I(N__47073));
    InMux I__10788 (
            .O(N__47079),
            .I(N__47073));
    InMux I__10787 (
            .O(N__47078),
            .I(N__47070));
    LocalMux I__10786 (
            .O(N__47073),
            .I(N__47067));
    LocalMux I__10785 (
            .O(N__47070),
            .I(\current_shift_inst.un4_control_input1_7 ));
    Odrv4 I__10784 (
            .O(N__47067),
            .I(\current_shift_inst.un4_control_input1_7 ));
    InMux I__10783 (
            .O(N__47062),
            .I(N__47059));
    LocalMux I__10782 (
            .O(N__47059),
            .I(N__47056));
    Span4Mux_v I__10781 (
            .O(N__47056),
            .I(N__47053));
    Odrv4 I__10780 (
            .O(N__47053),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_7 ));
    InMux I__10779 (
            .O(N__47050),
            .I(N__47047));
    LocalMux I__10778 (
            .O(N__47047),
            .I(N__47044));
    Span4Mux_h I__10777 (
            .O(N__47044),
            .I(N__47041));
    Span4Mux_h I__10776 (
            .O(N__47041),
            .I(N__47038));
    Odrv4 I__10775 (
            .O(N__47038),
            .I(\current_shift_inst.un38_control_input_0_s0_11 ));
    InMux I__10774 (
            .O(N__47035),
            .I(N__47032));
    LocalMux I__10773 (
            .O(N__47032),
            .I(N__47029));
    Span4Mux_h I__10772 (
            .O(N__47029),
            .I(N__47026));
    Span4Mux_v I__10771 (
            .O(N__47026),
            .I(N__47023));
    Odrv4 I__10770 (
            .O(N__47023),
            .I(\current_shift_inst.un38_control_input_0_s1_11 ));
    InMux I__10769 (
            .O(N__47020),
            .I(N__47017));
    LocalMux I__10768 (
            .O(N__47017),
            .I(N__47014));
    Odrv12 I__10767 (
            .O(N__47014),
            .I(\current_shift_inst.control_input_1_axb_5 ));
    InMux I__10766 (
            .O(N__47011),
            .I(N__47008));
    LocalMux I__10765 (
            .O(N__47008),
            .I(N__47005));
    Span4Mux_v I__10764 (
            .O(N__47005),
            .I(N__47002));
    Span4Mux_h I__10763 (
            .O(N__47002),
            .I(N__46999));
    Odrv4 I__10762 (
            .O(N__46999),
            .I(\current_shift_inst.un38_control_input_0_s0_13 ));
    CascadeMux I__10761 (
            .O(N__46996),
            .I(N__46988));
    InMux I__10760 (
            .O(N__46995),
            .I(N__46981));
    InMux I__10759 (
            .O(N__46994),
            .I(N__46981));
    InMux I__10758 (
            .O(N__46993),
            .I(N__46981));
    CascadeMux I__10757 (
            .O(N__46992),
            .I(N__46976));
    CascadeMux I__10756 (
            .O(N__46991),
            .I(N__46966));
    InMux I__10755 (
            .O(N__46988),
            .I(N__46962));
    LocalMux I__10754 (
            .O(N__46981),
            .I(N__46959));
    InMux I__10753 (
            .O(N__46980),
            .I(N__46950));
    InMux I__10752 (
            .O(N__46979),
            .I(N__46950));
    InMux I__10751 (
            .O(N__46976),
            .I(N__46950));
    InMux I__10750 (
            .O(N__46975),
            .I(N__46950));
    InMux I__10749 (
            .O(N__46974),
            .I(N__46937));
    InMux I__10748 (
            .O(N__46973),
            .I(N__46937));
    InMux I__10747 (
            .O(N__46972),
            .I(N__46937));
    InMux I__10746 (
            .O(N__46971),
            .I(N__46937));
    InMux I__10745 (
            .O(N__46970),
            .I(N__46937));
    InMux I__10744 (
            .O(N__46969),
            .I(N__46937));
    InMux I__10743 (
            .O(N__46966),
            .I(N__46932));
    InMux I__10742 (
            .O(N__46965),
            .I(N__46932));
    LocalMux I__10741 (
            .O(N__46962),
            .I(N__46921));
    Span4Mux_h I__10740 (
            .O(N__46959),
            .I(N__46918));
    LocalMux I__10739 (
            .O(N__46950),
            .I(N__46915));
    LocalMux I__10738 (
            .O(N__46937),
            .I(N__46912));
    LocalMux I__10737 (
            .O(N__46932),
            .I(N__46909));
    CascadeMux I__10736 (
            .O(N__46931),
            .I(N__46906));
    CascadeMux I__10735 (
            .O(N__46930),
            .I(N__46903));
    CascadeMux I__10734 (
            .O(N__46929),
            .I(N__46898));
    InMux I__10733 (
            .O(N__46928),
            .I(N__46886));
    InMux I__10732 (
            .O(N__46927),
            .I(N__46886));
    InMux I__10731 (
            .O(N__46926),
            .I(N__46886));
    InMux I__10730 (
            .O(N__46925),
            .I(N__46886));
    InMux I__10729 (
            .O(N__46924),
            .I(N__46886));
    Span4Mux_v I__10728 (
            .O(N__46921),
            .I(N__46881));
    Span4Mux_v I__10727 (
            .O(N__46918),
            .I(N__46881));
    Span4Mux_h I__10726 (
            .O(N__46915),
            .I(N__46878));
    Span4Mux_h I__10725 (
            .O(N__46912),
            .I(N__46873));
    Span4Mux_h I__10724 (
            .O(N__46909),
            .I(N__46873));
    InMux I__10723 (
            .O(N__46906),
            .I(N__46860));
    InMux I__10722 (
            .O(N__46903),
            .I(N__46860));
    InMux I__10721 (
            .O(N__46902),
            .I(N__46860));
    InMux I__10720 (
            .O(N__46901),
            .I(N__46860));
    InMux I__10719 (
            .O(N__46898),
            .I(N__46860));
    InMux I__10718 (
            .O(N__46897),
            .I(N__46860));
    LocalMux I__10717 (
            .O(N__46886),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    Odrv4 I__10716 (
            .O(N__46881),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    Odrv4 I__10715 (
            .O(N__46878),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    Odrv4 I__10714 (
            .O(N__46873),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    LocalMux I__10713 (
            .O(N__46860),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    InMux I__10712 (
            .O(N__46849),
            .I(N__46846));
    LocalMux I__10711 (
            .O(N__46846),
            .I(N__46843));
    Span4Mux_h I__10710 (
            .O(N__46843),
            .I(N__46840));
    Span4Mux_v I__10709 (
            .O(N__46840),
            .I(N__46837));
    Odrv4 I__10708 (
            .O(N__46837),
            .I(\current_shift_inst.un38_control_input_0_s1_13 ));
    InMux I__10707 (
            .O(N__46834),
            .I(N__46831));
    LocalMux I__10706 (
            .O(N__46831),
            .I(N__46828));
    Odrv12 I__10705 (
            .O(N__46828),
            .I(\current_shift_inst.control_input_1_axb_7 ));
    InMux I__10704 (
            .O(N__46825),
            .I(N__46822));
    LocalMux I__10703 (
            .O(N__46822),
            .I(\current_shift_inst.un4_control_input_1_axb_3 ));
    InMux I__10702 (
            .O(N__46819),
            .I(N__46804));
    InMux I__10701 (
            .O(N__46818),
            .I(N__46804));
    InMux I__10700 (
            .O(N__46817),
            .I(N__46791));
    InMux I__10699 (
            .O(N__46816),
            .I(N__46791));
    InMux I__10698 (
            .O(N__46815),
            .I(N__46788));
    InMux I__10697 (
            .O(N__46814),
            .I(N__46785));
    InMux I__10696 (
            .O(N__46813),
            .I(N__46774));
    InMux I__10695 (
            .O(N__46812),
            .I(N__46774));
    InMux I__10694 (
            .O(N__46811),
            .I(N__46774));
    InMux I__10693 (
            .O(N__46810),
            .I(N__46774));
    InMux I__10692 (
            .O(N__46809),
            .I(N__46774));
    LocalMux I__10691 (
            .O(N__46804),
            .I(N__46768));
    InMux I__10690 (
            .O(N__46803),
            .I(N__46765));
    InMux I__10689 (
            .O(N__46802),
            .I(N__46762));
    InMux I__10688 (
            .O(N__46801),
            .I(N__46759));
    InMux I__10687 (
            .O(N__46800),
            .I(N__46753));
    InMux I__10686 (
            .O(N__46799),
            .I(N__46750));
    InMux I__10685 (
            .O(N__46798),
            .I(N__46746));
    CascadeMux I__10684 (
            .O(N__46797),
            .I(N__46736));
    InMux I__10683 (
            .O(N__46796),
            .I(N__46733));
    LocalMux I__10682 (
            .O(N__46791),
            .I(N__46724));
    LocalMux I__10681 (
            .O(N__46788),
            .I(N__46724));
    LocalMux I__10680 (
            .O(N__46785),
            .I(N__46724));
    LocalMux I__10679 (
            .O(N__46774),
            .I(N__46724));
    InMux I__10678 (
            .O(N__46773),
            .I(N__46717));
    InMux I__10677 (
            .O(N__46772),
            .I(N__46717));
    InMux I__10676 (
            .O(N__46771),
            .I(N__46717));
    Span4Mux_v I__10675 (
            .O(N__46768),
            .I(N__46708));
    LocalMux I__10674 (
            .O(N__46765),
            .I(N__46708));
    LocalMux I__10673 (
            .O(N__46762),
            .I(N__46708));
    LocalMux I__10672 (
            .O(N__46759),
            .I(N__46708));
    InMux I__10671 (
            .O(N__46758),
            .I(N__46671));
    InMux I__10670 (
            .O(N__46757),
            .I(N__46671));
    InMux I__10669 (
            .O(N__46756),
            .I(N__46671));
    LocalMux I__10668 (
            .O(N__46753),
            .I(N__46668));
    LocalMux I__10667 (
            .O(N__46750),
            .I(N__46665));
    InMux I__10666 (
            .O(N__46749),
            .I(N__46662));
    LocalMux I__10665 (
            .O(N__46746),
            .I(N__46659));
    InMux I__10664 (
            .O(N__46745),
            .I(N__46652));
    InMux I__10663 (
            .O(N__46744),
            .I(N__46652));
    InMux I__10662 (
            .O(N__46743),
            .I(N__46652));
    CascadeMux I__10661 (
            .O(N__46742),
            .I(N__46648));
    InMux I__10660 (
            .O(N__46741),
            .I(N__46644));
    InMux I__10659 (
            .O(N__46740),
            .I(N__46639));
    InMux I__10658 (
            .O(N__46739),
            .I(N__46639));
    InMux I__10657 (
            .O(N__46736),
            .I(N__46636));
    LocalMux I__10656 (
            .O(N__46733),
            .I(N__46633));
    Span4Mux_v I__10655 (
            .O(N__46724),
            .I(N__46628));
    LocalMux I__10654 (
            .O(N__46717),
            .I(N__46628));
    Span4Mux_v I__10653 (
            .O(N__46708),
            .I(N__46625));
    InMux I__10652 (
            .O(N__46707),
            .I(N__46622));
    InMux I__10651 (
            .O(N__46706),
            .I(N__46617));
    InMux I__10650 (
            .O(N__46705),
            .I(N__46617));
    InMux I__10649 (
            .O(N__46704),
            .I(N__46614));
    InMux I__10648 (
            .O(N__46703),
            .I(N__46609));
    InMux I__10647 (
            .O(N__46702),
            .I(N__46609));
    InMux I__10646 (
            .O(N__46701),
            .I(N__46604));
    InMux I__10645 (
            .O(N__46700),
            .I(N__46604));
    InMux I__10644 (
            .O(N__46699),
            .I(N__46593));
    InMux I__10643 (
            .O(N__46698),
            .I(N__46593));
    InMux I__10642 (
            .O(N__46697),
            .I(N__46593));
    InMux I__10641 (
            .O(N__46696),
            .I(N__46593));
    InMux I__10640 (
            .O(N__46695),
            .I(N__46593));
    InMux I__10639 (
            .O(N__46694),
            .I(N__46586));
    InMux I__10638 (
            .O(N__46693),
            .I(N__46586));
    InMux I__10637 (
            .O(N__46692),
            .I(N__46586));
    InMux I__10636 (
            .O(N__46691),
            .I(N__46577));
    InMux I__10635 (
            .O(N__46690),
            .I(N__46577));
    InMux I__10634 (
            .O(N__46689),
            .I(N__46577));
    InMux I__10633 (
            .O(N__46688),
            .I(N__46577));
    InMux I__10632 (
            .O(N__46687),
            .I(N__46566));
    InMux I__10631 (
            .O(N__46686),
            .I(N__46566));
    InMux I__10630 (
            .O(N__46685),
            .I(N__46566));
    InMux I__10629 (
            .O(N__46684),
            .I(N__46566));
    InMux I__10628 (
            .O(N__46683),
            .I(N__46566));
    InMux I__10627 (
            .O(N__46682),
            .I(N__46561));
    InMux I__10626 (
            .O(N__46681),
            .I(N__46561));
    InMux I__10625 (
            .O(N__46680),
            .I(N__46554));
    InMux I__10624 (
            .O(N__46679),
            .I(N__46554));
    InMux I__10623 (
            .O(N__46678),
            .I(N__46554));
    LocalMux I__10622 (
            .O(N__46671),
            .I(N__46551));
    Span4Mux_v I__10621 (
            .O(N__46668),
            .I(N__46544));
    Span4Mux_h I__10620 (
            .O(N__46665),
            .I(N__46544));
    LocalMux I__10619 (
            .O(N__46662),
            .I(N__46544));
    Span4Mux_h I__10618 (
            .O(N__46659),
            .I(N__46539));
    LocalMux I__10617 (
            .O(N__46652),
            .I(N__46539));
    InMux I__10616 (
            .O(N__46651),
            .I(N__46532));
    InMux I__10615 (
            .O(N__46648),
            .I(N__46532));
    InMux I__10614 (
            .O(N__46647),
            .I(N__46532));
    LocalMux I__10613 (
            .O(N__46644),
            .I(N__46522));
    LocalMux I__10612 (
            .O(N__46639),
            .I(N__46522));
    LocalMux I__10611 (
            .O(N__46636),
            .I(N__46517));
    Span4Mux_h I__10610 (
            .O(N__46633),
            .I(N__46517));
    Span4Mux_h I__10609 (
            .O(N__46628),
            .I(N__46514));
    Sp12to4 I__10608 (
            .O(N__46625),
            .I(N__46507));
    LocalMux I__10607 (
            .O(N__46622),
            .I(N__46507));
    LocalMux I__10606 (
            .O(N__46617),
            .I(N__46507));
    LocalMux I__10605 (
            .O(N__46614),
            .I(N__46504));
    LocalMux I__10604 (
            .O(N__46609),
            .I(N__46501));
    LocalMux I__10603 (
            .O(N__46604),
            .I(N__46490));
    LocalMux I__10602 (
            .O(N__46593),
            .I(N__46490));
    LocalMux I__10601 (
            .O(N__46586),
            .I(N__46490));
    LocalMux I__10600 (
            .O(N__46577),
            .I(N__46490));
    LocalMux I__10599 (
            .O(N__46566),
            .I(N__46490));
    LocalMux I__10598 (
            .O(N__46561),
            .I(N__46485));
    LocalMux I__10597 (
            .O(N__46554),
            .I(N__46485));
    Span4Mux_h I__10596 (
            .O(N__46551),
            .I(N__46482));
    Span4Mux_h I__10595 (
            .O(N__46544),
            .I(N__46477));
    Span4Mux_h I__10594 (
            .O(N__46539),
            .I(N__46477));
    LocalMux I__10593 (
            .O(N__46532),
            .I(N__46474));
    InMux I__10592 (
            .O(N__46531),
            .I(N__46467));
    InMux I__10591 (
            .O(N__46530),
            .I(N__46467));
    InMux I__10590 (
            .O(N__46529),
            .I(N__46467));
    InMux I__10589 (
            .O(N__46528),
            .I(N__46462));
    InMux I__10588 (
            .O(N__46527),
            .I(N__46462));
    Span4Mux_h I__10587 (
            .O(N__46522),
            .I(N__46457));
    Span4Mux_h I__10586 (
            .O(N__46517),
            .I(N__46457));
    Sp12to4 I__10585 (
            .O(N__46514),
            .I(N__46452));
    Span12Mux_h I__10584 (
            .O(N__46507),
            .I(N__46452));
    Span4Mux_h I__10583 (
            .O(N__46504),
            .I(N__46443));
    Span4Mux_h I__10582 (
            .O(N__46501),
            .I(N__46443));
    Span4Mux_v I__10581 (
            .O(N__46490),
            .I(N__46443));
    Span4Mux_v I__10580 (
            .O(N__46485),
            .I(N__46443));
    Span4Mux_h I__10579 (
            .O(N__46482),
            .I(N__46440));
    Odrv4 I__10578 (
            .O(N__46477),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__10577 (
            .O(N__46474),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__10576 (
            .O(N__46467),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__10575 (
            .O(N__46462),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__10574 (
            .O(N__46457),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv12 I__10573 (
            .O(N__46452),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__10572 (
            .O(N__46443),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__10571 (
            .O(N__46440),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    CascadeMux I__10570 (
            .O(N__46423),
            .I(N__46415));
    CascadeMux I__10569 (
            .O(N__46422),
            .I(N__46412));
    CascadeMux I__10568 (
            .O(N__46421),
            .I(N__46409));
    CascadeMux I__10567 (
            .O(N__46420),
            .I(N__46403));
    CascadeMux I__10566 (
            .O(N__46419),
            .I(N__46400));
    CascadeMux I__10565 (
            .O(N__46418),
            .I(N__46397));
    InMux I__10564 (
            .O(N__46415),
            .I(N__46392));
    InMux I__10563 (
            .O(N__46412),
            .I(N__46392));
    InMux I__10562 (
            .O(N__46409),
            .I(N__46389));
    CascadeMux I__10561 (
            .O(N__46408),
            .I(N__46386));
    CascadeMux I__10560 (
            .O(N__46407),
            .I(N__46383));
    CascadeMux I__10559 (
            .O(N__46406),
            .I(N__46380));
    InMux I__10558 (
            .O(N__46403),
            .I(N__46363));
    InMux I__10557 (
            .O(N__46400),
            .I(N__46358));
    InMux I__10556 (
            .O(N__46397),
            .I(N__46358));
    LocalMux I__10555 (
            .O(N__46392),
            .I(N__46353));
    LocalMux I__10554 (
            .O(N__46389),
            .I(N__46353));
    InMux I__10553 (
            .O(N__46386),
            .I(N__46348));
    InMux I__10552 (
            .O(N__46383),
            .I(N__46348));
    InMux I__10551 (
            .O(N__46380),
            .I(N__46345));
    CascadeMux I__10550 (
            .O(N__46379),
            .I(N__46336));
    CascadeMux I__10549 (
            .O(N__46378),
            .I(N__46316));
    CascadeMux I__10548 (
            .O(N__46377),
            .I(N__46312));
    CascadeMux I__10547 (
            .O(N__46376),
            .I(N__46309));
    CascadeMux I__10546 (
            .O(N__46375),
            .I(N__46306));
    CascadeMux I__10545 (
            .O(N__46374),
            .I(N__46298));
    CascadeMux I__10544 (
            .O(N__46373),
            .I(N__46287));
    CascadeMux I__10543 (
            .O(N__46372),
            .I(N__46284));
    CascadeMux I__10542 (
            .O(N__46371),
            .I(N__46280));
    CascadeMux I__10541 (
            .O(N__46370),
            .I(N__46277));
    CascadeMux I__10540 (
            .O(N__46369),
            .I(N__46270));
    CascadeMux I__10539 (
            .O(N__46368),
            .I(N__46267));
    CascadeMux I__10538 (
            .O(N__46367),
            .I(N__46264));
    CascadeMux I__10537 (
            .O(N__46366),
            .I(N__46261));
    LocalMux I__10536 (
            .O(N__46363),
            .I(N__46250));
    LocalMux I__10535 (
            .O(N__46358),
            .I(N__46250));
    Span4Mux_h I__10534 (
            .O(N__46353),
            .I(N__46243));
    LocalMux I__10533 (
            .O(N__46348),
            .I(N__46243));
    LocalMux I__10532 (
            .O(N__46345),
            .I(N__46243));
    CascadeMux I__10531 (
            .O(N__46344),
            .I(N__46240));
    CascadeMux I__10530 (
            .O(N__46343),
            .I(N__46237));
    CascadeMux I__10529 (
            .O(N__46342),
            .I(N__46234));
    CascadeMux I__10528 (
            .O(N__46341),
            .I(N__46225));
    CascadeMux I__10527 (
            .O(N__46340),
            .I(N__46222));
    InMux I__10526 (
            .O(N__46339),
            .I(N__46219));
    InMux I__10525 (
            .O(N__46336),
            .I(N__46205));
    CascadeMux I__10524 (
            .O(N__46335),
            .I(N__46202));
    CascadeMux I__10523 (
            .O(N__46334),
            .I(N__46199));
    CascadeMux I__10522 (
            .O(N__46333),
            .I(N__46196));
    CascadeMux I__10521 (
            .O(N__46332),
            .I(N__46193));
    CascadeMux I__10520 (
            .O(N__46331),
            .I(N__46190));
    CascadeMux I__10519 (
            .O(N__46330),
            .I(N__46187));
    CascadeMux I__10518 (
            .O(N__46329),
            .I(N__46184));
    CascadeMux I__10517 (
            .O(N__46328),
            .I(N__46181));
    CascadeMux I__10516 (
            .O(N__46327),
            .I(N__46178));
    CascadeMux I__10515 (
            .O(N__46326),
            .I(N__46175));
    CascadeMux I__10514 (
            .O(N__46325),
            .I(N__46172));
    CascadeMux I__10513 (
            .O(N__46324),
            .I(N__46169));
    CascadeMux I__10512 (
            .O(N__46323),
            .I(N__46165));
    CascadeMux I__10511 (
            .O(N__46322),
            .I(N__46162));
    CascadeMux I__10510 (
            .O(N__46321),
            .I(N__46159));
    CascadeMux I__10509 (
            .O(N__46320),
            .I(N__46156));
    CascadeMux I__10508 (
            .O(N__46319),
            .I(N__46153));
    InMux I__10507 (
            .O(N__46316),
            .I(N__46149));
    InMux I__10506 (
            .O(N__46315),
            .I(N__46140));
    InMux I__10505 (
            .O(N__46312),
            .I(N__46140));
    InMux I__10504 (
            .O(N__46309),
            .I(N__46140));
    InMux I__10503 (
            .O(N__46306),
            .I(N__46140));
    CascadeMux I__10502 (
            .O(N__46305),
            .I(N__46137));
    CascadeMux I__10501 (
            .O(N__46304),
            .I(N__46134));
    CascadeMux I__10500 (
            .O(N__46303),
            .I(N__46131));
    CascadeMux I__10499 (
            .O(N__46302),
            .I(N__46128));
    InMux I__10498 (
            .O(N__46301),
            .I(N__46123));
    InMux I__10497 (
            .O(N__46298),
            .I(N__46123));
    CascadeMux I__10496 (
            .O(N__46297),
            .I(N__46120));
    CascadeMux I__10495 (
            .O(N__46296),
            .I(N__46117));
    CascadeMux I__10494 (
            .O(N__46295),
            .I(N__46114));
    CascadeMux I__10493 (
            .O(N__46294),
            .I(N__46111));
    CascadeMux I__10492 (
            .O(N__46293),
            .I(N__46108));
    CascadeMux I__10491 (
            .O(N__46292),
            .I(N__46105));
    CascadeMux I__10490 (
            .O(N__46291),
            .I(N__46102));
    CascadeMux I__10489 (
            .O(N__46290),
            .I(N__46099));
    InMux I__10488 (
            .O(N__46287),
            .I(N__46095));
    InMux I__10487 (
            .O(N__46284),
            .I(N__46086));
    InMux I__10486 (
            .O(N__46283),
            .I(N__46086));
    InMux I__10485 (
            .O(N__46280),
            .I(N__46086));
    InMux I__10484 (
            .O(N__46277),
            .I(N__46086));
    CascadeMux I__10483 (
            .O(N__46276),
            .I(N__46083));
    CascadeMux I__10482 (
            .O(N__46275),
            .I(N__46080));
    CascadeMux I__10481 (
            .O(N__46274),
            .I(N__46077));
    CascadeMux I__10480 (
            .O(N__46273),
            .I(N__46074));
    InMux I__10479 (
            .O(N__46270),
            .I(N__46065));
    InMux I__10478 (
            .O(N__46267),
            .I(N__46065));
    InMux I__10477 (
            .O(N__46264),
            .I(N__46065));
    InMux I__10476 (
            .O(N__46261),
            .I(N__46065));
    CascadeMux I__10475 (
            .O(N__46260),
            .I(N__46062));
    CascadeMux I__10474 (
            .O(N__46259),
            .I(N__46059));
    CascadeMux I__10473 (
            .O(N__46258),
            .I(N__46056));
    CascadeMux I__10472 (
            .O(N__46257),
            .I(N__46053));
    CascadeMux I__10471 (
            .O(N__46256),
            .I(N__46050));
    CascadeMux I__10470 (
            .O(N__46255),
            .I(N__46047));
    Span4Mux_v I__10469 (
            .O(N__46250),
            .I(N__46042));
    Span4Mux_v I__10468 (
            .O(N__46243),
            .I(N__46042));
    InMux I__10467 (
            .O(N__46240),
            .I(N__46039));
    InMux I__10466 (
            .O(N__46237),
            .I(N__46034));
    InMux I__10465 (
            .O(N__46234),
            .I(N__46034));
    InMux I__10464 (
            .O(N__46233),
            .I(N__46027));
    InMux I__10463 (
            .O(N__46232),
            .I(N__46027));
    InMux I__10462 (
            .O(N__46231),
            .I(N__46027));
    CascadeMux I__10461 (
            .O(N__46230),
            .I(N__46023));
    CascadeMux I__10460 (
            .O(N__46229),
            .I(N__46020));
    CascadeMux I__10459 (
            .O(N__46228),
            .I(N__46016));
    InMux I__10458 (
            .O(N__46225),
            .I(N__46011));
    InMux I__10457 (
            .O(N__46222),
            .I(N__46011));
    LocalMux I__10456 (
            .O(N__46219),
            .I(N__46008));
    CascadeMux I__10455 (
            .O(N__46218),
            .I(N__46003));
    CascadeMux I__10454 (
            .O(N__46217),
            .I(N__46000));
    CascadeMux I__10453 (
            .O(N__46216),
            .I(N__45988));
    CascadeMux I__10452 (
            .O(N__46215),
            .I(N__45985));
    CascadeMux I__10451 (
            .O(N__46214),
            .I(N__45982));
    CascadeMux I__10450 (
            .O(N__46213),
            .I(N__45978));
    CascadeMux I__10449 (
            .O(N__46212),
            .I(N__45975));
    CascadeMux I__10448 (
            .O(N__46211),
            .I(N__45972));
    CascadeMux I__10447 (
            .O(N__46210),
            .I(N__45968));
    CascadeMux I__10446 (
            .O(N__46209),
            .I(N__45964));
    CascadeMux I__10445 (
            .O(N__46208),
            .I(N__45960));
    LocalMux I__10444 (
            .O(N__46205),
            .I(N__45956));
    InMux I__10443 (
            .O(N__46202),
            .I(N__45949));
    InMux I__10442 (
            .O(N__46199),
            .I(N__45949));
    InMux I__10441 (
            .O(N__46196),
            .I(N__45949));
    InMux I__10440 (
            .O(N__46193),
            .I(N__45940));
    InMux I__10439 (
            .O(N__46190),
            .I(N__45940));
    InMux I__10438 (
            .O(N__46187),
            .I(N__45940));
    InMux I__10437 (
            .O(N__46184),
            .I(N__45940));
    InMux I__10436 (
            .O(N__46181),
            .I(N__45931));
    InMux I__10435 (
            .O(N__46178),
            .I(N__45931));
    InMux I__10434 (
            .O(N__46175),
            .I(N__45931));
    InMux I__10433 (
            .O(N__46172),
            .I(N__45931));
    InMux I__10432 (
            .O(N__46169),
            .I(N__45922));
    CascadeMux I__10431 (
            .O(N__46168),
            .I(N__45918));
    InMux I__10430 (
            .O(N__46165),
            .I(N__45913));
    InMux I__10429 (
            .O(N__46162),
            .I(N__45913));
    InMux I__10428 (
            .O(N__46159),
            .I(N__45906));
    InMux I__10427 (
            .O(N__46156),
            .I(N__45906));
    InMux I__10426 (
            .O(N__46153),
            .I(N__45906));
    InMux I__10425 (
            .O(N__46152),
            .I(N__45903));
    LocalMux I__10424 (
            .O(N__46149),
            .I(N__45898));
    LocalMux I__10423 (
            .O(N__46140),
            .I(N__45898));
    InMux I__10422 (
            .O(N__46137),
            .I(N__45889));
    InMux I__10421 (
            .O(N__46134),
            .I(N__45889));
    InMux I__10420 (
            .O(N__46131),
            .I(N__45889));
    InMux I__10419 (
            .O(N__46128),
            .I(N__45889));
    LocalMux I__10418 (
            .O(N__46123),
            .I(N__45886));
    InMux I__10417 (
            .O(N__46120),
            .I(N__45877));
    InMux I__10416 (
            .O(N__46117),
            .I(N__45877));
    InMux I__10415 (
            .O(N__46114),
            .I(N__45877));
    InMux I__10414 (
            .O(N__46111),
            .I(N__45877));
    InMux I__10413 (
            .O(N__46108),
            .I(N__45870));
    InMux I__10412 (
            .O(N__46105),
            .I(N__45870));
    InMux I__10411 (
            .O(N__46102),
            .I(N__45870));
    InMux I__10410 (
            .O(N__46099),
            .I(N__45865));
    InMux I__10409 (
            .O(N__46098),
            .I(N__45865));
    LocalMux I__10408 (
            .O(N__46095),
            .I(N__45860));
    LocalMux I__10407 (
            .O(N__46086),
            .I(N__45860));
    InMux I__10406 (
            .O(N__46083),
            .I(N__45851));
    InMux I__10405 (
            .O(N__46080),
            .I(N__45851));
    InMux I__10404 (
            .O(N__46077),
            .I(N__45851));
    InMux I__10403 (
            .O(N__46074),
            .I(N__45851));
    LocalMux I__10402 (
            .O(N__46065),
            .I(N__45848));
    InMux I__10401 (
            .O(N__46062),
            .I(N__45841));
    InMux I__10400 (
            .O(N__46059),
            .I(N__45841));
    InMux I__10399 (
            .O(N__46056),
            .I(N__45841));
    InMux I__10398 (
            .O(N__46053),
            .I(N__45834));
    InMux I__10397 (
            .O(N__46050),
            .I(N__45834));
    InMux I__10396 (
            .O(N__46047),
            .I(N__45834));
    Span4Mux_h I__10395 (
            .O(N__46042),
            .I(N__45825));
    LocalMux I__10394 (
            .O(N__46039),
            .I(N__45825));
    LocalMux I__10393 (
            .O(N__46034),
            .I(N__45825));
    LocalMux I__10392 (
            .O(N__46027),
            .I(N__45825));
    InMux I__10391 (
            .O(N__46026),
            .I(N__45822));
    InMux I__10390 (
            .O(N__46023),
            .I(N__45817));
    InMux I__10389 (
            .O(N__46020),
            .I(N__45817));
    CascadeMux I__10388 (
            .O(N__46019),
            .I(N__45814));
    InMux I__10387 (
            .O(N__46016),
            .I(N__45811));
    LocalMux I__10386 (
            .O(N__46011),
            .I(N__45806));
    Span4Mux_h I__10385 (
            .O(N__46008),
            .I(N__45806));
    InMux I__10384 (
            .O(N__46007),
            .I(N__45801));
    InMux I__10383 (
            .O(N__46006),
            .I(N__45801));
    InMux I__10382 (
            .O(N__46003),
            .I(N__45796));
    InMux I__10381 (
            .O(N__46000),
            .I(N__45796));
    InMux I__10380 (
            .O(N__45999),
            .I(N__45793));
    CascadeMux I__10379 (
            .O(N__45998),
            .I(N__45790));
    CascadeMux I__10378 (
            .O(N__45997),
            .I(N__45787));
    CascadeMux I__10377 (
            .O(N__45996),
            .I(N__45784));
    CascadeMux I__10376 (
            .O(N__45995),
            .I(N__45781));
    CascadeMux I__10375 (
            .O(N__45994),
            .I(N__45778));
    CascadeMux I__10374 (
            .O(N__45993),
            .I(N__45775));
    CascadeMux I__10373 (
            .O(N__45992),
            .I(N__45772));
    CascadeMux I__10372 (
            .O(N__45991),
            .I(N__45769));
    InMux I__10371 (
            .O(N__45988),
            .I(N__45764));
    InMux I__10370 (
            .O(N__45985),
            .I(N__45764));
    InMux I__10369 (
            .O(N__45982),
            .I(N__45753));
    InMux I__10368 (
            .O(N__45981),
            .I(N__45753));
    InMux I__10367 (
            .O(N__45978),
            .I(N__45753));
    InMux I__10366 (
            .O(N__45975),
            .I(N__45753));
    InMux I__10365 (
            .O(N__45972),
            .I(N__45753));
    InMux I__10364 (
            .O(N__45971),
            .I(N__45738));
    InMux I__10363 (
            .O(N__45968),
            .I(N__45738));
    InMux I__10362 (
            .O(N__45967),
            .I(N__45738));
    InMux I__10361 (
            .O(N__45964),
            .I(N__45738));
    InMux I__10360 (
            .O(N__45963),
            .I(N__45738));
    InMux I__10359 (
            .O(N__45960),
            .I(N__45738));
    InMux I__10358 (
            .O(N__45959),
            .I(N__45738));
    Span4Mux_h I__10357 (
            .O(N__45956),
            .I(N__45729));
    LocalMux I__10356 (
            .O(N__45949),
            .I(N__45729));
    LocalMux I__10355 (
            .O(N__45940),
            .I(N__45729));
    LocalMux I__10354 (
            .O(N__45931),
            .I(N__45729));
    CascadeMux I__10353 (
            .O(N__45930),
            .I(N__45726));
    CascadeMux I__10352 (
            .O(N__45929),
            .I(N__45723));
    CascadeMux I__10351 (
            .O(N__45928),
            .I(N__45720));
    CascadeMux I__10350 (
            .O(N__45927),
            .I(N__45717));
    CascadeMux I__10349 (
            .O(N__45926),
            .I(N__45714));
    CascadeMux I__10348 (
            .O(N__45925),
            .I(N__45711));
    LocalMux I__10347 (
            .O(N__45922),
            .I(N__45708));
    InMux I__10346 (
            .O(N__45921),
            .I(N__45703));
    InMux I__10345 (
            .O(N__45918),
            .I(N__45703));
    LocalMux I__10344 (
            .O(N__45913),
            .I(N__45694));
    LocalMux I__10343 (
            .O(N__45906),
            .I(N__45694));
    LocalMux I__10342 (
            .O(N__45903),
            .I(N__45694));
    Span4Mux_v I__10341 (
            .O(N__45898),
            .I(N__45694));
    LocalMux I__10340 (
            .O(N__45889),
            .I(N__45673));
    Span4Mux_v I__10339 (
            .O(N__45886),
            .I(N__45673));
    LocalMux I__10338 (
            .O(N__45877),
            .I(N__45673));
    LocalMux I__10337 (
            .O(N__45870),
            .I(N__45673));
    LocalMux I__10336 (
            .O(N__45865),
            .I(N__45673));
    Span4Mux_v I__10335 (
            .O(N__45860),
            .I(N__45673));
    LocalMux I__10334 (
            .O(N__45851),
            .I(N__45673));
    Span4Mux_h I__10333 (
            .O(N__45848),
            .I(N__45673));
    LocalMux I__10332 (
            .O(N__45841),
            .I(N__45673));
    LocalMux I__10331 (
            .O(N__45834),
            .I(N__45673));
    Span4Mux_v I__10330 (
            .O(N__45825),
            .I(N__45670));
    LocalMux I__10329 (
            .O(N__45822),
            .I(N__45667));
    LocalMux I__10328 (
            .O(N__45817),
            .I(N__45664));
    InMux I__10327 (
            .O(N__45814),
            .I(N__45661));
    LocalMux I__10326 (
            .O(N__45811),
            .I(N__45656));
    Span4Mux_h I__10325 (
            .O(N__45806),
            .I(N__45656));
    LocalMux I__10324 (
            .O(N__45801),
            .I(N__45649));
    LocalMux I__10323 (
            .O(N__45796),
            .I(N__45649));
    LocalMux I__10322 (
            .O(N__45793),
            .I(N__45649));
    InMux I__10321 (
            .O(N__45790),
            .I(N__45640));
    InMux I__10320 (
            .O(N__45787),
            .I(N__45640));
    InMux I__10319 (
            .O(N__45784),
            .I(N__45640));
    InMux I__10318 (
            .O(N__45781),
            .I(N__45640));
    InMux I__10317 (
            .O(N__45778),
            .I(N__45631));
    InMux I__10316 (
            .O(N__45775),
            .I(N__45631));
    InMux I__10315 (
            .O(N__45772),
            .I(N__45631));
    InMux I__10314 (
            .O(N__45769),
            .I(N__45631));
    LocalMux I__10313 (
            .O(N__45764),
            .I(N__45622));
    LocalMux I__10312 (
            .O(N__45753),
            .I(N__45622));
    LocalMux I__10311 (
            .O(N__45738),
            .I(N__45622));
    Span4Mux_h I__10310 (
            .O(N__45729),
            .I(N__45622));
    InMux I__10309 (
            .O(N__45726),
            .I(N__45615));
    InMux I__10308 (
            .O(N__45723),
            .I(N__45615));
    InMux I__10307 (
            .O(N__45720),
            .I(N__45615));
    InMux I__10306 (
            .O(N__45717),
            .I(N__45608));
    InMux I__10305 (
            .O(N__45714),
            .I(N__45608));
    InMux I__10304 (
            .O(N__45711),
            .I(N__45608));
    Span4Mux_h I__10303 (
            .O(N__45708),
            .I(N__45599));
    LocalMux I__10302 (
            .O(N__45703),
            .I(N__45599));
    Span4Mux_v I__10301 (
            .O(N__45694),
            .I(N__45599));
    Span4Mux_v I__10300 (
            .O(N__45673),
            .I(N__45599));
    Odrv4 I__10299 (
            .O(N__45670),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv12 I__10298 (
            .O(N__45667),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv12 I__10297 (
            .O(N__45664),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10296 (
            .O(N__45661),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__10295 (
            .O(N__45656),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv12 I__10294 (
            .O(N__45649),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10293 (
            .O(N__45640),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10292 (
            .O(N__45631),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__10291 (
            .O(N__45622),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10290 (
            .O(N__45615),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10289 (
            .O(N__45608),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__10288 (
            .O(N__45599),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    InMux I__10287 (
            .O(N__45574),
            .I(N__45571));
    LocalMux I__10286 (
            .O(N__45571),
            .I(N__45567));
    InMux I__10285 (
            .O(N__45570),
            .I(N__45564));
    Span4Mux_v I__10284 (
            .O(N__45567),
            .I(N__45560));
    LocalMux I__10283 (
            .O(N__45564),
            .I(N__45557));
    InMux I__10282 (
            .O(N__45563),
            .I(N__45554));
    Odrv4 I__10281 (
            .O(N__45560),
            .I(\current_shift_inst.un4_control_input1_5 ));
    Odrv4 I__10280 (
            .O(N__45557),
            .I(\current_shift_inst.un4_control_input1_5 ));
    LocalMux I__10279 (
            .O(N__45554),
            .I(\current_shift_inst.un4_control_input1_5 ));
    InMux I__10278 (
            .O(N__45547),
            .I(N__45544));
    LocalMux I__10277 (
            .O(N__45544),
            .I(N__45541));
    Span4Mux_h I__10276 (
            .O(N__45541),
            .I(N__45538));
    Span4Mux_v I__10275 (
            .O(N__45538),
            .I(N__45535));
    Odrv4 I__10274 (
            .O(N__45535),
            .I(\current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0 ));
    InMux I__10273 (
            .O(N__45532),
            .I(N__45529));
    LocalMux I__10272 (
            .O(N__45529),
            .I(N__45526));
    Span4Mux_h I__10271 (
            .O(N__45526),
            .I(N__45523));
    Span4Mux_v I__10270 (
            .O(N__45523),
            .I(N__45520));
    Odrv4 I__10269 (
            .O(N__45520),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7 ));
    InMux I__10268 (
            .O(N__45517),
            .I(N__45513));
    InMux I__10267 (
            .O(N__45516),
            .I(N__45510));
    LocalMux I__10266 (
            .O(N__45513),
            .I(N__45507));
    LocalMux I__10265 (
            .O(N__45510),
            .I(N__45504));
    Span4Mux_v I__10264 (
            .O(N__45507),
            .I(N__45500));
    Span4Mux_h I__10263 (
            .O(N__45504),
            .I(N__45497));
    InMux I__10262 (
            .O(N__45503),
            .I(N__45494));
    Odrv4 I__10261 (
            .O(N__45500),
            .I(\current_shift_inst.un4_control_input1_17 ));
    Odrv4 I__10260 (
            .O(N__45497),
            .I(\current_shift_inst.un4_control_input1_17 ));
    LocalMux I__10259 (
            .O(N__45494),
            .I(\current_shift_inst.un4_control_input1_17 ));
    CascadeMux I__10258 (
            .O(N__45487),
            .I(N__45484));
    InMux I__10257 (
            .O(N__45484),
            .I(N__45481));
    LocalMux I__10256 (
            .O(N__45481),
            .I(N__45478));
    Span4Mux_v I__10255 (
            .O(N__45478),
            .I(N__45475));
    Span4Mux_h I__10254 (
            .O(N__45475),
            .I(N__45472));
    Odrv4 I__10253 (
            .O(N__45472),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISST11_0_17 ));
    InMux I__10252 (
            .O(N__45469),
            .I(N__45466));
    LocalMux I__10251 (
            .O(N__45466),
            .I(N__45463));
    Span4Mux_h I__10250 (
            .O(N__45463),
            .I(N__45460));
    Odrv4 I__10249 (
            .O(N__45460),
            .I(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ));
    InMux I__10248 (
            .O(N__45457),
            .I(N__45454));
    LocalMux I__10247 (
            .O(N__45454),
            .I(N__45451));
    Span4Mux_v I__10246 (
            .O(N__45451),
            .I(N__45448));
    Span4Mux_h I__10245 (
            .O(N__45448),
            .I(N__45445));
    Odrv4 I__10244 (
            .O(N__45445),
            .I(\current_shift_inst.un38_control_input_axb_31_s0 ));
    InMux I__10243 (
            .O(N__45442),
            .I(N__45437));
    InMux I__10242 (
            .O(N__45441),
            .I(N__45434));
    InMux I__10241 (
            .O(N__45440),
            .I(N__45431));
    LocalMux I__10240 (
            .O(N__45437),
            .I(N__45428));
    LocalMux I__10239 (
            .O(N__45434),
            .I(N__45425));
    LocalMux I__10238 (
            .O(N__45431),
            .I(N__45422));
    Span4Mux_h I__10237 (
            .O(N__45428),
            .I(N__45419));
    Span4Mux_v I__10236 (
            .O(N__45425),
            .I(N__45414));
    Span4Mux_h I__10235 (
            .O(N__45422),
            .I(N__45414));
    Odrv4 I__10234 (
            .O(N__45419),
            .I(\current_shift_inst.un4_control_input1_19 ));
    Odrv4 I__10233 (
            .O(N__45414),
            .I(\current_shift_inst.un4_control_input1_19 ));
    InMux I__10232 (
            .O(N__45409),
            .I(N__45406));
    LocalMux I__10231 (
            .O(N__45406),
            .I(N__45403));
    Span4Mux_h I__10230 (
            .O(N__45403),
            .I(N__45400));
    Odrv4 I__10229 (
            .O(N__45400),
            .I(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ));
    InMux I__10228 (
            .O(N__45397),
            .I(N__45394));
    LocalMux I__10227 (
            .O(N__45394),
            .I(N__45391));
    Span4Mux_h I__10226 (
            .O(N__45391),
            .I(N__45387));
    CascadeMux I__10225 (
            .O(N__45390),
            .I(N__45383));
    Span4Mux_h I__10224 (
            .O(N__45387),
            .I(N__45380));
    InMux I__10223 (
            .O(N__45386),
            .I(N__45377));
    InMux I__10222 (
            .O(N__45383),
            .I(N__45374));
    Odrv4 I__10221 (
            .O(N__45380),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    LocalMux I__10220 (
            .O(N__45377),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    LocalMux I__10219 (
            .O(N__45374),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    CascadeMux I__10218 (
            .O(N__45367),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ));
    InMux I__10217 (
            .O(N__45364),
            .I(N__45361));
    LocalMux I__10216 (
            .O(N__45361),
            .I(N__45357));
    InMux I__10215 (
            .O(N__45360),
            .I(N__45354));
    Span4Mux_v I__10214 (
            .O(N__45357),
            .I(N__45351));
    LocalMux I__10213 (
            .O(N__45354),
            .I(N__45348));
    Span4Mux_h I__10212 (
            .O(N__45351),
            .I(N__45343));
    Span4Mux_v I__10211 (
            .O(N__45348),
            .I(N__45343));
    Odrv4 I__10210 (
            .O(N__45343),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ));
    InMux I__10209 (
            .O(N__45340),
            .I(N__45335));
    InMux I__10208 (
            .O(N__45339),
            .I(N__45332));
    InMux I__10207 (
            .O(N__45338),
            .I(N__45329));
    LocalMux I__10206 (
            .O(N__45335),
            .I(N__45324));
    LocalMux I__10205 (
            .O(N__45332),
            .I(N__45324));
    LocalMux I__10204 (
            .O(N__45329),
            .I(N__45316));
    Span4Mux_h I__10203 (
            .O(N__45324),
            .I(N__45316));
    InMux I__10202 (
            .O(N__45323),
            .I(N__45311));
    InMux I__10201 (
            .O(N__45322),
            .I(N__45311));
    CascadeMux I__10200 (
            .O(N__45321),
            .I(N__45298));
    Span4Mux_v I__10199 (
            .O(N__45316),
            .I(N__45291));
    LocalMux I__10198 (
            .O(N__45311),
            .I(N__45291));
    InMux I__10197 (
            .O(N__45310),
            .I(N__45282));
    InMux I__10196 (
            .O(N__45309),
            .I(N__45282));
    InMux I__10195 (
            .O(N__45308),
            .I(N__45282));
    InMux I__10194 (
            .O(N__45307),
            .I(N__45282));
    InMux I__10193 (
            .O(N__45306),
            .I(N__45272));
    InMux I__10192 (
            .O(N__45305),
            .I(N__45272));
    InMux I__10191 (
            .O(N__45304),
            .I(N__45272));
    InMux I__10190 (
            .O(N__45303),
            .I(N__45265));
    InMux I__10189 (
            .O(N__45302),
            .I(N__45265));
    InMux I__10188 (
            .O(N__45301),
            .I(N__45265));
    InMux I__10187 (
            .O(N__45298),
            .I(N__45262));
    InMux I__10186 (
            .O(N__45297),
            .I(N__45257));
    InMux I__10185 (
            .O(N__45296),
            .I(N__45257));
    Span4Mux_h I__10184 (
            .O(N__45291),
            .I(N__45252));
    LocalMux I__10183 (
            .O(N__45282),
            .I(N__45252));
    InMux I__10182 (
            .O(N__45281),
            .I(N__45246));
    InMux I__10181 (
            .O(N__45280),
            .I(N__45243));
    InMux I__10180 (
            .O(N__45279),
            .I(N__45240));
    LocalMux I__10179 (
            .O(N__45272),
            .I(N__45232));
    LocalMux I__10178 (
            .O(N__45265),
            .I(N__45229));
    LocalMux I__10177 (
            .O(N__45262),
            .I(N__45224));
    LocalMux I__10176 (
            .O(N__45257),
            .I(N__45224));
    Span4Mux_v I__10175 (
            .O(N__45252),
            .I(N__45219));
    InMux I__10174 (
            .O(N__45251),
            .I(N__45212));
    InMux I__10173 (
            .O(N__45250),
            .I(N__45212));
    InMux I__10172 (
            .O(N__45249),
            .I(N__45212));
    LocalMux I__10171 (
            .O(N__45246),
            .I(N__45208));
    LocalMux I__10170 (
            .O(N__45243),
            .I(N__45205));
    LocalMux I__10169 (
            .O(N__45240),
            .I(N__45202));
    InMux I__10168 (
            .O(N__45239),
            .I(N__45191));
    InMux I__10167 (
            .O(N__45238),
            .I(N__45191));
    InMux I__10166 (
            .O(N__45237),
            .I(N__45191));
    InMux I__10165 (
            .O(N__45236),
            .I(N__45191));
    InMux I__10164 (
            .O(N__45235),
            .I(N__45191));
    Span4Mux_h I__10163 (
            .O(N__45232),
            .I(N__45188));
    Span4Mux_v I__10162 (
            .O(N__45229),
            .I(N__45183));
    Span4Mux_h I__10161 (
            .O(N__45224),
            .I(N__45183));
    InMux I__10160 (
            .O(N__45223),
            .I(N__45178));
    InMux I__10159 (
            .O(N__45222),
            .I(N__45178));
    Sp12to4 I__10158 (
            .O(N__45219),
            .I(N__45173));
    LocalMux I__10157 (
            .O(N__45212),
            .I(N__45173));
    InMux I__10156 (
            .O(N__45211),
            .I(N__45170));
    Span4Mux_h I__10155 (
            .O(N__45208),
            .I(N__45163));
    Span4Mux_v I__10154 (
            .O(N__45205),
            .I(N__45163));
    Span4Mux_v I__10153 (
            .O(N__45202),
            .I(N__45163));
    LocalMux I__10152 (
            .O(N__45191),
            .I(N__45158));
    Span4Mux_h I__10151 (
            .O(N__45188),
            .I(N__45158));
    Span4Mux_h I__10150 (
            .O(N__45183),
            .I(N__45155));
    LocalMux I__10149 (
            .O(N__45178),
            .I(N__45150));
    Span12Mux_h I__10148 (
            .O(N__45173),
            .I(N__45150));
    LocalMux I__10147 (
            .O(N__45170),
            .I(\current_shift_inst.PI_CTRL.N_74 ));
    Odrv4 I__10146 (
            .O(N__45163),
            .I(\current_shift_inst.PI_CTRL.N_74 ));
    Odrv4 I__10145 (
            .O(N__45158),
            .I(\current_shift_inst.PI_CTRL.N_74 ));
    Odrv4 I__10144 (
            .O(N__45155),
            .I(\current_shift_inst.PI_CTRL.N_74 ));
    Odrv12 I__10143 (
            .O(N__45150),
            .I(\current_shift_inst.PI_CTRL.N_74 ));
    CascadeMux I__10142 (
            .O(N__45139),
            .I(N__45127));
    InMux I__10141 (
            .O(N__45138),
            .I(N__45113));
    InMux I__10140 (
            .O(N__45137),
            .I(N__45105));
    InMux I__10139 (
            .O(N__45136),
            .I(N__45105));
    InMux I__10138 (
            .O(N__45135),
            .I(N__45105));
    InMux I__10137 (
            .O(N__45134),
            .I(N__45102));
    InMux I__10136 (
            .O(N__45133),
            .I(N__45099));
    InMux I__10135 (
            .O(N__45132),
            .I(N__45092));
    InMux I__10134 (
            .O(N__45131),
            .I(N__45092));
    InMux I__10133 (
            .O(N__45130),
            .I(N__45092));
    InMux I__10132 (
            .O(N__45127),
            .I(N__45085));
    InMux I__10131 (
            .O(N__45126),
            .I(N__45085));
    InMux I__10130 (
            .O(N__45125),
            .I(N__45085));
    InMux I__10129 (
            .O(N__45124),
            .I(N__45082));
    InMux I__10128 (
            .O(N__45123),
            .I(N__45077));
    InMux I__10127 (
            .O(N__45122),
            .I(N__45077));
    InMux I__10126 (
            .O(N__45121),
            .I(N__45068));
    InMux I__10125 (
            .O(N__45120),
            .I(N__45068));
    InMux I__10124 (
            .O(N__45119),
            .I(N__45068));
    InMux I__10123 (
            .O(N__45118),
            .I(N__45068));
    InMux I__10122 (
            .O(N__45117),
            .I(N__45057));
    InMux I__10121 (
            .O(N__45116),
            .I(N__45054));
    LocalMux I__10120 (
            .O(N__45113),
            .I(N__45051));
    InMux I__10119 (
            .O(N__45112),
            .I(N__45048));
    LocalMux I__10118 (
            .O(N__45105),
            .I(N__45043));
    LocalMux I__10117 (
            .O(N__45102),
            .I(N__45038));
    LocalMux I__10116 (
            .O(N__45099),
            .I(N__45038));
    LocalMux I__10115 (
            .O(N__45092),
            .I(N__45033));
    LocalMux I__10114 (
            .O(N__45085),
            .I(N__45033));
    LocalMux I__10113 (
            .O(N__45082),
            .I(N__45030));
    LocalMux I__10112 (
            .O(N__45077),
            .I(N__45027));
    LocalMux I__10111 (
            .O(N__45068),
            .I(N__45024));
    InMux I__10110 (
            .O(N__45067),
            .I(N__45021));
    InMux I__10109 (
            .O(N__45066),
            .I(N__45016));
    InMux I__10108 (
            .O(N__45065),
            .I(N__45016));
    InMux I__10107 (
            .O(N__45064),
            .I(N__45005));
    InMux I__10106 (
            .O(N__45063),
            .I(N__45005));
    InMux I__10105 (
            .O(N__45062),
            .I(N__45005));
    InMux I__10104 (
            .O(N__45061),
            .I(N__45005));
    InMux I__10103 (
            .O(N__45060),
            .I(N__45005));
    LocalMux I__10102 (
            .O(N__45057),
            .I(N__45000));
    LocalMux I__10101 (
            .O(N__45054),
            .I(N__45000));
    Span4Mux_h I__10100 (
            .O(N__45051),
            .I(N__44995));
    LocalMux I__10099 (
            .O(N__45048),
            .I(N__44995));
    InMux I__10098 (
            .O(N__45047),
            .I(N__44990));
    InMux I__10097 (
            .O(N__45046),
            .I(N__44990));
    Span4Mux_v I__10096 (
            .O(N__45043),
            .I(N__44983));
    Span4Mux_v I__10095 (
            .O(N__45038),
            .I(N__44983));
    Span4Mux_v I__10094 (
            .O(N__45033),
            .I(N__44983));
    Span4Mux_v I__10093 (
            .O(N__45030),
            .I(N__44976));
    Span4Mux_v I__10092 (
            .O(N__45027),
            .I(N__44976));
    Span4Mux_v I__10091 (
            .O(N__45024),
            .I(N__44976));
    LocalMux I__10090 (
            .O(N__45021),
            .I(N__44973));
    LocalMux I__10089 (
            .O(N__45016),
            .I(N__44966));
    LocalMux I__10088 (
            .O(N__45005),
            .I(N__44966));
    Span4Mux_h I__10087 (
            .O(N__45000),
            .I(N__44966));
    Span4Mux_h I__10086 (
            .O(N__44995),
            .I(N__44963));
    LocalMux I__10085 (
            .O(N__44990),
            .I(N__44956));
    Sp12to4 I__10084 (
            .O(N__44983),
            .I(N__44956));
    Sp12to4 I__10083 (
            .O(N__44976),
            .I(N__44956));
    Odrv4 I__10082 (
            .O(N__44973),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    Odrv4 I__10081 (
            .O(N__44966),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    Odrv4 I__10080 (
            .O(N__44963),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    Odrv12 I__10079 (
            .O(N__44956),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    InMux I__10078 (
            .O(N__44947),
            .I(N__44944));
    LocalMux I__10077 (
            .O(N__44944),
            .I(N__44941));
    Span4Mux_h I__10076 (
            .O(N__44941),
            .I(N__44938));
    Odrv4 I__10075 (
            .O(N__44938),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ));
    CascadeMux I__10074 (
            .O(N__44935),
            .I(N__44930));
    CascadeMux I__10073 (
            .O(N__44934),
            .I(N__44927));
    CascadeMux I__10072 (
            .O(N__44933),
            .I(N__44924));
    InMux I__10071 (
            .O(N__44930),
            .I(N__44906));
    InMux I__10070 (
            .O(N__44927),
            .I(N__44906));
    InMux I__10069 (
            .O(N__44924),
            .I(N__44903));
    CascadeMux I__10068 (
            .O(N__44923),
            .I(N__44900));
    CascadeMux I__10067 (
            .O(N__44922),
            .I(N__44897));
    CascadeMux I__10066 (
            .O(N__44921),
            .I(N__44894));
    CascadeMux I__10065 (
            .O(N__44920),
            .I(N__44891));
    CascadeMux I__10064 (
            .O(N__44919),
            .I(N__44888));
    CascadeMux I__10063 (
            .O(N__44918),
            .I(N__44885));
    CascadeMux I__10062 (
            .O(N__44917),
            .I(N__44880));
    CascadeMux I__10061 (
            .O(N__44916),
            .I(N__44877));
    CascadeMux I__10060 (
            .O(N__44915),
            .I(N__44874));
    CascadeMux I__10059 (
            .O(N__44914),
            .I(N__44871));
    InMux I__10058 (
            .O(N__44913),
            .I(N__44868));
    CascadeMux I__10057 (
            .O(N__44912),
            .I(N__44862));
    CascadeMux I__10056 (
            .O(N__44911),
            .I(N__44859));
    LocalMux I__10055 (
            .O(N__44906),
            .I(N__44856));
    LocalMux I__10054 (
            .O(N__44903),
            .I(N__44853));
    InMux I__10053 (
            .O(N__44900),
            .I(N__44849));
    InMux I__10052 (
            .O(N__44897),
            .I(N__44842));
    InMux I__10051 (
            .O(N__44894),
            .I(N__44842));
    InMux I__10050 (
            .O(N__44891),
            .I(N__44842));
    InMux I__10049 (
            .O(N__44888),
            .I(N__44837));
    InMux I__10048 (
            .O(N__44885),
            .I(N__44837));
    CascadeMux I__10047 (
            .O(N__44884),
            .I(N__44834));
    CascadeMux I__10046 (
            .O(N__44883),
            .I(N__44829));
    InMux I__10045 (
            .O(N__44880),
            .I(N__44826));
    InMux I__10044 (
            .O(N__44877),
            .I(N__44823));
    InMux I__10043 (
            .O(N__44874),
            .I(N__44818));
    InMux I__10042 (
            .O(N__44871),
            .I(N__44818));
    LocalMux I__10041 (
            .O(N__44868),
            .I(N__44815));
    InMux I__10040 (
            .O(N__44867),
            .I(N__44812));
    CascadeMux I__10039 (
            .O(N__44866),
            .I(N__44803));
    CascadeMux I__10038 (
            .O(N__44865),
            .I(N__44800));
    InMux I__10037 (
            .O(N__44862),
            .I(N__44794));
    InMux I__10036 (
            .O(N__44859),
            .I(N__44794));
    Span4Mux_h I__10035 (
            .O(N__44856),
            .I(N__44789));
    Span4Mux_h I__10034 (
            .O(N__44853),
            .I(N__44789));
    InMux I__10033 (
            .O(N__44852),
            .I(N__44786));
    LocalMux I__10032 (
            .O(N__44849),
            .I(N__44783));
    LocalMux I__10031 (
            .O(N__44842),
            .I(N__44778));
    LocalMux I__10030 (
            .O(N__44837),
            .I(N__44778));
    InMux I__10029 (
            .O(N__44834),
            .I(N__44775));
    CascadeMux I__10028 (
            .O(N__44833),
            .I(N__44772));
    CascadeMux I__10027 (
            .O(N__44832),
            .I(N__44769));
    InMux I__10026 (
            .O(N__44829),
            .I(N__44765));
    LocalMux I__10025 (
            .O(N__44826),
            .I(N__44754));
    LocalMux I__10024 (
            .O(N__44823),
            .I(N__44754));
    LocalMux I__10023 (
            .O(N__44818),
            .I(N__44754));
    Span4Mux_h I__10022 (
            .O(N__44815),
            .I(N__44754));
    LocalMux I__10021 (
            .O(N__44812),
            .I(N__44754));
    CascadeMux I__10020 (
            .O(N__44811),
            .I(N__44751));
    CascadeMux I__10019 (
            .O(N__44810),
            .I(N__44748));
    CascadeMux I__10018 (
            .O(N__44809),
            .I(N__44745));
    CascadeMux I__10017 (
            .O(N__44808),
            .I(N__44742));
    CascadeMux I__10016 (
            .O(N__44807),
            .I(N__44739));
    CascadeMux I__10015 (
            .O(N__44806),
            .I(N__44736));
    InMux I__10014 (
            .O(N__44803),
            .I(N__44731));
    InMux I__10013 (
            .O(N__44800),
            .I(N__44731));
    InMux I__10012 (
            .O(N__44799),
            .I(N__44728));
    LocalMux I__10011 (
            .O(N__44794),
            .I(N__44721));
    Span4Mux_v I__10010 (
            .O(N__44789),
            .I(N__44721));
    LocalMux I__10009 (
            .O(N__44786),
            .I(N__44721));
    Span4Mux_v I__10008 (
            .O(N__44783),
            .I(N__44714));
    Span4Mux_v I__10007 (
            .O(N__44778),
            .I(N__44714));
    LocalMux I__10006 (
            .O(N__44775),
            .I(N__44714));
    InMux I__10005 (
            .O(N__44772),
            .I(N__44711));
    InMux I__10004 (
            .O(N__44769),
            .I(N__44708));
    InMux I__10003 (
            .O(N__44768),
            .I(N__44705));
    LocalMux I__10002 (
            .O(N__44765),
            .I(N__44702));
    Span4Mux_h I__10001 (
            .O(N__44754),
            .I(N__44699));
    InMux I__10000 (
            .O(N__44751),
            .I(N__44694));
    InMux I__9999 (
            .O(N__44748),
            .I(N__44694));
    InMux I__9998 (
            .O(N__44745),
            .I(N__44689));
    InMux I__9997 (
            .O(N__44742),
            .I(N__44689));
    InMux I__9996 (
            .O(N__44739),
            .I(N__44684));
    InMux I__9995 (
            .O(N__44736),
            .I(N__44684));
    LocalMux I__9994 (
            .O(N__44731),
            .I(N__44675));
    LocalMux I__9993 (
            .O(N__44728),
            .I(N__44675));
    Span4Mux_v I__9992 (
            .O(N__44721),
            .I(N__44675));
    Span4Mux_h I__9991 (
            .O(N__44714),
            .I(N__44675));
    LocalMux I__9990 (
            .O(N__44711),
            .I(N__44664));
    LocalMux I__9989 (
            .O(N__44708),
            .I(N__44664));
    LocalMux I__9988 (
            .O(N__44705),
            .I(N__44664));
    Span4Mux_h I__9987 (
            .O(N__44702),
            .I(N__44664));
    Span4Mux_h I__9986 (
            .O(N__44699),
            .I(N__44664));
    LocalMux I__9985 (
            .O(N__44694),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__9984 (
            .O(N__44689),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__9983 (
            .O(N__44684),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__9982 (
            .O(N__44675),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__9981 (
            .O(N__44664),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    InMux I__9980 (
            .O(N__44653),
            .I(N__44647));
    InMux I__9979 (
            .O(N__44652),
            .I(N__44644));
    CascadeMux I__9978 (
            .O(N__44651),
            .I(N__44641));
    InMux I__9977 (
            .O(N__44650),
            .I(N__44638));
    LocalMux I__9976 (
            .O(N__44647),
            .I(N__44635));
    LocalMux I__9975 (
            .O(N__44644),
            .I(N__44632));
    InMux I__9974 (
            .O(N__44641),
            .I(N__44629));
    LocalMux I__9973 (
            .O(N__44638),
            .I(N__44626));
    Span4Mux_h I__9972 (
            .O(N__44635),
            .I(N__44622));
    Span4Mux_h I__9971 (
            .O(N__44632),
            .I(N__44619));
    LocalMux I__9970 (
            .O(N__44629),
            .I(N__44614));
    Span4Mux_h I__9969 (
            .O(N__44626),
            .I(N__44614));
    InMux I__9968 (
            .O(N__44625),
            .I(N__44611));
    Span4Mux_h I__9967 (
            .O(N__44622),
            .I(N__44606));
    Span4Mux_h I__9966 (
            .O(N__44619),
            .I(N__44606));
    Span4Mux_h I__9965 (
            .O(N__44614),
            .I(N__44603));
    LocalMux I__9964 (
            .O(N__44611),
            .I(N__44600));
    Odrv4 I__9963 (
            .O(N__44606),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv4 I__9962 (
            .O(N__44603),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv4 I__9961 (
            .O(N__44600),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    CascadeMux I__9960 (
            .O(N__44593),
            .I(N__44590));
    InMux I__9959 (
            .O(N__44590),
            .I(N__44587));
    LocalMux I__9958 (
            .O(N__44587),
            .I(N__44584));
    Odrv4 I__9957 (
            .O(N__44584),
            .I(\current_shift_inst.PI_CTRL.integrator_i_26 ));
    CascadeMux I__9956 (
            .O(N__44581),
            .I(N__44578));
    InMux I__9955 (
            .O(N__44578),
            .I(N__44574));
    InMux I__9954 (
            .O(N__44577),
            .I(N__44570));
    LocalMux I__9953 (
            .O(N__44574),
            .I(N__44567));
    InMux I__9952 (
            .O(N__44573),
            .I(N__44564));
    LocalMux I__9951 (
            .O(N__44570),
            .I(N__44559));
    Span4Mux_h I__9950 (
            .O(N__44567),
            .I(N__44556));
    LocalMux I__9949 (
            .O(N__44564),
            .I(N__44553));
    InMux I__9948 (
            .O(N__44563),
            .I(N__44550));
    InMux I__9947 (
            .O(N__44562),
            .I(N__44547));
    Span4Mux_h I__9946 (
            .O(N__44559),
            .I(N__44544));
    Odrv4 I__9945 (
            .O(N__44556),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv4 I__9944 (
            .O(N__44553),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    LocalMux I__9943 (
            .O(N__44550),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    LocalMux I__9942 (
            .O(N__44547),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv4 I__9941 (
            .O(N__44544),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    CascadeMux I__9940 (
            .O(N__44533),
            .I(N__44530));
    InMux I__9939 (
            .O(N__44530),
            .I(N__44527));
    LocalMux I__9938 (
            .O(N__44527),
            .I(N__44524));
    Odrv4 I__9937 (
            .O(N__44524),
            .I(\current_shift_inst.PI_CTRL.integrator_i_24 ));
    InMux I__9936 (
            .O(N__44521),
            .I(N__44517));
    CascadeMux I__9935 (
            .O(N__44520),
            .I(N__44514));
    LocalMux I__9934 (
            .O(N__44517),
            .I(N__44510));
    InMux I__9933 (
            .O(N__44514),
            .I(N__44507));
    InMux I__9932 (
            .O(N__44513),
            .I(N__44504));
    Span4Mux_v I__9931 (
            .O(N__44510),
            .I(N__44501));
    LocalMux I__9930 (
            .O(N__44507),
            .I(N__44498));
    LocalMux I__9929 (
            .O(N__44504),
            .I(N__44495));
    Span4Mux_h I__9928 (
            .O(N__44501),
            .I(N__44490));
    Span4Mux_h I__9927 (
            .O(N__44498),
            .I(N__44490));
    Span12Mux_h I__9926 (
            .O(N__44495),
            .I(N__44486));
    Span4Mux_h I__9925 (
            .O(N__44490),
            .I(N__44483));
    InMux I__9924 (
            .O(N__44489),
            .I(N__44480));
    Odrv12 I__9923 (
            .O(N__44486),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    Odrv4 I__9922 (
            .O(N__44483),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    LocalMux I__9921 (
            .O(N__44480),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    CascadeMux I__9920 (
            .O(N__44473),
            .I(N__44470));
    InMux I__9919 (
            .O(N__44470),
            .I(N__44467));
    LocalMux I__9918 (
            .O(N__44467),
            .I(N__44464));
    Odrv4 I__9917 (
            .O(N__44464),
            .I(\current_shift_inst.PI_CTRL.integrator_i_28 ));
    CascadeMux I__9916 (
            .O(N__44461),
            .I(N__44458));
    InMux I__9915 (
            .O(N__44458),
            .I(N__44455));
    LocalMux I__9914 (
            .O(N__44455),
            .I(N__44450));
    InMux I__9913 (
            .O(N__44454),
            .I(N__44447));
    InMux I__9912 (
            .O(N__44453),
            .I(N__44444));
    Span4Mux_v I__9911 (
            .O(N__44450),
            .I(N__44438));
    LocalMux I__9910 (
            .O(N__44447),
            .I(N__44438));
    LocalMux I__9909 (
            .O(N__44444),
            .I(N__44435));
    InMux I__9908 (
            .O(N__44443),
            .I(N__44432));
    Span4Mux_h I__9907 (
            .O(N__44438),
            .I(N__44428));
    Span4Mux_h I__9906 (
            .O(N__44435),
            .I(N__44425));
    LocalMux I__9905 (
            .O(N__44432),
            .I(N__44422));
    InMux I__9904 (
            .O(N__44431),
            .I(N__44419));
    Span4Mux_h I__9903 (
            .O(N__44428),
            .I(N__44416));
    Odrv4 I__9902 (
            .O(N__44425),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    Odrv12 I__9901 (
            .O(N__44422),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    LocalMux I__9900 (
            .O(N__44419),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    Odrv4 I__9899 (
            .O(N__44416),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    CascadeMux I__9898 (
            .O(N__44407),
            .I(N__44404));
    InMux I__9897 (
            .O(N__44404),
            .I(N__44401));
    LocalMux I__9896 (
            .O(N__44401),
            .I(N__44398));
    Odrv4 I__9895 (
            .O(N__44398),
            .I(\current_shift_inst.PI_CTRL.integrator_i_23 ));
    InMux I__9894 (
            .O(N__44395),
            .I(N__44392));
    LocalMux I__9893 (
            .O(N__44392),
            .I(N__44389));
    Span4Mux_h I__9892 (
            .O(N__44389),
            .I(N__44386));
    Odrv4 I__9891 (
            .O(N__44386),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    InMux I__9890 (
            .O(N__44383),
            .I(N__44380));
    LocalMux I__9889 (
            .O(N__44380),
            .I(N__44377));
    Span4Mux_h I__9888 (
            .O(N__44377),
            .I(N__44374));
    Odrv4 I__9887 (
            .O(N__44374),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    CascadeMux I__9886 (
            .O(N__44371),
            .I(N__44368));
    InMux I__9885 (
            .O(N__44368),
            .I(N__44365));
    LocalMux I__9884 (
            .O(N__44365),
            .I(N__44362));
    Span4Mux_h I__9883 (
            .O(N__44362),
            .I(N__44359));
    Odrv4 I__9882 (
            .O(N__44359),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    InMux I__9881 (
            .O(N__44356),
            .I(N__44353));
    LocalMux I__9880 (
            .O(N__44353),
            .I(N__44350));
    Span4Mux_v I__9879 (
            .O(N__44350),
            .I(N__44347));
    Odrv4 I__9878 (
            .O(N__44347),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    InMux I__9877 (
            .O(N__44344),
            .I(N__44341));
    LocalMux I__9876 (
            .O(N__44341),
            .I(N__44338));
    Span12Mux_h I__9875 (
            .O(N__44338),
            .I(N__44335));
    Odrv12 I__9874 (
            .O(N__44335),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19 ));
    InMux I__9873 (
            .O(N__44332),
            .I(N__44328));
    InMux I__9872 (
            .O(N__44331),
            .I(N__44324));
    LocalMux I__9871 (
            .O(N__44328),
            .I(N__44321));
    InMux I__9870 (
            .O(N__44327),
            .I(N__44318));
    LocalMux I__9869 (
            .O(N__44324),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    Odrv4 I__9868 (
            .O(N__44321),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__9867 (
            .O(N__44318),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    InMux I__9866 (
            .O(N__44311),
            .I(N__44307));
    InMux I__9865 (
            .O(N__44310),
            .I(N__44304));
    LocalMux I__9864 (
            .O(N__44307),
            .I(N__44298));
    LocalMux I__9863 (
            .O(N__44304),
            .I(N__44298));
    InMux I__9862 (
            .O(N__44303),
            .I(N__44295));
    Span4Mux_h I__9861 (
            .O(N__44298),
            .I(N__44292));
    LocalMux I__9860 (
            .O(N__44295),
            .I(N__44289));
    Span4Mux_h I__9859 (
            .O(N__44292),
            .I(N__44286));
    Odrv12 I__9858 (
            .O(N__44289),
            .I(\delay_measurement_inst.elapsed_time_tr_2 ));
    Odrv4 I__9857 (
            .O(N__44286),
            .I(\delay_measurement_inst.elapsed_time_tr_2 ));
    CascadeMux I__9856 (
            .O(N__44281),
            .I(N__44278));
    InMux I__9855 (
            .O(N__44278),
            .I(N__44275));
    LocalMux I__9854 (
            .O(N__44275),
            .I(N__44272));
    Span4Mux_v I__9853 (
            .O(N__44272),
            .I(N__44269));
    Odrv4 I__9852 (
            .O(N__44269),
            .I(\current_shift_inst.un4_control_input_1_axb_27 ));
    InMux I__9851 (
            .O(N__44266),
            .I(N__44262));
    InMux I__9850 (
            .O(N__44265),
            .I(N__44259));
    LocalMux I__9849 (
            .O(N__44262),
            .I(N__44256));
    LocalMux I__9848 (
            .O(N__44259),
            .I(N__44253));
    Span4Mux_h I__9847 (
            .O(N__44256),
            .I(N__44249));
    Span12Mux_h I__9846 (
            .O(N__44253),
            .I(N__44246));
    InMux I__9845 (
            .O(N__44252),
            .I(N__44243));
    Odrv4 I__9844 (
            .O(N__44249),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_17 ));
    Odrv12 I__9843 (
            .O(N__44246),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_17 ));
    LocalMux I__9842 (
            .O(N__44243),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_17 ));
    InMux I__9841 (
            .O(N__44236),
            .I(N__44233));
    LocalMux I__9840 (
            .O(N__44233),
            .I(N__44230));
    Odrv12 I__9839 (
            .O(N__44230),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_17 ));
    InMux I__9838 (
            .O(N__44227),
            .I(N__44224));
    LocalMux I__9837 (
            .O(N__44224),
            .I(N__44221));
    Odrv4 I__9836 (
            .O(N__44221),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIKOBPZ0Z_17 ));
    CascadeMux I__9835 (
            .O(N__44218),
            .I(N__44215));
    InMux I__9834 (
            .O(N__44215),
            .I(N__44212));
    LocalMux I__9833 (
            .O(N__44212),
            .I(N__44209));
    Span4Mux_h I__9832 (
            .O(N__44209),
            .I(N__44206));
    Odrv4 I__9831 (
            .O(N__44206),
            .I(\current_shift_inst.PI_CTRL.integrator_i_10 ));
    CascadeMux I__9830 (
            .O(N__44203),
            .I(N__44198));
    InMux I__9829 (
            .O(N__44202),
            .I(N__44195));
    InMux I__9828 (
            .O(N__44201),
            .I(N__44192));
    InMux I__9827 (
            .O(N__44198),
            .I(N__44189));
    LocalMux I__9826 (
            .O(N__44195),
            .I(N__44186));
    LocalMux I__9825 (
            .O(N__44192),
            .I(N__44183));
    LocalMux I__9824 (
            .O(N__44189),
            .I(N__44180));
    Span4Mux_h I__9823 (
            .O(N__44186),
            .I(N__44173));
    Span4Mux_v I__9822 (
            .O(N__44183),
            .I(N__44173));
    Span4Mux_h I__9821 (
            .O(N__44180),
            .I(N__44170));
    InMux I__9820 (
            .O(N__44179),
            .I(N__44167));
    InMux I__9819 (
            .O(N__44178),
            .I(N__44164));
    Span4Mux_h I__9818 (
            .O(N__44173),
            .I(N__44161));
    Odrv4 I__9817 (
            .O(N__44170),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    LocalMux I__9816 (
            .O(N__44167),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    LocalMux I__9815 (
            .O(N__44164),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    Odrv4 I__9814 (
            .O(N__44161),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    CascadeMux I__9813 (
            .O(N__44152),
            .I(N__44149));
    InMux I__9812 (
            .O(N__44149),
            .I(N__44146));
    LocalMux I__9811 (
            .O(N__44146),
            .I(N__44143));
    Odrv4 I__9810 (
            .O(N__44143),
            .I(\current_shift_inst.PI_CTRL.integrator_i_7 ));
    CascadeMux I__9809 (
            .O(N__44140),
            .I(N__44136));
    InMux I__9808 (
            .O(N__44139),
            .I(N__44132));
    InMux I__9807 (
            .O(N__44136),
            .I(N__44127));
    InMux I__9806 (
            .O(N__44135),
            .I(N__44127));
    LocalMux I__9805 (
            .O(N__44132),
            .I(N__44123));
    LocalMux I__9804 (
            .O(N__44127),
            .I(N__44120));
    CascadeMux I__9803 (
            .O(N__44126),
            .I(N__44116));
    Span4Mux_h I__9802 (
            .O(N__44123),
            .I(N__44111));
    Span4Mux_h I__9801 (
            .O(N__44120),
            .I(N__44111));
    InMux I__9800 (
            .O(N__44119),
            .I(N__44108));
    InMux I__9799 (
            .O(N__44116),
            .I(N__44105));
    Span4Mux_h I__9798 (
            .O(N__44111),
            .I(N__44102));
    LocalMux I__9797 (
            .O(N__44108),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    LocalMux I__9796 (
            .O(N__44105),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    Odrv4 I__9795 (
            .O(N__44102),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    CascadeMux I__9794 (
            .O(N__44095),
            .I(N__44092));
    InMux I__9793 (
            .O(N__44092),
            .I(N__44089));
    LocalMux I__9792 (
            .O(N__44089),
            .I(N__44086));
    Odrv4 I__9791 (
            .O(N__44086),
            .I(\current_shift_inst.PI_CTRL.integrator_i_13 ));
    InMux I__9790 (
            .O(N__44083),
            .I(N__44074));
    InMux I__9789 (
            .O(N__44082),
            .I(N__44063));
    InMux I__9788 (
            .O(N__44081),
            .I(N__44060));
    InMux I__9787 (
            .O(N__44080),
            .I(N__44057));
    InMux I__9786 (
            .O(N__44079),
            .I(N__44046));
    InMux I__9785 (
            .O(N__44078),
            .I(N__44043));
    InMux I__9784 (
            .O(N__44077),
            .I(N__44040));
    LocalMux I__9783 (
            .O(N__44074),
            .I(N__44037));
    InMux I__9782 (
            .O(N__44073),
            .I(N__44020));
    InMux I__9781 (
            .O(N__44072),
            .I(N__44020));
    InMux I__9780 (
            .O(N__44071),
            .I(N__44020));
    InMux I__9779 (
            .O(N__44070),
            .I(N__44020));
    InMux I__9778 (
            .O(N__44069),
            .I(N__44020));
    InMux I__9777 (
            .O(N__44068),
            .I(N__44020));
    InMux I__9776 (
            .O(N__44067),
            .I(N__44020));
    InMux I__9775 (
            .O(N__44066),
            .I(N__44020));
    LocalMux I__9774 (
            .O(N__44063),
            .I(N__44010));
    LocalMux I__9773 (
            .O(N__44060),
            .I(N__44010));
    LocalMux I__9772 (
            .O(N__44057),
            .I(N__44010));
    InMux I__9771 (
            .O(N__44056),
            .I(N__43999));
    InMux I__9770 (
            .O(N__44055),
            .I(N__43999));
    InMux I__9769 (
            .O(N__44054),
            .I(N__43999));
    InMux I__9768 (
            .O(N__44053),
            .I(N__43999));
    InMux I__9767 (
            .O(N__44052),
            .I(N__43999));
    InMux I__9766 (
            .O(N__44051),
            .I(N__43993));
    InMux I__9765 (
            .O(N__44050),
            .I(N__43988));
    InMux I__9764 (
            .O(N__44049),
            .I(N__43988));
    LocalMux I__9763 (
            .O(N__44046),
            .I(N__43977));
    LocalMux I__9762 (
            .O(N__44043),
            .I(N__43974));
    LocalMux I__9761 (
            .O(N__44040),
            .I(N__43967));
    Span4Mux_v I__9760 (
            .O(N__44037),
            .I(N__43967));
    LocalMux I__9759 (
            .O(N__44020),
            .I(N__43967));
    InMux I__9758 (
            .O(N__44019),
            .I(N__43962));
    InMux I__9757 (
            .O(N__44018),
            .I(N__43962));
    InMux I__9756 (
            .O(N__44017),
            .I(N__43959));
    Span4Mux_v I__9755 (
            .O(N__44010),
            .I(N__43954));
    LocalMux I__9754 (
            .O(N__43999),
            .I(N__43954));
    InMux I__9753 (
            .O(N__43998),
            .I(N__43949));
    InMux I__9752 (
            .O(N__43997),
            .I(N__43949));
    InMux I__9751 (
            .O(N__43996),
            .I(N__43946));
    LocalMux I__9750 (
            .O(N__43993),
            .I(N__43941));
    LocalMux I__9749 (
            .O(N__43988),
            .I(N__43941));
    InMux I__9748 (
            .O(N__43987),
            .I(N__43928));
    InMux I__9747 (
            .O(N__43986),
            .I(N__43928));
    InMux I__9746 (
            .O(N__43985),
            .I(N__43928));
    InMux I__9745 (
            .O(N__43984),
            .I(N__43928));
    InMux I__9744 (
            .O(N__43983),
            .I(N__43928));
    InMux I__9743 (
            .O(N__43982),
            .I(N__43928));
    InMux I__9742 (
            .O(N__43981),
            .I(N__43923));
    InMux I__9741 (
            .O(N__43980),
            .I(N__43923));
    Span4Mux_h I__9740 (
            .O(N__43977),
            .I(N__43920));
    Span4Mux_v I__9739 (
            .O(N__43974),
            .I(N__43913));
    Span4Mux_h I__9738 (
            .O(N__43967),
            .I(N__43913));
    LocalMux I__9737 (
            .O(N__43962),
            .I(N__43913));
    LocalMux I__9736 (
            .O(N__43959),
            .I(N__43908));
    Span4Mux_h I__9735 (
            .O(N__43954),
            .I(N__43908));
    LocalMux I__9734 (
            .O(N__43949),
            .I(N__43901));
    LocalMux I__9733 (
            .O(N__43946),
            .I(N__43901));
    Span4Mux_v I__9732 (
            .O(N__43941),
            .I(N__43901));
    LocalMux I__9731 (
            .O(N__43928),
            .I(N__43898));
    LocalMux I__9730 (
            .O(N__43923),
            .I(N__43891));
    Span4Mux_v I__9729 (
            .O(N__43920),
            .I(N__43891));
    Span4Mux_h I__9728 (
            .O(N__43913),
            .I(N__43891));
    Span4Mux_v I__9727 (
            .O(N__43908),
            .I(N__43888));
    Span4Mux_v I__9726 (
            .O(N__43901),
            .I(N__43885));
    Span4Mux_h I__9725 (
            .O(N__43898),
            .I(N__43882));
    Odrv4 I__9724 (
            .O(N__43891),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_26 ));
    Odrv4 I__9723 (
            .O(N__43888),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_26 ));
    Odrv4 I__9722 (
            .O(N__43885),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_26 ));
    Odrv4 I__9721 (
            .O(N__43882),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_26 ));
    InMux I__9720 (
            .O(N__43873),
            .I(N__43869));
    InMux I__9719 (
            .O(N__43872),
            .I(N__43866));
    LocalMux I__9718 (
            .O(N__43869),
            .I(N__43863));
    LocalMux I__9717 (
            .O(N__43866),
            .I(N__43860));
    Span4Mux_v I__9716 (
            .O(N__43863),
            .I(N__43856));
    Span4Mux_h I__9715 (
            .O(N__43860),
            .I(N__43853));
    InMux I__9714 (
            .O(N__43859),
            .I(N__43850));
    Span4Mux_h I__9713 (
            .O(N__43856),
            .I(N__43845));
    Span4Mux_h I__9712 (
            .O(N__43853),
            .I(N__43845));
    LocalMux I__9711 (
            .O(N__43850),
            .I(N__43842));
    Odrv4 I__9710 (
            .O(N__43845),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    Odrv4 I__9709 (
            .O(N__43842),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    InMux I__9708 (
            .O(N__43837),
            .I(N__43834));
    LocalMux I__9707 (
            .O(N__43834),
            .I(N__43831));
    Span4Mux_h I__9706 (
            .O(N__43831),
            .I(N__43828));
    Odrv4 I__9705 (
            .O(N__43828),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_14 ));
    InMux I__9704 (
            .O(N__43825),
            .I(N__43822));
    LocalMux I__9703 (
            .O(N__43822),
            .I(N__43819));
    Span4Mux_v I__9702 (
            .O(N__43819),
            .I(N__43816));
    Odrv4 I__9701 (
            .O(N__43816),
            .I(\current_shift_inst.PI_CTRL.error_control_RNI898PZ0Z_14 ));
    InMux I__9700 (
            .O(N__43813),
            .I(N__43810));
    LocalMux I__9699 (
            .O(N__43810),
            .I(N__43807));
    Span4Mux_h I__9698 (
            .O(N__43807),
            .I(N__43804));
    Odrv4 I__9697 (
            .O(N__43804),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ));
    InMux I__9696 (
            .O(N__43801),
            .I(N__43798));
    LocalMux I__9695 (
            .O(N__43798),
            .I(N__43794));
    InMux I__9694 (
            .O(N__43797),
            .I(N__43790));
    Span4Mux_v I__9693 (
            .O(N__43794),
            .I(N__43786));
    CascadeMux I__9692 (
            .O(N__43793),
            .I(N__43782));
    LocalMux I__9691 (
            .O(N__43790),
            .I(N__43779));
    InMux I__9690 (
            .O(N__43789),
            .I(N__43776));
    Span4Mux_h I__9689 (
            .O(N__43786),
            .I(N__43773));
    InMux I__9688 (
            .O(N__43785),
            .I(N__43770));
    InMux I__9687 (
            .O(N__43782),
            .I(N__43767));
    Span12Mux_s9_v I__9686 (
            .O(N__43779),
            .I(N__43762));
    LocalMux I__9685 (
            .O(N__43776),
            .I(N__43762));
    Span4Mux_h I__9684 (
            .O(N__43773),
            .I(N__43757));
    LocalMux I__9683 (
            .O(N__43770),
            .I(N__43757));
    LocalMux I__9682 (
            .O(N__43767),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    Odrv12 I__9681 (
            .O(N__43762),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    Odrv4 I__9680 (
            .O(N__43757),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    InMux I__9679 (
            .O(N__43750),
            .I(N__43747));
    LocalMux I__9678 (
            .O(N__43747),
            .I(N__43744));
    Span4Mux_h I__9677 (
            .O(N__43744),
            .I(N__43741));
    Odrv4 I__9676 (
            .O(N__43741),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ));
    InMux I__9675 (
            .O(N__43738),
            .I(N__43735));
    LocalMux I__9674 (
            .O(N__43735),
            .I(N__43732));
    Span4Mux_v I__9673 (
            .O(N__43732),
            .I(N__43729));
    Odrv4 I__9672 (
            .O(N__43729),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ));
    InMux I__9671 (
            .O(N__43726),
            .I(N__43723));
    LocalMux I__9670 (
            .O(N__43723),
            .I(N__43720));
    Odrv12 I__9669 (
            .O(N__43720),
            .I(\current_shift_inst.un4_control_input_1_axb_26 ));
    CascadeMux I__9668 (
            .O(N__43717),
            .I(N__43714));
    InMux I__9667 (
            .O(N__43714),
            .I(N__43711));
    LocalMux I__9666 (
            .O(N__43711),
            .I(N__43708));
    Odrv4 I__9665 (
            .O(N__43708),
            .I(\current_shift_inst.un4_control_input_1_axb_28 ));
    InMux I__9664 (
            .O(N__43705),
            .I(N__43702));
    LocalMux I__9663 (
            .O(N__43702),
            .I(N__43698));
    InMux I__9662 (
            .O(N__43701),
            .I(N__43695));
    Span4Mux_v I__9661 (
            .O(N__43698),
            .I(N__43689));
    LocalMux I__9660 (
            .O(N__43695),
            .I(N__43689));
    InMux I__9659 (
            .O(N__43694),
            .I(N__43686));
    Odrv4 I__9658 (
            .O(N__43689),
            .I(\current_shift_inst.un4_control_input1_26 ));
    LocalMux I__9657 (
            .O(N__43686),
            .I(\current_shift_inst.un4_control_input1_26 ));
    InMux I__9656 (
            .O(N__43681),
            .I(N__43678));
    LocalMux I__9655 (
            .O(N__43678),
            .I(N__43675));
    Odrv12 I__9654 (
            .O(N__43675),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ));
    InMux I__9653 (
            .O(N__43672),
            .I(N__43669));
    LocalMux I__9652 (
            .O(N__43669),
            .I(N__43666));
    Odrv12 I__9651 (
            .O(N__43666),
            .I(\current_shift_inst.un4_control_input_1_axb_29 ));
    InMux I__9650 (
            .O(N__43663),
            .I(N__43658));
    InMux I__9649 (
            .O(N__43662),
            .I(N__43654));
    InMux I__9648 (
            .O(N__43661),
            .I(N__43651));
    LocalMux I__9647 (
            .O(N__43658),
            .I(N__43648));
    InMux I__9646 (
            .O(N__43657),
            .I(N__43645));
    LocalMux I__9645 (
            .O(N__43654),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    LocalMux I__9644 (
            .O(N__43651),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    Odrv12 I__9643 (
            .O(N__43648),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    LocalMux I__9642 (
            .O(N__43645),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    InMux I__9641 (
            .O(N__43636),
            .I(N__43633));
    LocalMux I__9640 (
            .O(N__43633),
            .I(N__43629));
    InMux I__9639 (
            .O(N__43632),
            .I(N__43626));
    Span4Mux_v I__9638 (
            .O(N__43629),
            .I(N__43620));
    LocalMux I__9637 (
            .O(N__43626),
            .I(N__43620));
    InMux I__9636 (
            .O(N__43625),
            .I(N__43617));
    Span4Mux_h I__9635 (
            .O(N__43620),
            .I(N__43613));
    LocalMux I__9634 (
            .O(N__43617),
            .I(N__43609));
    InMux I__9633 (
            .O(N__43616),
            .I(N__43606));
    Span4Mux_h I__9632 (
            .O(N__43613),
            .I(N__43603));
    InMux I__9631 (
            .O(N__43612),
            .I(N__43600));
    Odrv4 I__9630 (
            .O(N__43609),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    LocalMux I__9629 (
            .O(N__43606),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    Odrv4 I__9628 (
            .O(N__43603),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    LocalMux I__9627 (
            .O(N__43600),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    InMux I__9626 (
            .O(N__43591),
            .I(N__43585));
    InMux I__9625 (
            .O(N__43590),
            .I(N__43582));
    CascadeMux I__9624 (
            .O(N__43589),
            .I(N__43579));
    CascadeMux I__9623 (
            .O(N__43588),
            .I(N__43576));
    LocalMux I__9622 (
            .O(N__43585),
            .I(N__43573));
    LocalMux I__9621 (
            .O(N__43582),
            .I(N__43570));
    InMux I__9620 (
            .O(N__43579),
            .I(N__43566));
    InMux I__9619 (
            .O(N__43576),
            .I(N__43563));
    Span12Mux_v I__9618 (
            .O(N__43573),
            .I(N__43560));
    Span4Mux_h I__9617 (
            .O(N__43570),
            .I(N__43557));
    InMux I__9616 (
            .O(N__43569),
            .I(N__43554));
    LocalMux I__9615 (
            .O(N__43566),
            .I(N__43551));
    LocalMux I__9614 (
            .O(N__43563),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    Odrv12 I__9613 (
            .O(N__43560),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    Odrv4 I__9612 (
            .O(N__43557),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    LocalMux I__9611 (
            .O(N__43554),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    Odrv4 I__9610 (
            .O(N__43551),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    CascadeMux I__9609 (
            .O(N__43540),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_ ));
    InMux I__9608 (
            .O(N__43537),
            .I(N__43532));
    CascadeMux I__9607 (
            .O(N__43536),
            .I(N__43529));
    InMux I__9606 (
            .O(N__43535),
            .I(N__43524));
    LocalMux I__9605 (
            .O(N__43532),
            .I(N__43521));
    InMux I__9604 (
            .O(N__43529),
            .I(N__43516));
    InMux I__9603 (
            .O(N__43528),
            .I(N__43516));
    InMux I__9602 (
            .O(N__43527),
            .I(N__43513));
    LocalMux I__9601 (
            .O(N__43524),
            .I(N__43508));
    Span12Mux_s7_v I__9600 (
            .O(N__43521),
            .I(N__43508));
    LocalMux I__9599 (
            .O(N__43516),
            .I(N__43505));
    LocalMux I__9598 (
            .O(N__43513),
            .I(N__43502));
    Odrv12 I__9597 (
            .O(N__43508),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    Odrv4 I__9596 (
            .O(N__43505),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    Odrv4 I__9595 (
            .O(N__43502),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    InMux I__9594 (
            .O(N__43495),
            .I(N__43492));
    LocalMux I__9593 (
            .O(N__43492),
            .I(N__43489));
    Odrv12 I__9592 (
            .O(N__43489),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_3 ));
    InMux I__9591 (
            .O(N__43486),
            .I(N__43483));
    LocalMux I__9590 (
            .O(N__43483),
            .I(N__43480));
    Odrv4 I__9589 (
            .O(N__43480),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ));
    CascadeMux I__9588 (
            .O(N__43477),
            .I(N__43474));
    InMux I__9587 (
            .O(N__43474),
            .I(N__43471));
    LocalMux I__9586 (
            .O(N__43471),
            .I(N__43465));
    InMux I__9585 (
            .O(N__43470),
            .I(N__43462));
    InMux I__9584 (
            .O(N__43469),
            .I(N__43459));
    InMux I__9583 (
            .O(N__43468),
            .I(N__43456));
    Span4Mux_h I__9582 (
            .O(N__43465),
            .I(N__43453));
    LocalMux I__9581 (
            .O(N__43462),
            .I(N__43447));
    LocalMux I__9580 (
            .O(N__43459),
            .I(N__43447));
    LocalMux I__9579 (
            .O(N__43456),
            .I(N__43442));
    Sp12to4 I__9578 (
            .O(N__43453),
            .I(N__43442));
    InMux I__9577 (
            .O(N__43452),
            .I(N__43439));
    Span12Mux_h I__9576 (
            .O(N__43447),
            .I(N__43436));
    Odrv12 I__9575 (
            .O(N__43442),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    LocalMux I__9574 (
            .O(N__43439),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    Odrv12 I__9573 (
            .O(N__43436),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    InMux I__9572 (
            .O(N__43429),
            .I(N__43426));
    LocalMux I__9571 (
            .O(N__43426),
            .I(N__43423));
    Span4Mux_v I__9570 (
            .O(N__43423),
            .I(N__43420));
    Odrv4 I__9569 (
            .O(N__43420),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ));
    InMux I__9568 (
            .O(N__43417),
            .I(N__43414));
    LocalMux I__9567 (
            .O(N__43414),
            .I(N__43411));
    Odrv4 I__9566 (
            .O(N__43411),
            .I(\current_shift_inst.un4_control_input_1_axb_21 ));
    InMux I__9565 (
            .O(N__43408),
            .I(N__43405));
    LocalMux I__9564 (
            .O(N__43405),
            .I(N__43402));
    Odrv4 I__9563 (
            .O(N__43402),
            .I(\current_shift_inst.un4_control_input_1_axb_22 ));
    InMux I__9562 (
            .O(N__43399),
            .I(N__43396));
    LocalMux I__9561 (
            .O(N__43396),
            .I(N__43393));
    Odrv4 I__9560 (
            .O(N__43393),
            .I(\current_shift_inst.un4_control_input_1_axb_17 ));
    InMux I__9559 (
            .O(N__43390),
            .I(N__43387));
    LocalMux I__9558 (
            .O(N__43387),
            .I(\current_shift_inst.un4_control_input_1_axb_25 ));
    InMux I__9557 (
            .O(N__43384),
            .I(N__43381));
    LocalMux I__9556 (
            .O(N__43381),
            .I(N__43378));
    Odrv4 I__9555 (
            .O(N__43378),
            .I(\current_shift_inst.un4_control_input_1_axb_20 ));
    InMux I__9554 (
            .O(N__43375),
            .I(N__43372));
    LocalMux I__9553 (
            .O(N__43372),
            .I(N__43368));
    InMux I__9552 (
            .O(N__43371),
            .I(N__43365));
    Span4Mux_v I__9551 (
            .O(N__43368),
            .I(N__43359));
    LocalMux I__9550 (
            .O(N__43365),
            .I(N__43359));
    InMux I__9549 (
            .O(N__43364),
            .I(N__43356));
    Odrv4 I__9548 (
            .O(N__43359),
            .I(\current_shift_inst.un4_control_input1_18 ));
    LocalMux I__9547 (
            .O(N__43356),
            .I(\current_shift_inst.un4_control_input1_18 ));
    InMux I__9546 (
            .O(N__43351),
            .I(N__43348));
    LocalMux I__9545 (
            .O(N__43348),
            .I(N__43345));
    Odrv12 I__9544 (
            .O(N__43345),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18 ));
    InMux I__9543 (
            .O(N__43342),
            .I(N__43339));
    LocalMux I__9542 (
            .O(N__43339),
            .I(N__43336));
    Odrv4 I__9541 (
            .O(N__43336),
            .I(\current_shift_inst.un4_control_input_1_axb_19 ));
    InMux I__9540 (
            .O(N__43333),
            .I(N__43330));
    LocalMux I__9539 (
            .O(N__43330),
            .I(N__43327));
    Odrv4 I__9538 (
            .O(N__43327),
            .I(\current_shift_inst.un4_control_input_1_axb_24 ));
    InMux I__9537 (
            .O(N__43324),
            .I(N__43321));
    LocalMux I__9536 (
            .O(N__43321),
            .I(N__43317));
    InMux I__9535 (
            .O(N__43320),
            .I(N__43314));
    Span4Mux_v I__9534 (
            .O(N__43317),
            .I(N__43308));
    LocalMux I__9533 (
            .O(N__43314),
            .I(N__43308));
    InMux I__9532 (
            .O(N__43313),
            .I(N__43305));
    Odrv4 I__9531 (
            .O(N__43308),
            .I(\current_shift_inst.un4_control_input1_28 ));
    LocalMux I__9530 (
            .O(N__43305),
            .I(\current_shift_inst.un4_control_input1_28 ));
    InMux I__9529 (
            .O(N__43300),
            .I(N__43297));
    LocalMux I__9528 (
            .O(N__43297),
            .I(N__43294));
    Odrv12 I__9527 (
            .O(N__43294),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ));
    InMux I__9526 (
            .O(N__43291),
            .I(bfn_17_18_0_));
    InMux I__9525 (
            .O(N__43288),
            .I(N__43284));
    InMux I__9524 (
            .O(N__43287),
            .I(N__43281));
    LocalMux I__9523 (
            .O(N__43284),
            .I(N__43277));
    LocalMux I__9522 (
            .O(N__43281),
            .I(N__43274));
    InMux I__9521 (
            .O(N__43280),
            .I(N__43271));
    Span4Mux_h I__9520 (
            .O(N__43277),
            .I(N__43268));
    Span4Mux_v I__9519 (
            .O(N__43274),
            .I(N__43263));
    LocalMux I__9518 (
            .O(N__43271),
            .I(N__43263));
    Odrv4 I__9517 (
            .O(N__43268),
            .I(\current_shift_inst.un4_control_input1_27 ));
    Odrv4 I__9516 (
            .O(N__43263),
            .I(\current_shift_inst.un4_control_input1_27 ));
    InMux I__9515 (
            .O(N__43258),
            .I(\current_shift_inst.un4_control_input_1_cry_25 ));
    InMux I__9514 (
            .O(N__43255),
            .I(\current_shift_inst.un4_control_input_1_cry_26 ));
    InMux I__9513 (
            .O(N__43252),
            .I(N__43249));
    LocalMux I__9512 (
            .O(N__43249),
            .I(N__43246));
    Span4Mux_v I__9511 (
            .O(N__43246),
            .I(N__43243));
    Span4Mux_h I__9510 (
            .O(N__43243),
            .I(N__43238));
    InMux I__9509 (
            .O(N__43242),
            .I(N__43233));
    InMux I__9508 (
            .O(N__43241),
            .I(N__43233));
    Odrv4 I__9507 (
            .O(N__43238),
            .I(\current_shift_inst.un4_control_input1_29 ));
    LocalMux I__9506 (
            .O(N__43233),
            .I(\current_shift_inst.un4_control_input1_29 ));
    InMux I__9505 (
            .O(N__43228),
            .I(\current_shift_inst.un4_control_input_1_cry_27 ));
    InMux I__9504 (
            .O(N__43225),
            .I(N__43221));
    InMux I__9503 (
            .O(N__43224),
            .I(N__43218));
    LocalMux I__9502 (
            .O(N__43221),
            .I(N__43212));
    LocalMux I__9501 (
            .O(N__43218),
            .I(N__43212));
    InMux I__9500 (
            .O(N__43217),
            .I(N__43209));
    Odrv4 I__9499 (
            .O(N__43212),
            .I(\current_shift_inst.un4_control_input1_30 ));
    LocalMux I__9498 (
            .O(N__43209),
            .I(\current_shift_inst.un4_control_input1_30 ));
    InMux I__9497 (
            .O(N__43204),
            .I(\current_shift_inst.un4_control_input_1_cry_28 ));
    InMux I__9496 (
            .O(N__43201),
            .I(\current_shift_inst.un4_control_input1_31 ));
    InMux I__9495 (
            .O(N__43198),
            .I(N__43195));
    LocalMux I__9494 (
            .O(N__43195),
            .I(N__43192));
    Odrv4 I__9493 (
            .O(N__43192),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    CascadeMux I__9492 (
            .O(N__43189),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO_cascade_ ));
    InMux I__9491 (
            .O(N__43186),
            .I(N__43183));
    LocalMux I__9490 (
            .O(N__43183),
            .I(N__43180));
    Odrv4 I__9489 (
            .O(N__43180),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ));
    InMux I__9488 (
            .O(N__43177),
            .I(N__43174));
    LocalMux I__9487 (
            .O(N__43174),
            .I(\current_shift_inst.un4_control_input_1_axb_18 ));
    InMux I__9486 (
            .O(N__43171),
            .I(N__43167));
    InMux I__9485 (
            .O(N__43170),
            .I(N__43164));
    LocalMux I__9484 (
            .O(N__43167),
            .I(N__43158));
    LocalMux I__9483 (
            .O(N__43164),
            .I(N__43158));
    InMux I__9482 (
            .O(N__43163),
            .I(N__43155));
    Odrv4 I__9481 (
            .O(N__43158),
            .I(\current_shift_inst.un4_control_input1_24 ));
    LocalMux I__9480 (
            .O(N__43155),
            .I(\current_shift_inst.un4_control_input1_24 ));
    CascadeMux I__9479 (
            .O(N__43150),
            .I(N__43147));
    InMux I__9478 (
            .O(N__43147),
            .I(N__43144));
    LocalMux I__9477 (
            .O(N__43144),
            .I(N__43141));
    Odrv12 I__9476 (
            .O(N__43141),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ));
    InMux I__9475 (
            .O(N__43138),
            .I(bfn_17_17_0_));
    InMux I__9474 (
            .O(N__43135),
            .I(\current_shift_inst.un4_control_input_1_cry_17 ));
    InMux I__9473 (
            .O(N__43132),
            .I(N__43129));
    LocalMux I__9472 (
            .O(N__43129),
            .I(N__43124));
    InMux I__9471 (
            .O(N__43128),
            .I(N__43119));
    InMux I__9470 (
            .O(N__43127),
            .I(N__43119));
    Odrv4 I__9469 (
            .O(N__43124),
            .I(\current_shift_inst.un4_control_input1_20 ));
    LocalMux I__9468 (
            .O(N__43119),
            .I(\current_shift_inst.un4_control_input1_20 ));
    InMux I__9467 (
            .O(N__43114),
            .I(\current_shift_inst.un4_control_input_1_cry_18 ));
    InMux I__9466 (
            .O(N__43111),
            .I(N__43108));
    LocalMux I__9465 (
            .O(N__43108),
            .I(N__43103));
    InMux I__9464 (
            .O(N__43107),
            .I(N__43098));
    InMux I__9463 (
            .O(N__43106),
            .I(N__43098));
    Odrv4 I__9462 (
            .O(N__43103),
            .I(\current_shift_inst.un4_control_input1_21 ));
    LocalMux I__9461 (
            .O(N__43098),
            .I(\current_shift_inst.un4_control_input1_21 ));
    InMux I__9460 (
            .O(N__43093),
            .I(\current_shift_inst.un4_control_input_1_cry_19 ));
    InMux I__9459 (
            .O(N__43090),
            .I(N__43086));
    InMux I__9458 (
            .O(N__43089),
            .I(N__43083));
    LocalMux I__9457 (
            .O(N__43086),
            .I(N__43080));
    LocalMux I__9456 (
            .O(N__43083),
            .I(N__43077));
    Span4Mux_v I__9455 (
            .O(N__43080),
            .I(N__43071));
    Span4Mux_h I__9454 (
            .O(N__43077),
            .I(N__43071));
    InMux I__9453 (
            .O(N__43076),
            .I(N__43068));
    Odrv4 I__9452 (
            .O(N__43071),
            .I(\current_shift_inst.un4_control_input1_22 ));
    LocalMux I__9451 (
            .O(N__43068),
            .I(\current_shift_inst.un4_control_input1_22 ));
    InMux I__9450 (
            .O(N__43063),
            .I(\current_shift_inst.un4_control_input_1_cry_20 ));
    InMux I__9449 (
            .O(N__43060),
            .I(N__43057));
    LocalMux I__9448 (
            .O(N__43057),
            .I(N__43054));
    Span4Mux_v I__9447 (
            .O(N__43054),
            .I(N__43050));
    InMux I__9446 (
            .O(N__43053),
            .I(N__43047));
    Span4Mux_h I__9445 (
            .O(N__43050),
            .I(N__43042));
    LocalMux I__9444 (
            .O(N__43047),
            .I(N__43042));
    Span4Mux_v I__9443 (
            .O(N__43042),
            .I(N__43038));
    InMux I__9442 (
            .O(N__43041),
            .I(N__43035));
    Odrv4 I__9441 (
            .O(N__43038),
            .I(\current_shift_inst.un4_control_input1_23 ));
    LocalMux I__9440 (
            .O(N__43035),
            .I(\current_shift_inst.un4_control_input1_23 ));
    InMux I__9439 (
            .O(N__43030),
            .I(\current_shift_inst.un4_control_input_1_cry_21 ));
    InMux I__9438 (
            .O(N__43027),
            .I(\current_shift_inst.un4_control_input_1_cry_22 ));
    InMux I__9437 (
            .O(N__43024),
            .I(N__43021));
    LocalMux I__9436 (
            .O(N__43021),
            .I(N__43018));
    Span4Mux_h I__9435 (
            .O(N__43018),
            .I(N__43013));
    InMux I__9434 (
            .O(N__43017),
            .I(N__43008));
    InMux I__9433 (
            .O(N__43016),
            .I(N__43008));
    Odrv4 I__9432 (
            .O(N__43013),
            .I(\current_shift_inst.un4_control_input1_25 ));
    LocalMux I__9431 (
            .O(N__43008),
            .I(\current_shift_inst.un4_control_input1_25 ));
    InMux I__9430 (
            .O(N__43003),
            .I(\current_shift_inst.un4_control_input_1_cry_23 ));
    InMux I__9429 (
            .O(N__43000),
            .I(N__42996));
    InMux I__9428 (
            .O(N__42999),
            .I(N__42993));
    LocalMux I__9427 (
            .O(N__42996),
            .I(N__42990));
    LocalMux I__9426 (
            .O(N__42993),
            .I(N__42987));
    Span4Mux_v I__9425 (
            .O(N__42990),
            .I(N__42981));
    Span4Mux_h I__9424 (
            .O(N__42987),
            .I(N__42981));
    InMux I__9423 (
            .O(N__42986),
            .I(N__42978));
    Odrv4 I__9422 (
            .O(N__42981),
            .I(\current_shift_inst.un4_control_input1_9 ));
    LocalMux I__9421 (
            .O(N__42978),
            .I(\current_shift_inst.un4_control_input1_9 ));
    InMux I__9420 (
            .O(N__42973),
            .I(\current_shift_inst.un4_control_input_1_cry_7 ));
    InMux I__9419 (
            .O(N__42970),
            .I(N__42967));
    LocalMux I__9418 (
            .O(N__42967),
            .I(N__42964));
    Span4Mux_h I__9417 (
            .O(N__42964),
            .I(N__42961));
    Span4Mux_h I__9416 (
            .O(N__42961),
            .I(N__42956));
    InMux I__9415 (
            .O(N__42960),
            .I(N__42953));
    InMux I__9414 (
            .O(N__42959),
            .I(N__42950));
    Odrv4 I__9413 (
            .O(N__42956),
            .I(\current_shift_inst.un4_control_input1_10 ));
    LocalMux I__9412 (
            .O(N__42953),
            .I(\current_shift_inst.un4_control_input1_10 ));
    LocalMux I__9411 (
            .O(N__42950),
            .I(\current_shift_inst.un4_control_input1_10 ));
    InMux I__9410 (
            .O(N__42943),
            .I(bfn_17_16_0_));
    InMux I__9409 (
            .O(N__42940),
            .I(N__42937));
    LocalMux I__9408 (
            .O(N__42937),
            .I(N__42933));
    InMux I__9407 (
            .O(N__42936),
            .I(N__42930));
    Span4Mux_v I__9406 (
            .O(N__42933),
            .I(N__42926));
    LocalMux I__9405 (
            .O(N__42930),
            .I(N__42923));
    InMux I__9404 (
            .O(N__42929),
            .I(N__42920));
    Odrv4 I__9403 (
            .O(N__42926),
            .I(\current_shift_inst.un4_control_input1_11 ));
    Odrv12 I__9402 (
            .O(N__42923),
            .I(\current_shift_inst.un4_control_input1_11 ));
    LocalMux I__9401 (
            .O(N__42920),
            .I(\current_shift_inst.un4_control_input1_11 ));
    InMux I__9400 (
            .O(N__42913),
            .I(\current_shift_inst.un4_control_input_1_cry_9 ));
    InMux I__9399 (
            .O(N__42910),
            .I(\current_shift_inst.un4_control_input_1_cry_10 ));
    InMux I__9398 (
            .O(N__42907),
            .I(N__42904));
    LocalMux I__9397 (
            .O(N__42904),
            .I(N__42901));
    Span4Mux_h I__9396 (
            .O(N__42901),
            .I(N__42896));
    InMux I__9395 (
            .O(N__42900),
            .I(N__42893));
    InMux I__9394 (
            .O(N__42899),
            .I(N__42890));
    Odrv4 I__9393 (
            .O(N__42896),
            .I(\current_shift_inst.un4_control_input1_13 ));
    LocalMux I__9392 (
            .O(N__42893),
            .I(\current_shift_inst.un4_control_input1_13 ));
    LocalMux I__9391 (
            .O(N__42890),
            .I(\current_shift_inst.un4_control_input1_13 ));
    InMux I__9390 (
            .O(N__42883),
            .I(\current_shift_inst.un4_control_input_1_cry_11 ));
    InMux I__9389 (
            .O(N__42880),
            .I(N__42877));
    LocalMux I__9388 (
            .O(N__42877),
            .I(N__42873));
    InMux I__9387 (
            .O(N__42876),
            .I(N__42870));
    Span4Mux_h I__9386 (
            .O(N__42873),
            .I(N__42866));
    LocalMux I__9385 (
            .O(N__42870),
            .I(N__42863));
    InMux I__9384 (
            .O(N__42869),
            .I(N__42860));
    Odrv4 I__9383 (
            .O(N__42866),
            .I(\current_shift_inst.un4_control_input1_14 ));
    Odrv4 I__9382 (
            .O(N__42863),
            .I(\current_shift_inst.un4_control_input1_14 ));
    LocalMux I__9381 (
            .O(N__42860),
            .I(\current_shift_inst.un4_control_input1_14 ));
    InMux I__9380 (
            .O(N__42853),
            .I(\current_shift_inst.un4_control_input_1_cry_12 ));
    InMux I__9379 (
            .O(N__42850),
            .I(N__42847));
    LocalMux I__9378 (
            .O(N__42847),
            .I(N__42843));
    InMux I__9377 (
            .O(N__42846),
            .I(N__42840));
    Span4Mux_v I__9376 (
            .O(N__42843),
            .I(N__42836));
    LocalMux I__9375 (
            .O(N__42840),
            .I(N__42833));
    InMux I__9374 (
            .O(N__42839),
            .I(N__42830));
    Odrv4 I__9373 (
            .O(N__42836),
            .I(\current_shift_inst.un4_control_input1_15 ));
    Odrv12 I__9372 (
            .O(N__42833),
            .I(\current_shift_inst.un4_control_input1_15 ));
    LocalMux I__9371 (
            .O(N__42830),
            .I(\current_shift_inst.un4_control_input1_15 ));
    InMux I__9370 (
            .O(N__42823),
            .I(\current_shift_inst.un4_control_input_1_cry_13 ));
    InMux I__9369 (
            .O(N__42820),
            .I(N__42816));
    InMux I__9368 (
            .O(N__42819),
            .I(N__42813));
    LocalMux I__9367 (
            .O(N__42816),
            .I(N__42810));
    LocalMux I__9366 (
            .O(N__42813),
            .I(N__42807));
    Span4Mux_v I__9365 (
            .O(N__42810),
            .I(N__42801));
    Span4Mux_h I__9364 (
            .O(N__42807),
            .I(N__42801));
    InMux I__9363 (
            .O(N__42806),
            .I(N__42798));
    Odrv4 I__9362 (
            .O(N__42801),
            .I(\current_shift_inst.un4_control_input1_16 ));
    LocalMux I__9361 (
            .O(N__42798),
            .I(\current_shift_inst.un4_control_input1_16 ));
    InMux I__9360 (
            .O(N__42793),
            .I(\current_shift_inst.un4_control_input_1_cry_14 ));
    InMux I__9359 (
            .O(N__42790),
            .I(\current_shift_inst.un4_control_input_1_cry_15 ));
    InMux I__9358 (
            .O(N__42787),
            .I(N__42749));
    InMux I__9357 (
            .O(N__42786),
            .I(N__42749));
    InMux I__9356 (
            .O(N__42785),
            .I(N__42749));
    InMux I__9355 (
            .O(N__42784),
            .I(N__42749));
    InMux I__9354 (
            .O(N__42783),
            .I(N__42740));
    InMux I__9353 (
            .O(N__42782),
            .I(N__42740));
    InMux I__9352 (
            .O(N__42781),
            .I(N__42740));
    InMux I__9351 (
            .O(N__42780),
            .I(N__42740));
    InMux I__9350 (
            .O(N__42779),
            .I(N__42731));
    InMux I__9349 (
            .O(N__42778),
            .I(N__42731));
    InMux I__9348 (
            .O(N__42777),
            .I(N__42731));
    InMux I__9347 (
            .O(N__42776),
            .I(N__42731));
    InMux I__9346 (
            .O(N__42775),
            .I(N__42722));
    InMux I__9345 (
            .O(N__42774),
            .I(N__42722));
    InMux I__9344 (
            .O(N__42773),
            .I(N__42722));
    InMux I__9343 (
            .O(N__42772),
            .I(N__42722));
    InMux I__9342 (
            .O(N__42771),
            .I(N__42713));
    InMux I__9341 (
            .O(N__42770),
            .I(N__42713));
    InMux I__9340 (
            .O(N__42769),
            .I(N__42713));
    InMux I__9339 (
            .O(N__42768),
            .I(N__42713));
    InMux I__9338 (
            .O(N__42767),
            .I(N__42704));
    InMux I__9337 (
            .O(N__42766),
            .I(N__42704));
    InMux I__9336 (
            .O(N__42765),
            .I(N__42704));
    InMux I__9335 (
            .O(N__42764),
            .I(N__42704));
    InMux I__9334 (
            .O(N__42763),
            .I(N__42699));
    InMux I__9333 (
            .O(N__42762),
            .I(N__42699));
    InMux I__9332 (
            .O(N__42761),
            .I(N__42690));
    InMux I__9331 (
            .O(N__42760),
            .I(N__42690));
    InMux I__9330 (
            .O(N__42759),
            .I(N__42690));
    InMux I__9329 (
            .O(N__42758),
            .I(N__42690));
    LocalMux I__9328 (
            .O(N__42749),
            .I(N__42687));
    LocalMux I__9327 (
            .O(N__42740),
            .I(N__42680));
    LocalMux I__9326 (
            .O(N__42731),
            .I(N__42680));
    LocalMux I__9325 (
            .O(N__42722),
            .I(N__42680));
    LocalMux I__9324 (
            .O(N__42713),
            .I(N__42671));
    LocalMux I__9323 (
            .O(N__42704),
            .I(N__42671));
    LocalMux I__9322 (
            .O(N__42699),
            .I(N__42671));
    LocalMux I__9321 (
            .O(N__42690),
            .I(N__42671));
    Span4Mux_v I__9320 (
            .O(N__42687),
            .I(N__42664));
    Span4Mux_v I__9319 (
            .O(N__42680),
            .I(N__42664));
    Span4Mux_v I__9318 (
            .O(N__42671),
            .I(N__42664));
    Span4Mux_v I__9317 (
            .O(N__42664),
            .I(N__42661));
    Odrv4 I__9316 (
            .O(N__42661),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    InMux I__9315 (
            .O(N__42658),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ));
    InMux I__9314 (
            .O(N__42655),
            .I(N__42651));
    InMux I__9313 (
            .O(N__42654),
            .I(N__42648));
    LocalMux I__9312 (
            .O(N__42651),
            .I(N__42645));
    LocalMux I__9311 (
            .O(N__42648),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    Odrv4 I__9310 (
            .O(N__42645),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    CEMux I__9309 (
            .O(N__42640),
            .I(N__42635));
    CEMux I__9308 (
            .O(N__42639),
            .I(N__42632));
    CEMux I__9307 (
            .O(N__42638),
            .I(N__42629));
    LocalMux I__9306 (
            .O(N__42635),
            .I(N__42624));
    LocalMux I__9305 (
            .O(N__42632),
            .I(N__42624));
    LocalMux I__9304 (
            .O(N__42629),
            .I(N__42620));
    Span4Mux_v I__9303 (
            .O(N__42624),
            .I(N__42617));
    CEMux I__9302 (
            .O(N__42623),
            .I(N__42614));
    Span4Mux_v I__9301 (
            .O(N__42620),
            .I(N__42607));
    Span4Mux_h I__9300 (
            .O(N__42617),
            .I(N__42607));
    LocalMux I__9299 (
            .O(N__42614),
            .I(N__42607));
    Span4Mux_v I__9298 (
            .O(N__42607),
            .I(N__42604));
    Odrv4 I__9297 (
            .O(N__42604),
            .I(\delay_measurement_inst.delay_tr_timer.N_305_i ));
    InMux I__9296 (
            .O(N__42601),
            .I(N__42598));
    LocalMux I__9295 (
            .O(N__42598),
            .I(\current_shift_inst.un4_control_input_1_axb_1 ));
    CascadeMux I__9294 (
            .O(N__42595),
            .I(N__42592));
    InMux I__9293 (
            .O(N__42592),
            .I(N__42583));
    InMux I__9292 (
            .O(N__42591),
            .I(N__42583));
    InMux I__9291 (
            .O(N__42590),
            .I(N__42583));
    LocalMux I__9290 (
            .O(N__42583),
            .I(\current_shift_inst.un4_control_input1_2 ));
    InMux I__9289 (
            .O(N__42580),
            .I(\current_shift_inst.un4_control_input_1_cry_1 ));
    InMux I__9288 (
            .O(N__42577),
            .I(N__42568));
    InMux I__9287 (
            .O(N__42576),
            .I(N__42568));
    InMux I__9286 (
            .O(N__42575),
            .I(N__42568));
    LocalMux I__9285 (
            .O(N__42568),
            .I(\current_shift_inst.un4_control_input1_4 ));
    InMux I__9284 (
            .O(N__42565),
            .I(\current_shift_inst.un4_control_input_1_cry_2 ));
    InMux I__9283 (
            .O(N__42562),
            .I(\current_shift_inst.un4_control_input_1_cry_3 ));
    InMux I__9282 (
            .O(N__42559),
            .I(N__42555));
    InMux I__9281 (
            .O(N__42558),
            .I(N__42552));
    LocalMux I__9280 (
            .O(N__42555),
            .I(N__42548));
    LocalMux I__9279 (
            .O(N__42552),
            .I(N__42545));
    InMux I__9278 (
            .O(N__42551),
            .I(N__42542));
    Odrv4 I__9277 (
            .O(N__42548),
            .I(\current_shift_inst.un4_control_input1_6 ));
    Odrv12 I__9276 (
            .O(N__42545),
            .I(\current_shift_inst.un4_control_input1_6 ));
    LocalMux I__9275 (
            .O(N__42542),
            .I(\current_shift_inst.un4_control_input1_6 ));
    InMux I__9274 (
            .O(N__42535),
            .I(\current_shift_inst.un4_control_input_1_cry_4 ));
    InMux I__9273 (
            .O(N__42532),
            .I(\current_shift_inst.un4_control_input_1_cry_5 ));
    InMux I__9272 (
            .O(N__42529),
            .I(\current_shift_inst.un4_control_input_1_cry_6 ));
    InMux I__9271 (
            .O(N__42526),
            .I(N__42519));
    InMux I__9270 (
            .O(N__42525),
            .I(N__42519));
    InMux I__9269 (
            .O(N__42524),
            .I(N__42516));
    LocalMux I__9268 (
            .O(N__42519),
            .I(N__42513));
    LocalMux I__9267 (
            .O(N__42516),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    Odrv4 I__9266 (
            .O(N__42513),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    InMux I__9265 (
            .O(N__42508),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ));
    InMux I__9264 (
            .O(N__42505),
            .I(N__42498));
    InMux I__9263 (
            .O(N__42504),
            .I(N__42498));
    InMux I__9262 (
            .O(N__42503),
            .I(N__42495));
    LocalMux I__9261 (
            .O(N__42498),
            .I(N__42492));
    LocalMux I__9260 (
            .O(N__42495),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    Odrv12 I__9259 (
            .O(N__42492),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    InMux I__9258 (
            .O(N__42487),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ));
    CascadeMux I__9257 (
            .O(N__42484),
            .I(N__42480));
    CascadeMux I__9256 (
            .O(N__42483),
            .I(N__42477));
    InMux I__9255 (
            .O(N__42480),
            .I(N__42471));
    InMux I__9254 (
            .O(N__42477),
            .I(N__42471));
    InMux I__9253 (
            .O(N__42476),
            .I(N__42468));
    LocalMux I__9252 (
            .O(N__42471),
            .I(N__42465));
    LocalMux I__9251 (
            .O(N__42468),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    Odrv12 I__9250 (
            .O(N__42465),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    InMux I__9249 (
            .O(N__42460),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ));
    CascadeMux I__9248 (
            .O(N__42457),
            .I(N__42453));
    CascadeMux I__9247 (
            .O(N__42456),
            .I(N__42450));
    InMux I__9246 (
            .O(N__42453),
            .I(N__42444));
    InMux I__9245 (
            .O(N__42450),
            .I(N__42444));
    InMux I__9244 (
            .O(N__42449),
            .I(N__42441));
    LocalMux I__9243 (
            .O(N__42444),
            .I(N__42438));
    LocalMux I__9242 (
            .O(N__42441),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    Odrv12 I__9241 (
            .O(N__42438),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    InMux I__9240 (
            .O(N__42433),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ));
    InMux I__9239 (
            .O(N__42430),
            .I(N__42426));
    InMux I__9238 (
            .O(N__42429),
            .I(N__42422));
    LocalMux I__9237 (
            .O(N__42426),
            .I(N__42419));
    InMux I__9236 (
            .O(N__42425),
            .I(N__42416));
    LocalMux I__9235 (
            .O(N__42422),
            .I(N__42411));
    Span4Mux_v I__9234 (
            .O(N__42419),
            .I(N__42411));
    LocalMux I__9233 (
            .O(N__42416),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    Odrv4 I__9232 (
            .O(N__42411),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    InMux I__9231 (
            .O(N__42406),
            .I(bfn_17_14_0_));
    InMux I__9230 (
            .O(N__42403),
            .I(N__42399));
    InMux I__9229 (
            .O(N__42402),
            .I(N__42396));
    LocalMux I__9228 (
            .O(N__42399),
            .I(N__42393));
    LocalMux I__9227 (
            .O(N__42396),
            .I(N__42387));
    Span4Mux_v I__9226 (
            .O(N__42393),
            .I(N__42387));
    InMux I__9225 (
            .O(N__42392),
            .I(N__42384));
    Span4Mux_h I__9224 (
            .O(N__42387),
            .I(N__42381));
    LocalMux I__9223 (
            .O(N__42384),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    Odrv4 I__9222 (
            .O(N__42381),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    InMux I__9221 (
            .O(N__42376),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ));
    CascadeMux I__9220 (
            .O(N__42373),
            .I(N__42369));
    CascadeMux I__9219 (
            .O(N__42372),
            .I(N__42366));
    InMux I__9218 (
            .O(N__42369),
            .I(N__42360));
    InMux I__9217 (
            .O(N__42366),
            .I(N__42360));
    InMux I__9216 (
            .O(N__42365),
            .I(N__42357));
    LocalMux I__9215 (
            .O(N__42360),
            .I(N__42354));
    LocalMux I__9214 (
            .O(N__42357),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    Odrv4 I__9213 (
            .O(N__42354),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    InMux I__9212 (
            .O(N__42349),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ));
    CascadeMux I__9211 (
            .O(N__42346),
            .I(N__42342));
    CascadeMux I__9210 (
            .O(N__42345),
            .I(N__42339));
    InMux I__9209 (
            .O(N__42342),
            .I(N__42333));
    InMux I__9208 (
            .O(N__42339),
            .I(N__42333));
    InMux I__9207 (
            .O(N__42338),
            .I(N__42330));
    LocalMux I__9206 (
            .O(N__42333),
            .I(N__42327));
    LocalMux I__9205 (
            .O(N__42330),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    Odrv4 I__9204 (
            .O(N__42327),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    InMux I__9203 (
            .O(N__42322),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ));
    InMux I__9202 (
            .O(N__42319),
            .I(N__42315));
    InMux I__9201 (
            .O(N__42318),
            .I(N__42312));
    LocalMux I__9200 (
            .O(N__42315),
            .I(N__42309));
    LocalMux I__9199 (
            .O(N__42312),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    Odrv12 I__9198 (
            .O(N__42309),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    InMux I__9197 (
            .O(N__42304),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ));
    InMux I__9196 (
            .O(N__42301),
            .I(N__42295));
    InMux I__9195 (
            .O(N__42300),
            .I(N__42295));
    LocalMux I__9194 (
            .O(N__42295),
            .I(N__42291));
    InMux I__9193 (
            .O(N__42294),
            .I(N__42288));
    Span4Mux_h I__9192 (
            .O(N__42291),
            .I(N__42285));
    LocalMux I__9191 (
            .O(N__42288),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    Odrv4 I__9190 (
            .O(N__42285),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    InMux I__9189 (
            .O(N__42280),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ));
    InMux I__9188 (
            .O(N__42277),
            .I(N__42270));
    InMux I__9187 (
            .O(N__42276),
            .I(N__42270));
    InMux I__9186 (
            .O(N__42275),
            .I(N__42267));
    LocalMux I__9185 (
            .O(N__42270),
            .I(N__42264));
    LocalMux I__9184 (
            .O(N__42267),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    Odrv4 I__9183 (
            .O(N__42264),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    InMux I__9182 (
            .O(N__42259),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ));
    CascadeMux I__9181 (
            .O(N__42256),
            .I(N__42252));
    CascadeMux I__9180 (
            .O(N__42255),
            .I(N__42249));
    InMux I__9179 (
            .O(N__42252),
            .I(N__42243));
    InMux I__9178 (
            .O(N__42249),
            .I(N__42243));
    InMux I__9177 (
            .O(N__42248),
            .I(N__42240));
    LocalMux I__9176 (
            .O(N__42243),
            .I(N__42237));
    LocalMux I__9175 (
            .O(N__42240),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    Odrv12 I__9174 (
            .O(N__42237),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    InMux I__9173 (
            .O(N__42232),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ));
    CascadeMux I__9172 (
            .O(N__42229),
            .I(N__42225));
    CascadeMux I__9171 (
            .O(N__42228),
            .I(N__42222));
    InMux I__9170 (
            .O(N__42225),
            .I(N__42216));
    InMux I__9169 (
            .O(N__42222),
            .I(N__42216));
    InMux I__9168 (
            .O(N__42221),
            .I(N__42213));
    LocalMux I__9167 (
            .O(N__42216),
            .I(N__42210));
    LocalMux I__9166 (
            .O(N__42213),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    Odrv12 I__9165 (
            .O(N__42210),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    InMux I__9164 (
            .O(N__42205),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ));
    InMux I__9163 (
            .O(N__42202),
            .I(N__42198));
    InMux I__9162 (
            .O(N__42201),
            .I(N__42195));
    LocalMux I__9161 (
            .O(N__42198),
            .I(N__42192));
    LocalMux I__9160 (
            .O(N__42195),
            .I(N__42186));
    Span4Mux_v I__9159 (
            .O(N__42192),
            .I(N__42186));
    InMux I__9158 (
            .O(N__42191),
            .I(N__42183));
    Span4Mux_h I__9157 (
            .O(N__42186),
            .I(N__42180));
    LocalMux I__9156 (
            .O(N__42183),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    Odrv4 I__9155 (
            .O(N__42180),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    InMux I__9154 (
            .O(N__42175),
            .I(bfn_17_13_0_));
    InMux I__9153 (
            .O(N__42172),
            .I(N__42168));
    InMux I__9152 (
            .O(N__42171),
            .I(N__42164));
    LocalMux I__9151 (
            .O(N__42168),
            .I(N__42161));
    InMux I__9150 (
            .O(N__42167),
            .I(N__42158));
    LocalMux I__9149 (
            .O(N__42164),
            .I(N__42153));
    Span4Mux_v I__9148 (
            .O(N__42161),
            .I(N__42153));
    LocalMux I__9147 (
            .O(N__42158),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    Odrv4 I__9146 (
            .O(N__42153),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    InMux I__9145 (
            .O(N__42148),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ));
    CascadeMux I__9144 (
            .O(N__42145),
            .I(N__42141));
    CascadeMux I__9143 (
            .O(N__42144),
            .I(N__42138));
    InMux I__9142 (
            .O(N__42141),
            .I(N__42132));
    InMux I__9141 (
            .O(N__42138),
            .I(N__42132));
    InMux I__9140 (
            .O(N__42137),
            .I(N__42129));
    LocalMux I__9139 (
            .O(N__42132),
            .I(N__42126));
    LocalMux I__9138 (
            .O(N__42129),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    Odrv4 I__9137 (
            .O(N__42126),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    InMux I__9136 (
            .O(N__42121),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ));
    CascadeMux I__9135 (
            .O(N__42118),
            .I(N__42114));
    CascadeMux I__9134 (
            .O(N__42117),
            .I(N__42111));
    InMux I__9133 (
            .O(N__42114),
            .I(N__42105));
    InMux I__9132 (
            .O(N__42111),
            .I(N__42105));
    InMux I__9131 (
            .O(N__42110),
            .I(N__42102));
    LocalMux I__9130 (
            .O(N__42105),
            .I(N__42099));
    LocalMux I__9129 (
            .O(N__42102),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    Odrv4 I__9128 (
            .O(N__42099),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    InMux I__9127 (
            .O(N__42094),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ));
    CascadeMux I__9126 (
            .O(N__42091),
            .I(N__42087));
    CascadeMux I__9125 (
            .O(N__42090),
            .I(N__42084));
    InMux I__9124 (
            .O(N__42087),
            .I(N__42078));
    InMux I__9123 (
            .O(N__42084),
            .I(N__42078));
    InMux I__9122 (
            .O(N__42083),
            .I(N__42075));
    LocalMux I__9121 (
            .O(N__42078),
            .I(N__42072));
    LocalMux I__9120 (
            .O(N__42075),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    Odrv12 I__9119 (
            .O(N__42072),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    InMux I__9118 (
            .O(N__42067),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ));
    InMux I__9117 (
            .O(N__42064),
            .I(N__42057));
    InMux I__9116 (
            .O(N__42063),
            .I(N__42057));
    InMux I__9115 (
            .O(N__42062),
            .I(N__42054));
    LocalMux I__9114 (
            .O(N__42057),
            .I(N__42051));
    LocalMux I__9113 (
            .O(N__42054),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    Odrv12 I__9112 (
            .O(N__42051),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    InMux I__9111 (
            .O(N__42046),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ));
    InMux I__9110 (
            .O(N__42043),
            .I(N__42037));
    InMux I__9109 (
            .O(N__42042),
            .I(N__42037));
    LocalMux I__9108 (
            .O(N__42037),
            .I(N__42033));
    InMux I__9107 (
            .O(N__42036),
            .I(N__42030));
    Span4Mux_h I__9106 (
            .O(N__42033),
            .I(N__42027));
    LocalMux I__9105 (
            .O(N__42030),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    Odrv4 I__9104 (
            .O(N__42027),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    InMux I__9103 (
            .O(N__42022),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ));
    CascadeMux I__9102 (
            .O(N__42019),
            .I(N__42015));
    CascadeMux I__9101 (
            .O(N__42018),
            .I(N__42012));
    InMux I__9100 (
            .O(N__42015),
            .I(N__42006));
    InMux I__9099 (
            .O(N__42012),
            .I(N__42006));
    InMux I__9098 (
            .O(N__42011),
            .I(N__42003));
    LocalMux I__9097 (
            .O(N__42006),
            .I(N__42000));
    LocalMux I__9096 (
            .O(N__42003),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    Odrv12 I__9095 (
            .O(N__42000),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    InMux I__9094 (
            .O(N__41995),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ));
    CascadeMux I__9093 (
            .O(N__41992),
            .I(N__41988));
    CascadeMux I__9092 (
            .O(N__41991),
            .I(N__41985));
    InMux I__9091 (
            .O(N__41988),
            .I(N__41979));
    InMux I__9090 (
            .O(N__41985),
            .I(N__41979));
    InMux I__9089 (
            .O(N__41984),
            .I(N__41976));
    LocalMux I__9088 (
            .O(N__41979),
            .I(N__41973));
    LocalMux I__9087 (
            .O(N__41976),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    Odrv4 I__9086 (
            .O(N__41973),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    InMux I__9085 (
            .O(N__41968),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ));
    InMux I__9084 (
            .O(N__41965),
            .I(N__41961));
    InMux I__9083 (
            .O(N__41964),
            .I(N__41957));
    LocalMux I__9082 (
            .O(N__41961),
            .I(N__41954));
    InMux I__9081 (
            .O(N__41960),
            .I(N__41951));
    LocalMux I__9080 (
            .O(N__41957),
            .I(N__41946));
    Span4Mux_v I__9079 (
            .O(N__41954),
            .I(N__41946));
    LocalMux I__9078 (
            .O(N__41951),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    Odrv4 I__9077 (
            .O(N__41946),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    InMux I__9076 (
            .O(N__41941),
            .I(bfn_17_12_0_));
    InMux I__9075 (
            .O(N__41938),
            .I(N__41934));
    InMux I__9074 (
            .O(N__41937),
            .I(N__41931));
    LocalMux I__9073 (
            .O(N__41934),
            .I(N__41928));
    LocalMux I__9072 (
            .O(N__41931),
            .I(N__41922));
    Span4Mux_v I__9071 (
            .O(N__41928),
            .I(N__41922));
    InMux I__9070 (
            .O(N__41927),
            .I(N__41919));
    Span4Mux_h I__9069 (
            .O(N__41922),
            .I(N__41916));
    LocalMux I__9068 (
            .O(N__41919),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    Odrv4 I__9067 (
            .O(N__41916),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    InMux I__9066 (
            .O(N__41911),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ));
    CascadeMux I__9065 (
            .O(N__41908),
            .I(N__41904));
    CascadeMux I__9064 (
            .O(N__41907),
            .I(N__41901));
    InMux I__9063 (
            .O(N__41904),
            .I(N__41895));
    InMux I__9062 (
            .O(N__41901),
            .I(N__41895));
    InMux I__9061 (
            .O(N__41900),
            .I(N__41892));
    LocalMux I__9060 (
            .O(N__41895),
            .I(N__41889));
    LocalMux I__9059 (
            .O(N__41892),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    Odrv4 I__9058 (
            .O(N__41889),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    InMux I__9057 (
            .O(N__41884),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ));
    CascadeMux I__9056 (
            .O(N__41881),
            .I(N__41877));
    CascadeMux I__9055 (
            .O(N__41880),
            .I(N__41874));
    InMux I__9054 (
            .O(N__41877),
            .I(N__41868));
    InMux I__9053 (
            .O(N__41874),
            .I(N__41868));
    InMux I__9052 (
            .O(N__41873),
            .I(N__41865));
    LocalMux I__9051 (
            .O(N__41868),
            .I(N__41862));
    LocalMux I__9050 (
            .O(N__41865),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    Odrv4 I__9049 (
            .O(N__41862),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    InMux I__9048 (
            .O(N__41857),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ));
    InMux I__9047 (
            .O(N__41854),
            .I(N__41851));
    LocalMux I__9046 (
            .O(N__41851),
            .I(N__41848));
    Span4Mux_v I__9045 (
            .O(N__41848),
            .I(N__41845));
    Odrv4 I__9044 (
            .O(N__41845),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_21 ));
    InMux I__9043 (
            .O(N__41842),
            .I(N__41838));
    InMux I__9042 (
            .O(N__41841),
            .I(N__41835));
    LocalMux I__9041 (
            .O(N__41838),
            .I(N__41832));
    LocalMux I__9040 (
            .O(N__41835),
            .I(N__41829));
    Span4Mux_h I__9039 (
            .O(N__41832),
            .I(N__41825));
    Span4Mux_h I__9038 (
            .O(N__41829),
            .I(N__41822));
    InMux I__9037 (
            .O(N__41828),
            .I(N__41819));
    Odrv4 I__9036 (
            .O(N__41825),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_21 ));
    Odrv4 I__9035 (
            .O(N__41822),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_21 ));
    LocalMux I__9034 (
            .O(N__41819),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_21 ));
    InMux I__9033 (
            .O(N__41812),
            .I(N__41809));
    LocalMux I__9032 (
            .O(N__41809),
            .I(\current_shift_inst.PI_CTRL.error_control_RNI9BAQZ0Z_21 ));
    InMux I__9031 (
            .O(N__41806),
            .I(N__41803));
    LocalMux I__9030 (
            .O(N__41803),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ));
    CascadeMux I__9029 (
            .O(N__41800),
            .I(N__41796));
    InMux I__9028 (
            .O(N__41799),
            .I(N__41793));
    InMux I__9027 (
            .O(N__41796),
            .I(N__41790));
    LocalMux I__9026 (
            .O(N__41793),
            .I(N__41786));
    LocalMux I__9025 (
            .O(N__41790),
            .I(N__41783));
    InMux I__9024 (
            .O(N__41789),
            .I(N__41780));
    Span4Mux_v I__9023 (
            .O(N__41786),
            .I(N__41775));
    Span4Mux_h I__9022 (
            .O(N__41783),
            .I(N__41770));
    LocalMux I__9021 (
            .O(N__41780),
            .I(N__41770));
    InMux I__9020 (
            .O(N__41779),
            .I(N__41767));
    CascadeMux I__9019 (
            .O(N__41778),
            .I(N__41764));
    Span4Mux_h I__9018 (
            .O(N__41775),
            .I(N__41757));
    Span4Mux_v I__9017 (
            .O(N__41770),
            .I(N__41757));
    LocalMux I__9016 (
            .O(N__41767),
            .I(N__41757));
    InMux I__9015 (
            .O(N__41764),
            .I(N__41754));
    Span4Mux_h I__9014 (
            .O(N__41757),
            .I(N__41751));
    LocalMux I__9013 (
            .O(N__41754),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    Odrv4 I__9012 (
            .O(N__41751),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    InMux I__9011 (
            .O(N__41746),
            .I(N__41743));
    LocalMux I__9010 (
            .O(N__41743),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ));
    CascadeMux I__9009 (
            .O(N__41740),
            .I(N__41736));
    InMux I__9008 (
            .O(N__41739),
            .I(N__41733));
    InMux I__9007 (
            .O(N__41736),
            .I(N__41730));
    LocalMux I__9006 (
            .O(N__41733),
            .I(N__41725));
    LocalMux I__9005 (
            .O(N__41730),
            .I(N__41722));
    InMux I__9004 (
            .O(N__41729),
            .I(N__41719));
    InMux I__9003 (
            .O(N__41728),
            .I(N__41715));
    Span4Mux_v I__9002 (
            .O(N__41725),
            .I(N__41712));
    Span4Mux_v I__9001 (
            .O(N__41722),
            .I(N__41709));
    LocalMux I__9000 (
            .O(N__41719),
            .I(N__41706));
    InMux I__8999 (
            .O(N__41718),
            .I(N__41703));
    LocalMux I__8998 (
            .O(N__41715),
            .I(N__41700));
    Span4Mux_h I__8997 (
            .O(N__41712),
            .I(N__41691));
    Span4Mux_h I__8996 (
            .O(N__41709),
            .I(N__41691));
    Span4Mux_v I__8995 (
            .O(N__41706),
            .I(N__41691));
    LocalMux I__8994 (
            .O(N__41703),
            .I(N__41691));
    Span4Mux_h I__8993 (
            .O(N__41700),
            .I(N__41688));
    Span4Mux_h I__8992 (
            .O(N__41691),
            .I(N__41685));
    Odrv4 I__8991 (
            .O(N__41688),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv4 I__8990 (
            .O(N__41685),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    InMux I__8989 (
            .O(N__41680),
            .I(N__41677));
    LocalMux I__8988 (
            .O(N__41677),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ));
    CascadeMux I__8987 (
            .O(N__41674),
            .I(N__41671));
    InMux I__8986 (
            .O(N__41671),
            .I(N__41667));
    InMux I__8985 (
            .O(N__41670),
            .I(N__41664));
    LocalMux I__8984 (
            .O(N__41667),
            .I(N__41659));
    LocalMux I__8983 (
            .O(N__41664),
            .I(N__41656));
    InMux I__8982 (
            .O(N__41663),
            .I(N__41651));
    InMux I__8981 (
            .O(N__41662),
            .I(N__41651));
    Span4Mux_h I__8980 (
            .O(N__41659),
            .I(N__41644));
    Span4Mux_h I__8979 (
            .O(N__41656),
            .I(N__41644));
    LocalMux I__8978 (
            .O(N__41651),
            .I(N__41644));
    Span4Mux_h I__8977 (
            .O(N__41644),
            .I(N__41641));
    Span4Mux_h I__8976 (
            .O(N__41641),
            .I(N__41637));
    InMux I__8975 (
            .O(N__41640),
            .I(N__41634));
    Odrv4 I__8974 (
            .O(N__41637),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    LocalMux I__8973 (
            .O(N__41634),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    CascadeMux I__8972 (
            .O(N__41629),
            .I(N__41626));
    InMux I__8971 (
            .O(N__41626),
            .I(N__41623));
    LocalMux I__8970 (
            .O(N__41623),
            .I(N__41620));
    Odrv4 I__8969 (
            .O(N__41620),
            .I(\current_shift_inst.PI_CTRL.integrator_i_12 ));
    InMux I__8968 (
            .O(N__41617),
            .I(bfn_17_11_0_));
    InMux I__8967 (
            .O(N__41614),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ));
    CascadeMux I__8966 (
            .O(N__41611),
            .I(N__41607));
    CascadeMux I__8965 (
            .O(N__41610),
            .I(N__41604));
    InMux I__8964 (
            .O(N__41607),
            .I(N__41598));
    InMux I__8963 (
            .O(N__41604),
            .I(N__41598));
    InMux I__8962 (
            .O(N__41603),
            .I(N__41595));
    LocalMux I__8961 (
            .O(N__41598),
            .I(N__41592));
    LocalMux I__8960 (
            .O(N__41595),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    Odrv4 I__8959 (
            .O(N__41592),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    InMux I__8958 (
            .O(N__41587),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ));
    InMux I__8957 (
            .O(N__41584),
            .I(N__41581));
    LocalMux I__8956 (
            .O(N__41581),
            .I(N__41578));
    Span4Mux_h I__8955 (
            .O(N__41578),
            .I(N__41575));
    Odrv4 I__8954 (
            .O(N__41575),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ));
    InMux I__8953 (
            .O(N__41572),
            .I(N__41568));
    InMux I__8952 (
            .O(N__41571),
            .I(N__41565));
    LocalMux I__8951 (
            .O(N__41568),
            .I(N__41562));
    LocalMux I__8950 (
            .O(N__41565),
            .I(N__41559));
    Span4Mux_h I__8949 (
            .O(N__41562),
            .I(N__41555));
    Span4Mux_h I__8948 (
            .O(N__41559),
            .I(N__41552));
    InMux I__8947 (
            .O(N__41558),
            .I(N__41549));
    Odrv4 I__8946 (
            .O(N__41555),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_18 ));
    Odrv4 I__8945 (
            .O(N__41552),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_18 ));
    LocalMux I__8944 (
            .O(N__41549),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_18 ));
    InMux I__8943 (
            .O(N__41542),
            .I(N__41539));
    LocalMux I__8942 (
            .O(N__41539),
            .I(N__41536));
    Span4Mux_h I__8941 (
            .O(N__41536),
            .I(N__41533));
    Odrv4 I__8940 (
            .O(N__41533),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_18 ));
    InMux I__8939 (
            .O(N__41530),
            .I(N__41527));
    LocalMux I__8938 (
            .O(N__41527),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIOTCPZ0Z_18 ));
    CascadeMux I__8937 (
            .O(N__41524),
            .I(N__41520));
    InMux I__8936 (
            .O(N__41523),
            .I(N__41516));
    InMux I__8935 (
            .O(N__41520),
            .I(N__41509));
    InMux I__8934 (
            .O(N__41519),
            .I(N__41509));
    LocalMux I__8933 (
            .O(N__41516),
            .I(N__41506));
    InMux I__8932 (
            .O(N__41515),
            .I(N__41501));
    InMux I__8931 (
            .O(N__41514),
            .I(N__41501));
    LocalMux I__8930 (
            .O(N__41509),
            .I(N__41498));
    Span4Mux_v I__8929 (
            .O(N__41506),
            .I(N__41495));
    LocalMux I__8928 (
            .O(N__41501),
            .I(N__41492));
    Span4Mux_h I__8927 (
            .O(N__41498),
            .I(N__41489));
    Odrv4 I__8926 (
            .O(N__41495),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    Odrv4 I__8925 (
            .O(N__41492),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    Odrv4 I__8924 (
            .O(N__41489),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    CascadeMux I__8923 (
            .O(N__41482),
            .I(N__41479));
    InMux I__8922 (
            .O(N__41479),
            .I(N__41476));
    LocalMux I__8921 (
            .O(N__41476),
            .I(\current_shift_inst.PI_CTRL.integrator_i_14 ));
    CascadeMux I__8920 (
            .O(N__41473),
            .I(N__41470));
    InMux I__8919 (
            .O(N__41470),
            .I(N__41467));
    LocalMux I__8918 (
            .O(N__41467),
            .I(\current_shift_inst.PI_CTRL.integrator_i_8 ));
    InMux I__8917 (
            .O(N__41464),
            .I(N__41461));
    LocalMux I__8916 (
            .O(N__41461),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ));
    InMux I__8915 (
            .O(N__41458),
            .I(N__41455));
    LocalMux I__8914 (
            .O(N__41455),
            .I(N__41450));
    InMux I__8913 (
            .O(N__41454),
            .I(N__41447));
    CascadeMux I__8912 (
            .O(N__41453),
            .I(N__41443));
    Span4Mux_v I__8911 (
            .O(N__41450),
            .I(N__41438));
    LocalMux I__8910 (
            .O(N__41447),
            .I(N__41438));
    InMux I__8909 (
            .O(N__41446),
            .I(N__41435));
    InMux I__8908 (
            .O(N__41443),
            .I(N__41432));
    Span4Mux_h I__8907 (
            .O(N__41438),
            .I(N__41429));
    LocalMux I__8906 (
            .O(N__41435),
            .I(N__41425));
    LocalMux I__8905 (
            .O(N__41432),
            .I(N__41420));
    Span4Mux_h I__8904 (
            .O(N__41429),
            .I(N__41420));
    InMux I__8903 (
            .O(N__41428),
            .I(N__41417));
    Odrv12 I__8902 (
            .O(N__41425),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    Odrv4 I__8901 (
            .O(N__41420),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    LocalMux I__8900 (
            .O(N__41417),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    InMux I__8899 (
            .O(N__41410),
            .I(N__41407));
    LocalMux I__8898 (
            .O(N__41407),
            .I(N__41404));
    Span4Mux_v I__8897 (
            .O(N__41404),
            .I(N__41401));
    Odrv4 I__8896 (
            .O(N__41401),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_25 ));
    InMux I__8895 (
            .O(N__41398),
            .I(N__41395));
    LocalMux I__8894 (
            .O(N__41395),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIGNFQZ0Z_25 ));
    InMux I__8893 (
            .O(N__41392),
            .I(N__41387));
    InMux I__8892 (
            .O(N__41391),
            .I(N__41382));
    InMux I__8891 (
            .O(N__41390),
            .I(N__41382));
    LocalMux I__8890 (
            .O(N__41387),
            .I(N__41379));
    LocalMux I__8889 (
            .O(N__41382),
            .I(N__41376));
    Span4Mux_h I__8888 (
            .O(N__41379),
            .I(N__41373));
    Span4Mux_h I__8887 (
            .O(N__41376),
            .I(N__41370));
    Odrv4 I__8886 (
            .O(N__41373),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_25 ));
    Odrv4 I__8885 (
            .O(N__41370),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_25 ));
    InMux I__8884 (
            .O(N__41365),
            .I(N__41362));
    LocalMux I__8883 (
            .O(N__41362),
            .I(N__41359));
    Span4Mux_h I__8882 (
            .O(N__41359),
            .I(N__41356));
    Odrv4 I__8881 (
            .O(N__41356),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ));
    InMux I__8880 (
            .O(N__41353),
            .I(N__41350));
    LocalMux I__8879 (
            .O(N__41350),
            .I(N__41347));
    Odrv4 I__8878 (
            .O(N__41347),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ));
    InMux I__8877 (
            .O(N__41344),
            .I(N__41341));
    LocalMux I__8876 (
            .O(N__41341),
            .I(N__41335));
    InMux I__8875 (
            .O(N__41340),
            .I(N__41332));
    InMux I__8874 (
            .O(N__41339),
            .I(N__41329));
    InMux I__8873 (
            .O(N__41338),
            .I(N__41326));
    Span4Mux_v I__8872 (
            .O(N__41335),
            .I(N__41323));
    LocalMux I__8871 (
            .O(N__41332),
            .I(N__41320));
    LocalMux I__8870 (
            .O(N__41329),
            .I(N__41316));
    LocalMux I__8869 (
            .O(N__41326),
            .I(N__41313));
    Span4Mux_h I__8868 (
            .O(N__41323),
            .I(N__41308));
    Span4Mux_v I__8867 (
            .O(N__41320),
            .I(N__41308));
    InMux I__8866 (
            .O(N__41319),
            .I(N__41305));
    Span4Mux_v I__8865 (
            .O(N__41316),
            .I(N__41302));
    Span4Mux_v I__8864 (
            .O(N__41313),
            .I(N__41299));
    Span4Mux_h I__8863 (
            .O(N__41308),
            .I(N__41294));
    LocalMux I__8862 (
            .O(N__41305),
            .I(N__41294));
    Span4Mux_h I__8861 (
            .O(N__41302),
            .I(N__41291));
    Odrv4 I__8860 (
            .O(N__41299),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    Odrv4 I__8859 (
            .O(N__41294),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    Odrv4 I__8858 (
            .O(N__41291),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    InMux I__8857 (
            .O(N__41284),
            .I(N__41281));
    LocalMux I__8856 (
            .O(N__41281),
            .I(N__41278));
    Odrv4 I__8855 (
            .O(N__41278),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ));
    InMux I__8854 (
            .O(N__41275),
            .I(N__41272));
    LocalMux I__8853 (
            .O(N__41272),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ));
    InMux I__8852 (
            .O(N__41269),
            .I(N__41266));
    LocalMux I__8851 (
            .O(N__41266),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ));
    InMux I__8850 (
            .O(N__41263),
            .I(N__41260));
    LocalMux I__8849 (
            .O(N__41260),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISST11_17 ));
    InMux I__8848 (
            .O(N__41257),
            .I(N__41253));
    InMux I__8847 (
            .O(N__41256),
            .I(N__41250));
    LocalMux I__8846 (
            .O(N__41253),
            .I(measured_delay_hc_29));
    LocalMux I__8845 (
            .O(N__41250),
            .I(measured_delay_hc_29));
    InMux I__8844 (
            .O(N__41245),
            .I(N__41241));
    InMux I__8843 (
            .O(N__41244),
            .I(N__41238));
    LocalMux I__8842 (
            .O(N__41241),
            .I(measured_delay_hc_30));
    LocalMux I__8841 (
            .O(N__41238),
            .I(measured_delay_hc_30));
    InMux I__8840 (
            .O(N__41233),
            .I(N__41229));
    InMux I__8839 (
            .O(N__41232),
            .I(N__41226));
    LocalMux I__8838 (
            .O(N__41229),
            .I(measured_delay_hc_27));
    LocalMux I__8837 (
            .O(N__41226),
            .I(measured_delay_hc_27));
    CascadeMux I__8836 (
            .O(N__41221),
            .I(N__41216));
    CascadeMux I__8835 (
            .O(N__41220),
            .I(N__41204));
    CascadeMux I__8834 (
            .O(N__41219),
            .I(N__41200));
    InMux I__8833 (
            .O(N__41216),
            .I(N__41188));
    InMux I__8832 (
            .O(N__41215),
            .I(N__41188));
    InMux I__8831 (
            .O(N__41214),
            .I(N__41188));
    InMux I__8830 (
            .O(N__41213),
            .I(N__41180));
    InMux I__8829 (
            .O(N__41212),
            .I(N__41177));
    CascadeMux I__8828 (
            .O(N__41211),
            .I(N__41174));
    CascadeMux I__8827 (
            .O(N__41210),
            .I(N__41171));
    CascadeMux I__8826 (
            .O(N__41209),
            .I(N__41166));
    CascadeMux I__8825 (
            .O(N__41208),
            .I(N__41163));
    CascadeMux I__8824 (
            .O(N__41207),
            .I(N__41160));
    InMux I__8823 (
            .O(N__41204),
            .I(N__41150));
    InMux I__8822 (
            .O(N__41203),
            .I(N__41143));
    InMux I__8821 (
            .O(N__41200),
            .I(N__41143));
    InMux I__8820 (
            .O(N__41199),
            .I(N__41143));
    InMux I__8819 (
            .O(N__41198),
            .I(N__41134));
    InMux I__8818 (
            .O(N__41197),
            .I(N__41134));
    InMux I__8817 (
            .O(N__41196),
            .I(N__41134));
    InMux I__8816 (
            .O(N__41195),
            .I(N__41134));
    LocalMux I__8815 (
            .O(N__41188),
            .I(N__41131));
    InMux I__8814 (
            .O(N__41187),
            .I(N__41128));
    InMux I__8813 (
            .O(N__41186),
            .I(N__41119));
    InMux I__8812 (
            .O(N__41185),
            .I(N__41119));
    InMux I__8811 (
            .O(N__41184),
            .I(N__41119));
    InMux I__8810 (
            .O(N__41183),
            .I(N__41119));
    LocalMux I__8809 (
            .O(N__41180),
            .I(N__41114));
    LocalMux I__8808 (
            .O(N__41177),
            .I(N__41114));
    InMux I__8807 (
            .O(N__41174),
            .I(N__41105));
    InMux I__8806 (
            .O(N__41171),
            .I(N__41105));
    InMux I__8805 (
            .O(N__41170),
            .I(N__41105));
    InMux I__8804 (
            .O(N__41169),
            .I(N__41105));
    InMux I__8803 (
            .O(N__41166),
            .I(N__41094));
    InMux I__8802 (
            .O(N__41163),
            .I(N__41094));
    InMux I__8801 (
            .O(N__41160),
            .I(N__41094));
    InMux I__8800 (
            .O(N__41159),
            .I(N__41094));
    InMux I__8799 (
            .O(N__41158),
            .I(N__41094));
    InMux I__8798 (
            .O(N__41157),
            .I(N__41083));
    InMux I__8797 (
            .O(N__41156),
            .I(N__41083));
    InMux I__8796 (
            .O(N__41155),
            .I(N__41083));
    InMux I__8795 (
            .O(N__41154),
            .I(N__41083));
    InMux I__8794 (
            .O(N__41153),
            .I(N__41083));
    LocalMux I__8793 (
            .O(N__41150),
            .I(N__41074));
    LocalMux I__8792 (
            .O(N__41143),
            .I(N__41074));
    LocalMux I__8791 (
            .O(N__41134),
            .I(N__41074));
    Span4Mux_h I__8790 (
            .O(N__41131),
            .I(N__41074));
    LocalMux I__8789 (
            .O(N__41128),
            .I(N__41071));
    LocalMux I__8788 (
            .O(N__41119),
            .I(N__41068));
    Span4Mux_h I__8787 (
            .O(N__41114),
            .I(N__41065));
    LocalMux I__8786 (
            .O(N__41105),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    LocalMux I__8785 (
            .O(N__41094),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    LocalMux I__8784 (
            .O(N__41083),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    Odrv4 I__8783 (
            .O(N__41074),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    Odrv12 I__8782 (
            .O(N__41071),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    Odrv12 I__8781 (
            .O(N__41068),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    Odrv4 I__8780 (
            .O(N__41065),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    InMux I__8779 (
            .O(N__41050),
            .I(N__41043));
    InMux I__8778 (
            .O(N__41049),
            .I(N__41025));
    InMux I__8777 (
            .O(N__41048),
            .I(N__41025));
    InMux I__8776 (
            .O(N__41047),
            .I(N__41025));
    InMux I__8775 (
            .O(N__41046),
            .I(N__41022));
    LocalMux I__8774 (
            .O(N__41043),
            .I(N__41009));
    InMux I__8773 (
            .O(N__41042),
            .I(N__41002));
    InMux I__8772 (
            .O(N__41041),
            .I(N__41002));
    InMux I__8771 (
            .O(N__41040),
            .I(N__41002));
    InMux I__8770 (
            .O(N__41039),
            .I(N__40993));
    InMux I__8769 (
            .O(N__41038),
            .I(N__40993));
    InMux I__8768 (
            .O(N__41037),
            .I(N__40993));
    InMux I__8767 (
            .O(N__41036),
            .I(N__40993));
    InMux I__8766 (
            .O(N__41035),
            .I(N__40984));
    InMux I__8765 (
            .O(N__41034),
            .I(N__40984));
    InMux I__8764 (
            .O(N__41033),
            .I(N__40984));
    InMux I__8763 (
            .O(N__41032),
            .I(N__40984));
    LocalMux I__8762 (
            .O(N__41025),
            .I(N__40975));
    LocalMux I__8761 (
            .O(N__41022),
            .I(N__40972));
    InMux I__8760 (
            .O(N__41021),
            .I(N__40959));
    InMux I__8759 (
            .O(N__41020),
            .I(N__40959));
    InMux I__8758 (
            .O(N__41019),
            .I(N__40959));
    InMux I__8757 (
            .O(N__41018),
            .I(N__40959));
    InMux I__8756 (
            .O(N__41017),
            .I(N__40959));
    InMux I__8755 (
            .O(N__41016),
            .I(N__40959));
    InMux I__8754 (
            .O(N__41015),
            .I(N__40950));
    InMux I__8753 (
            .O(N__41014),
            .I(N__40950));
    InMux I__8752 (
            .O(N__41013),
            .I(N__40950));
    InMux I__8751 (
            .O(N__41012),
            .I(N__40950));
    Span4Mux_h I__8750 (
            .O(N__41009),
            .I(N__40947));
    LocalMux I__8749 (
            .O(N__41002),
            .I(N__40944));
    LocalMux I__8748 (
            .O(N__40993),
            .I(N__40939));
    LocalMux I__8747 (
            .O(N__40984),
            .I(N__40939));
    InMux I__8746 (
            .O(N__40983),
            .I(N__40936));
    InMux I__8745 (
            .O(N__40982),
            .I(N__40925));
    InMux I__8744 (
            .O(N__40981),
            .I(N__40925));
    InMux I__8743 (
            .O(N__40980),
            .I(N__40925));
    InMux I__8742 (
            .O(N__40979),
            .I(N__40925));
    InMux I__8741 (
            .O(N__40978),
            .I(N__40925));
    Span4Mux_h I__8740 (
            .O(N__40975),
            .I(N__40916));
    Span4Mux_h I__8739 (
            .O(N__40972),
            .I(N__40916));
    LocalMux I__8738 (
            .O(N__40959),
            .I(N__40916));
    LocalMux I__8737 (
            .O(N__40950),
            .I(N__40916));
    Odrv4 I__8736 (
            .O(N__40947),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    Odrv12 I__8735 (
            .O(N__40944),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    Odrv12 I__8734 (
            .O(N__40939),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    LocalMux I__8733 (
            .O(N__40936),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    LocalMux I__8732 (
            .O(N__40925),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    Odrv4 I__8731 (
            .O(N__40916),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    InMux I__8730 (
            .O(N__40903),
            .I(N__40899));
    InMux I__8729 (
            .O(N__40902),
            .I(N__40896));
    LocalMux I__8728 (
            .O(N__40899),
            .I(measured_delay_hc_28));
    LocalMux I__8727 (
            .O(N__40896),
            .I(measured_delay_hc_28));
    InMux I__8726 (
            .O(N__40891),
            .I(N__40888));
    LocalMux I__8725 (
            .O(N__40888),
            .I(N__40885));
    Odrv4 I__8724 (
            .O(N__40885),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ));
    InMux I__8723 (
            .O(N__40882),
            .I(N__40878));
    CascadeMux I__8722 (
            .O(N__40881),
            .I(N__40874));
    LocalMux I__8721 (
            .O(N__40878),
            .I(N__40870));
    InMux I__8720 (
            .O(N__40877),
            .I(N__40867));
    InMux I__8719 (
            .O(N__40874),
            .I(N__40864));
    InMux I__8718 (
            .O(N__40873),
            .I(N__40861));
    Span4Mux_v I__8717 (
            .O(N__40870),
            .I(N__40858));
    LocalMux I__8716 (
            .O(N__40867),
            .I(N__40855));
    LocalMux I__8715 (
            .O(N__40864),
            .I(N__40851));
    LocalMux I__8714 (
            .O(N__40861),
            .I(N__40844));
    Span4Mux_h I__8713 (
            .O(N__40858),
            .I(N__40844));
    Span4Mux_v I__8712 (
            .O(N__40855),
            .I(N__40844));
    InMux I__8711 (
            .O(N__40854),
            .I(N__40841));
    Span12Mux_v I__8710 (
            .O(N__40851),
            .I(N__40838));
    Span4Mux_h I__8709 (
            .O(N__40844),
            .I(N__40833));
    LocalMux I__8708 (
            .O(N__40841),
            .I(N__40833));
    Odrv12 I__8707 (
            .O(N__40838),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    Odrv4 I__8706 (
            .O(N__40833),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    CascadeMux I__8705 (
            .O(N__40828),
            .I(N__40825));
    InMux I__8704 (
            .O(N__40825),
            .I(N__40822));
    LocalMux I__8703 (
            .O(N__40822),
            .I(N__40819));
    Span4Mux_v I__8702 (
            .O(N__40819),
            .I(N__40816));
    Odrv4 I__8701 (
            .O(N__40816),
            .I(\current_shift_inst.PI_CTRL.integrator_i_25 ));
    InMux I__8700 (
            .O(N__40813),
            .I(N__40810));
    LocalMux I__8699 (
            .O(N__40810),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI25021_19 ));
    InMux I__8698 (
            .O(N__40807),
            .I(N__40804));
    LocalMux I__8697 (
            .O(N__40804),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ));
    InMux I__8696 (
            .O(N__40801),
            .I(N__40798));
    LocalMux I__8695 (
            .O(N__40798),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ));
    InMux I__8694 (
            .O(N__40795),
            .I(N__40792));
    LocalMux I__8693 (
            .O(N__40792),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ));
    InMux I__8692 (
            .O(N__40789),
            .I(N__40786));
    LocalMux I__8691 (
            .O(N__40786),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ));
    InMux I__8690 (
            .O(N__40783),
            .I(N__40780));
    LocalMux I__8689 (
            .O(N__40780),
            .I(N__40777));
    Span4Mux_h I__8688 (
            .O(N__40777),
            .I(N__40773));
    InMux I__8687 (
            .O(N__40776),
            .I(N__40770));
    Odrv4 I__8686 (
            .O(N__40773),
            .I(\current_shift_inst.un4_control_input_0_31 ));
    LocalMux I__8685 (
            .O(N__40770),
            .I(\current_shift_inst.un4_control_input_0_31 ));
    InMux I__8684 (
            .O(N__40765),
            .I(N__40762));
    LocalMux I__8683 (
            .O(N__40762),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ));
    InMux I__8682 (
            .O(N__40759),
            .I(N__40756));
    LocalMux I__8681 (
            .O(N__40756),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ));
    InMux I__8680 (
            .O(N__40753),
            .I(N__40750));
    LocalMux I__8679 (
            .O(N__40750),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_16 ));
    CascadeMux I__8678 (
            .O(N__40747),
            .I(N__40744));
    InMux I__8677 (
            .O(N__40744),
            .I(N__40741));
    LocalMux I__8676 (
            .O(N__40741),
            .I(N__40738));
    Odrv4 I__8675 (
            .O(N__40738),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ));
    InMux I__8674 (
            .O(N__40735),
            .I(N__40732));
    LocalMux I__8673 (
            .O(N__40732),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11 ));
    InMux I__8672 (
            .O(N__40729),
            .I(N__40726));
    LocalMux I__8671 (
            .O(N__40726),
            .I(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ));
    InMux I__8670 (
            .O(N__40723),
            .I(N__40720));
    LocalMux I__8669 (
            .O(N__40720),
            .I(\current_shift_inst.elapsed_time_ns_1_RNID8O11_12 ));
    InMux I__8668 (
            .O(N__40717),
            .I(N__40714));
    LocalMux I__8667 (
            .O(N__40714),
            .I(\current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0 ));
    CascadeMux I__8666 (
            .O(N__40711),
            .I(N__40708));
    InMux I__8665 (
            .O(N__40708),
            .I(N__40705));
    LocalMux I__8664 (
            .O(N__40705),
            .I(N__40702));
    Odrv12 I__8663 (
            .O(N__40702),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ));
    InMux I__8662 (
            .O(N__40699),
            .I(N__40696));
    LocalMux I__8661 (
            .O(N__40696),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_18 ));
    InMux I__8660 (
            .O(N__40693),
            .I(N__40690));
    LocalMux I__8659 (
            .O(N__40690),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJO221_20 ));
    InMux I__8658 (
            .O(N__40687),
            .I(N__40684));
    LocalMux I__8657 (
            .O(N__40684),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_15 ));
    CascadeMux I__8656 (
            .O(N__40681),
            .I(N__40678));
    InMux I__8655 (
            .O(N__40678),
            .I(N__40675));
    LocalMux I__8654 (
            .O(N__40675),
            .I(N__40672));
    Span4Mux_h I__8653 (
            .O(N__40672),
            .I(N__40669));
    Odrv4 I__8652 (
            .O(N__40669),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ));
    InMux I__8651 (
            .O(N__40666),
            .I(N__40663));
    LocalMux I__8650 (
            .O(N__40663),
            .I(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ));
    InMux I__8649 (
            .O(N__40660),
            .I(N__40657));
    LocalMux I__8648 (
            .O(N__40657),
            .I(\current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0 ));
    InMux I__8647 (
            .O(N__40654),
            .I(N__40651));
    LocalMux I__8646 (
            .O(N__40651),
            .I(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ));
    CascadeMux I__8645 (
            .O(N__40648),
            .I(N__40645));
    InMux I__8644 (
            .O(N__40645),
            .I(N__40642));
    LocalMux I__8643 (
            .O(N__40642),
            .I(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ));
    InMux I__8642 (
            .O(N__40639),
            .I(N__40636));
    LocalMux I__8641 (
            .O(N__40636),
            .I(N__40633));
    Span4Mux_v I__8640 (
            .O(N__40633),
            .I(N__40630));
    Odrv4 I__8639 (
            .O(N__40630),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ));
    InMux I__8638 (
            .O(N__40627),
            .I(N__40624));
    LocalMux I__8637 (
            .O(N__40624),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_9 ));
    InMux I__8636 (
            .O(N__40621),
            .I(N__40618));
    LocalMux I__8635 (
            .O(N__40618),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14 ));
    InMux I__8634 (
            .O(N__40615),
            .I(N__40612));
    LocalMux I__8633 (
            .O(N__40612),
            .I(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ));
    InMux I__8632 (
            .O(N__40609),
            .I(N__40606));
    LocalMux I__8631 (
            .O(N__40606),
            .I(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ));
    InMux I__8630 (
            .O(N__40603),
            .I(N__40600));
    LocalMux I__8629 (
            .O(N__40600),
            .I(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ));
    InMux I__8628 (
            .O(N__40597),
            .I(N__40594));
    LocalMux I__8627 (
            .O(N__40594),
            .I(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ));
    InMux I__8626 (
            .O(N__40591),
            .I(N__40588));
    LocalMux I__8625 (
            .O(N__40588),
            .I(N__40585));
    Span4Mux_h I__8624 (
            .O(N__40585),
            .I(N__40582));
    Odrv4 I__8623 (
            .O(N__40582),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20 ));
    InMux I__8622 (
            .O(N__40579),
            .I(N__40576));
    LocalMux I__8621 (
            .O(N__40576),
            .I(N__40573));
    Span4Mux_v I__8620 (
            .O(N__40573),
            .I(N__40570));
    Odrv4 I__8619 (
            .O(N__40570),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10 ));
    InMux I__8618 (
            .O(N__40567),
            .I(N__40564));
    LocalMux I__8617 (
            .O(N__40564),
            .I(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ));
    InMux I__8616 (
            .O(N__40561),
            .I(N__40558));
    LocalMux I__8615 (
            .O(N__40558),
            .I(N__40555));
    Odrv4 I__8614 (
            .O(N__40555),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_13 ));
    InMux I__8613 (
            .O(N__40552),
            .I(N__40549));
    LocalMux I__8612 (
            .O(N__40549),
            .I(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ));
    InMux I__8611 (
            .O(N__40546),
            .I(N__40543));
    LocalMux I__8610 (
            .O(N__40543),
            .I(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ));
    InMux I__8609 (
            .O(N__40540),
            .I(N__40537));
    LocalMux I__8608 (
            .O(N__40537),
            .I(N__40534));
    Odrv4 I__8607 (
            .O(N__40534),
            .I(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ));
    InMux I__8606 (
            .O(N__40531),
            .I(N__40528));
    LocalMux I__8605 (
            .O(N__40528),
            .I(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ));
    InMux I__8604 (
            .O(N__40525),
            .I(N__40522));
    LocalMux I__8603 (
            .O(N__40522),
            .I(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ));
    InMux I__8602 (
            .O(N__40519),
            .I(N__40516));
    LocalMux I__8601 (
            .O(N__40516),
            .I(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ));
    InMux I__8600 (
            .O(N__40513),
            .I(N__40510));
    LocalMux I__8599 (
            .O(N__40510),
            .I(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ));
    InMux I__8598 (
            .O(N__40507),
            .I(N__40504));
    LocalMux I__8597 (
            .O(N__40504),
            .I(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ));
    InMux I__8596 (
            .O(N__40501),
            .I(N__40498));
    LocalMux I__8595 (
            .O(N__40498),
            .I(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ));
    InMux I__8594 (
            .O(N__40495),
            .I(N__40492));
    LocalMux I__8593 (
            .O(N__40492),
            .I(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ));
    InMux I__8592 (
            .O(N__40489),
            .I(N__40486));
    LocalMux I__8591 (
            .O(N__40486),
            .I(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ));
    InMux I__8590 (
            .O(N__40483),
            .I(N__40480));
    LocalMux I__8589 (
            .O(N__40480),
            .I(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ));
    InMux I__8588 (
            .O(N__40477),
            .I(N__40474));
    LocalMux I__8587 (
            .O(N__40474),
            .I(N__40471));
    Span4Mux_v I__8586 (
            .O(N__40471),
            .I(N__40468));
    Odrv4 I__8585 (
            .O(N__40468),
            .I(\current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0 ));
    InMux I__8584 (
            .O(N__40465),
            .I(N__40462));
    LocalMux I__8583 (
            .O(N__40462),
            .I(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ));
    InMux I__8582 (
            .O(N__40459),
            .I(N__40456));
    LocalMux I__8581 (
            .O(N__40456),
            .I(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ));
    InMux I__8580 (
            .O(N__40453),
            .I(N__40450));
    LocalMux I__8579 (
            .O(N__40450),
            .I(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ));
    CascadeMux I__8578 (
            .O(N__40447),
            .I(N__40444));
    InMux I__8577 (
            .O(N__40444),
            .I(N__40441));
    LocalMux I__8576 (
            .O(N__40441),
            .I(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ));
    InMux I__8575 (
            .O(N__40438),
            .I(N__40435));
    LocalMux I__8574 (
            .O(N__40435),
            .I(N__40432));
    Span4Mux_h I__8573 (
            .O(N__40432),
            .I(N__40429));
    Odrv4 I__8572 (
            .O(N__40429),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ));
    CascadeMux I__8571 (
            .O(N__40426),
            .I(N__40421));
    CascadeMux I__8570 (
            .O(N__40425),
            .I(N__40418));
    InMux I__8569 (
            .O(N__40424),
            .I(N__40412));
    InMux I__8568 (
            .O(N__40421),
            .I(N__40412));
    InMux I__8567 (
            .O(N__40418),
            .I(N__40409));
    CascadeMux I__8566 (
            .O(N__40417),
            .I(N__40406));
    LocalMux I__8565 (
            .O(N__40412),
            .I(N__40403));
    LocalMux I__8564 (
            .O(N__40409),
            .I(N__40400));
    InMux I__8563 (
            .O(N__40406),
            .I(N__40397));
    Span4Mux_h I__8562 (
            .O(N__40403),
            .I(N__40392));
    Span4Mux_h I__8561 (
            .O(N__40400),
            .I(N__40392));
    LocalMux I__8560 (
            .O(N__40397),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    Odrv4 I__8559 (
            .O(N__40392),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    InMux I__8558 (
            .O(N__40387),
            .I(N__40384));
    LocalMux I__8557 (
            .O(N__40384),
            .I(N__40381));
    Span4Mux_v I__8556 (
            .O(N__40381),
            .I(N__40378));
    Odrv4 I__8555 (
            .O(N__40378),
            .I(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ));
    InMux I__8554 (
            .O(N__40375),
            .I(N__40365));
    InMux I__8553 (
            .O(N__40374),
            .I(N__40365));
    InMux I__8552 (
            .O(N__40373),
            .I(N__40365));
    InMux I__8551 (
            .O(N__40372),
            .I(N__40362));
    LocalMux I__8550 (
            .O(N__40365),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    LocalMux I__8549 (
            .O(N__40362),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    InMux I__8548 (
            .O(N__40357),
            .I(N__40354));
    LocalMux I__8547 (
            .O(N__40354),
            .I(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ));
    CascadeMux I__8546 (
            .O(N__40351),
            .I(N__40348));
    InMux I__8545 (
            .O(N__40348),
            .I(N__40345));
    LocalMux I__8544 (
            .O(N__40345),
            .I(N__40342));
    Odrv4 I__8543 (
            .O(N__40342),
            .I(\current_shift_inst.PI_CTRL.integrator_i_18 ));
    InMux I__8542 (
            .O(N__40339),
            .I(N__40336));
    LocalMux I__8541 (
            .O(N__40336),
            .I(N__40333));
    Odrv12 I__8540 (
            .O(N__40333),
            .I(\current_shift_inst.PI_CTRL.integrator_i_19 ));
    InMux I__8539 (
            .O(N__40330),
            .I(N__40327));
    LocalMux I__8538 (
            .O(N__40327),
            .I(N__40322));
    InMux I__8537 (
            .O(N__40326),
            .I(N__40319));
    InMux I__8536 (
            .O(N__40325),
            .I(N__40316));
    Span4Mux_h I__8535 (
            .O(N__40322),
            .I(N__40313));
    LocalMux I__8534 (
            .O(N__40319),
            .I(N__40310));
    LocalMux I__8533 (
            .O(N__40316),
            .I(N__40307));
    Odrv4 I__8532 (
            .O(N__40313),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_24 ));
    Odrv4 I__8531 (
            .O(N__40310),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_24 ));
    Odrv4 I__8530 (
            .O(N__40307),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_24 ));
    InMux I__8529 (
            .O(N__40300),
            .I(N__40297));
    LocalMux I__8528 (
            .O(N__40297),
            .I(N__40294));
    Span4Mux_v I__8527 (
            .O(N__40294),
            .I(N__40291));
    Odrv4 I__8526 (
            .O(N__40291),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_24 ));
    InMux I__8525 (
            .O(N__40288),
            .I(N__40285));
    LocalMux I__8524 (
            .O(N__40285),
            .I(N__40282));
    Odrv4 I__8523 (
            .O(N__40282),
            .I(\current_shift_inst.PI_CTRL.error_control_RNICIEQZ0Z_24 ));
    InMux I__8522 (
            .O(N__40279),
            .I(N__40276));
    LocalMux I__8521 (
            .O(N__40276),
            .I(N__40273));
    Odrv4 I__8520 (
            .O(N__40273),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ));
    CascadeMux I__8519 (
            .O(N__40270),
            .I(N__40266));
    InMux I__8518 (
            .O(N__40269),
            .I(N__40263));
    InMux I__8517 (
            .O(N__40266),
            .I(N__40260));
    LocalMux I__8516 (
            .O(N__40263),
            .I(N__40255));
    LocalMux I__8515 (
            .O(N__40260),
            .I(N__40252));
    InMux I__8514 (
            .O(N__40259),
            .I(N__40249));
    CascadeMux I__8513 (
            .O(N__40258),
            .I(N__40246));
    Span4Mux_h I__8512 (
            .O(N__40255),
            .I(N__40241));
    Span4Mux_v I__8511 (
            .O(N__40252),
            .I(N__40241));
    LocalMux I__8510 (
            .O(N__40249),
            .I(N__40237));
    InMux I__8509 (
            .O(N__40246),
            .I(N__40234));
    Span4Mux_h I__8508 (
            .O(N__40241),
            .I(N__40231));
    InMux I__8507 (
            .O(N__40240),
            .I(N__40228));
    Span4Mux_h I__8506 (
            .O(N__40237),
            .I(N__40225));
    LocalMux I__8505 (
            .O(N__40234),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    Odrv4 I__8504 (
            .O(N__40231),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    LocalMux I__8503 (
            .O(N__40228),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    Odrv4 I__8502 (
            .O(N__40225),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    InMux I__8501 (
            .O(N__40216),
            .I(N__40213));
    LocalMux I__8500 (
            .O(N__40213),
            .I(N__40210));
    Odrv4 I__8499 (
            .O(N__40210),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ));
    CascadeMux I__8498 (
            .O(N__40207),
            .I(N__40202));
    InMux I__8497 (
            .O(N__40206),
            .I(N__40199));
    InMux I__8496 (
            .O(N__40205),
            .I(N__40196));
    InMux I__8495 (
            .O(N__40202),
            .I(N__40192));
    LocalMux I__8494 (
            .O(N__40199),
            .I(N__40189));
    LocalMux I__8493 (
            .O(N__40196),
            .I(N__40186));
    InMux I__8492 (
            .O(N__40195),
            .I(N__40183));
    LocalMux I__8491 (
            .O(N__40192),
            .I(N__40179));
    Span4Mux_h I__8490 (
            .O(N__40189),
            .I(N__40172));
    Span4Mux_v I__8489 (
            .O(N__40186),
            .I(N__40172));
    LocalMux I__8488 (
            .O(N__40183),
            .I(N__40172));
    InMux I__8487 (
            .O(N__40182),
            .I(N__40169));
    Span4Mux_v I__8486 (
            .O(N__40179),
            .I(N__40164));
    Span4Mux_h I__8485 (
            .O(N__40172),
            .I(N__40164));
    LocalMux I__8484 (
            .O(N__40169),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    Odrv4 I__8483 (
            .O(N__40164),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    InMux I__8482 (
            .O(N__40159),
            .I(N__40156));
    LocalMux I__8481 (
            .O(N__40156),
            .I(N__40153));
    Odrv4 I__8480 (
            .O(N__40153),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ));
    CascadeMux I__8479 (
            .O(N__40150),
            .I(N__40146));
    InMux I__8478 (
            .O(N__40149),
            .I(N__40143));
    InMux I__8477 (
            .O(N__40146),
            .I(N__40138));
    LocalMux I__8476 (
            .O(N__40143),
            .I(N__40135));
    InMux I__8475 (
            .O(N__40142),
            .I(N__40132));
    InMux I__8474 (
            .O(N__40141),
            .I(N__40129));
    LocalMux I__8473 (
            .O(N__40138),
            .I(N__40126));
    Span4Mux_v I__8472 (
            .O(N__40135),
            .I(N__40123));
    LocalMux I__8471 (
            .O(N__40132),
            .I(N__40118));
    LocalMux I__8470 (
            .O(N__40129),
            .I(N__40118));
    Span4Mux_v I__8469 (
            .O(N__40126),
            .I(N__40114));
    Span4Mux_h I__8468 (
            .O(N__40123),
            .I(N__40109));
    Span4Mux_v I__8467 (
            .O(N__40118),
            .I(N__40109));
    InMux I__8466 (
            .O(N__40117),
            .I(N__40106));
    Odrv4 I__8465 (
            .O(N__40114),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv4 I__8464 (
            .O(N__40109),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    LocalMux I__8463 (
            .O(N__40106),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    InMux I__8462 (
            .O(N__40099),
            .I(N__40096));
    LocalMux I__8461 (
            .O(N__40096),
            .I(N__40093));
    Span4Mux_h I__8460 (
            .O(N__40093),
            .I(N__40090));
    Odrv4 I__8459 (
            .O(N__40090),
            .I(\current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0 ));
    InMux I__8458 (
            .O(N__40087),
            .I(N__40084));
    LocalMux I__8457 (
            .O(N__40084),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNISPBJZ0 ));
    InMux I__8456 (
            .O(N__40081),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_25 ));
    InMux I__8455 (
            .O(N__40078),
            .I(N__40075));
    LocalMux I__8454 (
            .O(N__40075),
            .I(N__40072));
    Span4Mux_h I__8453 (
            .O(N__40072),
            .I(N__40069));
    Odrv4 I__8452 (
            .O(N__40069),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNILB5KZ0 ));
    CascadeMux I__8451 (
            .O(N__40066),
            .I(N__40063));
    InMux I__8450 (
            .O(N__40063),
            .I(N__40060));
    LocalMux I__8449 (
            .O(N__40060),
            .I(N__40057));
    Odrv4 I__8448 (
            .O(N__40057),
            .I(\current_shift_inst.PI_CTRL.integrator_i_27 ));
    InMux I__8447 (
            .O(N__40054),
            .I(N__40051));
    LocalMux I__8446 (
            .O(N__40051),
            .I(N__40048));
    Odrv12 I__8445 (
            .O(N__40048),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ));
    InMux I__8444 (
            .O(N__40045),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_26 ));
    InMux I__8443 (
            .O(N__40042),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_27 ));
    InMux I__8442 (
            .O(N__40039),
            .I(N__40036));
    LocalMux I__8441 (
            .O(N__40036),
            .I(N__40033));
    Odrv12 I__8440 (
            .O(N__40033),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ));
    InMux I__8439 (
            .O(N__40030),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_28 ));
    CascadeMux I__8438 (
            .O(N__40027),
            .I(N__40024));
    InMux I__8437 (
            .O(N__40024),
            .I(N__40021));
    LocalMux I__8436 (
            .O(N__40021),
            .I(N__40018));
    Span4Mux_h I__8435 (
            .O(N__40018),
            .I(N__40015));
    Odrv4 I__8434 (
            .O(N__40015),
            .I(\current_shift_inst.PI_CTRL.integrator_i_30 ));
    InMux I__8433 (
            .O(N__40012),
            .I(N__40009));
    LocalMux I__8432 (
            .O(N__40009),
            .I(N__40006));
    Odrv12 I__8431 (
            .O(N__40006),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ));
    InMux I__8430 (
            .O(N__40003),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_29 ));
    InMux I__8429 (
            .O(N__40000),
            .I(bfn_16_12_0_));
    InMux I__8428 (
            .O(N__39997),
            .I(N__39993));
    CascadeMux I__8427 (
            .O(N__39996),
            .I(N__39990));
    LocalMux I__8426 (
            .O(N__39993),
            .I(N__39986));
    InMux I__8425 (
            .O(N__39990),
            .I(N__39982));
    InMux I__8424 (
            .O(N__39989),
            .I(N__39979));
    Span4Mux_h I__8423 (
            .O(N__39986),
            .I(N__39976));
    InMux I__8422 (
            .O(N__39985),
            .I(N__39973));
    LocalMux I__8421 (
            .O(N__39982),
            .I(N__39970));
    LocalMux I__8420 (
            .O(N__39979),
            .I(N__39963));
    Span4Mux_h I__8419 (
            .O(N__39976),
            .I(N__39963));
    LocalMux I__8418 (
            .O(N__39973),
            .I(N__39963));
    Odrv4 I__8417 (
            .O(N__39970),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    Odrv4 I__8416 (
            .O(N__39963),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    InMux I__8415 (
            .O(N__39958),
            .I(N__39955));
    LocalMux I__8414 (
            .O(N__39955),
            .I(\current_shift_inst.PI_CTRL.integrator_i_29 ));
    CascadeMux I__8413 (
            .O(N__39952),
            .I(N__39949));
    InMux I__8412 (
            .O(N__39949),
            .I(N__39946));
    LocalMux I__8411 (
            .O(N__39946),
            .I(N__39943));
    Odrv4 I__8410 (
            .O(N__39943),
            .I(\current_shift_inst.PI_CTRL.integrator_i_20 ));
    CascadeMux I__8409 (
            .O(N__39940),
            .I(N__39936));
    InMux I__8408 (
            .O(N__39939),
            .I(N__39928));
    InMux I__8407 (
            .O(N__39936),
            .I(N__39928));
    InMux I__8406 (
            .O(N__39935),
            .I(N__39928));
    LocalMux I__8405 (
            .O(N__39928),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_i_0_26 ));
    InMux I__8404 (
            .O(N__39925),
            .I(N__39922));
    LocalMux I__8403 (
            .O(N__39922),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIDGBQZ0Z_22 ));
    InMux I__8402 (
            .O(N__39919),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_17 ));
    CascadeMux I__8401 (
            .O(N__39916),
            .I(N__39913));
    InMux I__8400 (
            .O(N__39913),
            .I(N__39910));
    LocalMux I__8399 (
            .O(N__39910),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIHLCQZ0Z_23 ));
    InMux I__8398 (
            .O(N__39907),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_18 ));
    InMux I__8397 (
            .O(N__39904),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_19 ));
    CascadeMux I__8396 (
            .O(N__39901),
            .I(N__39898));
    InMux I__8395 (
            .O(N__39898),
            .I(N__39895));
    LocalMux I__8394 (
            .O(N__39895),
            .I(N__39892));
    Span4Mux_v I__8393 (
            .O(N__39892),
            .I(N__39889));
    Odrv4 I__8392 (
            .O(N__39889),
            .I(\current_shift_inst.PI_CTRL.integrator_i_21 ));
    InMux I__8391 (
            .O(N__39886),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_20 ));
    InMux I__8390 (
            .O(N__39883),
            .I(N__39880));
    LocalMux I__8389 (
            .O(N__39880),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIKD7JZ0 ));
    CascadeMux I__8388 (
            .O(N__39877),
            .I(N__39874));
    InMux I__8387 (
            .O(N__39874),
            .I(N__39871));
    LocalMux I__8386 (
            .O(N__39871),
            .I(N__39868));
    Span4Mux_v I__8385 (
            .O(N__39868),
            .I(N__39865));
    Odrv4 I__8384 (
            .O(N__39865),
            .I(\current_shift_inst.PI_CTRL.integrator_i_22 ));
    InMux I__8383 (
            .O(N__39862),
            .I(N__39859));
    LocalMux I__8382 (
            .O(N__39859),
            .I(N__39856));
    Odrv12 I__8381 (
            .O(N__39856),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ));
    InMux I__8380 (
            .O(N__39853),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_21 ));
    InMux I__8379 (
            .O(N__39850),
            .I(N__39847));
    LocalMux I__8378 (
            .O(N__39847),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIMG8JZ0 ));
    InMux I__8377 (
            .O(N__39844),
            .I(bfn_16_11_0_));
    InMux I__8376 (
            .O(N__39841),
            .I(N__39838));
    LocalMux I__8375 (
            .O(N__39838),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIOJ9JZ0 ));
    InMux I__8374 (
            .O(N__39835),
            .I(N__39832));
    LocalMux I__8373 (
            .O(N__39832),
            .I(N__39829));
    Odrv12 I__8372 (
            .O(N__39829),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ));
    InMux I__8371 (
            .O(N__39826),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_23 ));
    InMux I__8370 (
            .O(N__39823),
            .I(N__39820));
    LocalMux I__8369 (
            .O(N__39820),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNIQMAJZ0 ));
    InMux I__8368 (
            .O(N__39817),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_24 ));
    InMux I__8367 (
            .O(N__39814),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_9 ));
    InMux I__8366 (
            .O(N__39811),
            .I(N__39808));
    LocalMux I__8365 (
            .O(N__39808),
            .I(\current_shift_inst.PI_CTRL.error_control_RNICE9PZ0Z_15 ));
    CascadeMux I__8364 (
            .O(N__39805),
            .I(N__39802));
    InMux I__8363 (
            .O(N__39802),
            .I(N__39799));
    LocalMux I__8362 (
            .O(N__39799),
            .I(\current_shift_inst.PI_CTRL.integrator_i_11 ));
    InMux I__8361 (
            .O(N__39796),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_10 ));
    InMux I__8360 (
            .O(N__39793),
            .I(N__39790));
    LocalMux I__8359 (
            .O(N__39790),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIGJAPZ0Z_16 ));
    InMux I__8358 (
            .O(N__39787),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_11 ));
    InMux I__8357 (
            .O(N__39784),
            .I(N__39781));
    LocalMux I__8356 (
            .O(N__39781),
            .I(N__39778));
    Span4Mux_h I__8355 (
            .O(N__39778),
            .I(N__39775));
    Odrv4 I__8354 (
            .O(N__39775),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ));
    InMux I__8353 (
            .O(N__39772),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_12 ));
    InMux I__8352 (
            .O(N__39769),
            .I(N__39766));
    LocalMux I__8351 (
            .O(N__39766),
            .I(N__39763));
    Span4Mux_h I__8350 (
            .O(N__39763),
            .I(N__39760));
    Odrv4 I__8349 (
            .O(N__39760),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ));
    InMux I__8348 (
            .O(N__39757),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_13 ));
    InMux I__8347 (
            .O(N__39754),
            .I(N__39751));
    LocalMux I__8346 (
            .O(N__39751),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIS2EPZ0Z_19 ));
    CascadeMux I__8345 (
            .O(N__39748),
            .I(N__39745));
    InMux I__8344 (
            .O(N__39745),
            .I(N__39742));
    LocalMux I__8343 (
            .O(N__39742),
            .I(N__39739));
    Odrv12 I__8342 (
            .O(N__39739),
            .I(\current_shift_inst.PI_CTRL.integrator_i_15 ));
    InMux I__8341 (
            .O(N__39736),
            .I(N__39733));
    LocalMux I__8340 (
            .O(N__39733),
            .I(N__39730));
    Span4Mux_h I__8339 (
            .O(N__39730),
            .I(N__39727));
    Odrv4 I__8338 (
            .O(N__39727),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ));
    InMux I__8337 (
            .O(N__39724),
            .I(bfn_16_10_0_));
    InMux I__8336 (
            .O(N__39721),
            .I(N__39718));
    LocalMux I__8335 (
            .O(N__39718),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIENGPZ0Z_20 ));
    CascadeMux I__8334 (
            .O(N__39715),
            .I(N__39712));
    InMux I__8333 (
            .O(N__39712),
            .I(N__39709));
    LocalMux I__8332 (
            .O(N__39709),
            .I(\current_shift_inst.PI_CTRL.integrator_i_16 ));
    InMux I__8331 (
            .O(N__39706),
            .I(N__39703));
    LocalMux I__8330 (
            .O(N__39703),
            .I(N__39700));
    Span4Mux_h I__8329 (
            .O(N__39700),
            .I(N__39697));
    Odrv4 I__8328 (
            .O(N__39697),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ));
    InMux I__8327 (
            .O(N__39694),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_15 ));
    CascadeMux I__8326 (
            .O(N__39691),
            .I(N__39688));
    InMux I__8325 (
            .O(N__39688),
            .I(N__39685));
    LocalMux I__8324 (
            .O(N__39685),
            .I(N__39682));
    Span4Mux_v I__8323 (
            .O(N__39682),
            .I(N__39679));
    Odrv4 I__8322 (
            .O(N__39679),
            .I(\current_shift_inst.PI_CTRL.integrator_i_17 ));
    InMux I__8321 (
            .O(N__39676),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_16 ));
    InMux I__8320 (
            .O(N__39673),
            .I(N__39670));
    LocalMux I__8319 (
            .O(N__39670),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIC46UZ0Z_6 ));
    CascadeMux I__8318 (
            .O(N__39667),
            .I(N__39664));
    InMux I__8317 (
            .O(N__39664),
            .I(N__39661));
    LocalMux I__8316 (
            .O(N__39661),
            .I(\current_shift_inst.PI_CTRL.integrator_i_2 ));
    InMux I__8315 (
            .O(N__39658),
            .I(N__39655));
    LocalMux I__8314 (
            .O(N__39655),
            .I(N__39652));
    Odrv4 I__8313 (
            .O(N__39652),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ));
    InMux I__8312 (
            .O(N__39649),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_1 ));
    InMux I__8311 (
            .O(N__39646),
            .I(N__39643));
    LocalMux I__8310 (
            .O(N__39643),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIG97UZ0Z_7 ));
    CascadeMux I__8309 (
            .O(N__39640),
            .I(N__39637));
    InMux I__8308 (
            .O(N__39637),
            .I(N__39634));
    LocalMux I__8307 (
            .O(N__39634),
            .I(\current_shift_inst.PI_CTRL.integrator_i_3 ));
    InMux I__8306 (
            .O(N__39631),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_2 ));
    InMux I__8305 (
            .O(N__39628),
            .I(N__39625));
    LocalMux I__8304 (
            .O(N__39625),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIKE8UZ0Z_8 ));
    CascadeMux I__8303 (
            .O(N__39622),
            .I(N__39619));
    InMux I__8302 (
            .O(N__39619),
            .I(N__39616));
    LocalMux I__8301 (
            .O(N__39616),
            .I(\current_shift_inst.PI_CTRL.integrator_i_4 ));
    InMux I__8300 (
            .O(N__39613),
            .I(N__39610));
    LocalMux I__8299 (
            .O(N__39610),
            .I(N__39607));
    Odrv4 I__8298 (
            .O(N__39607),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ));
    InMux I__8297 (
            .O(N__39604),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_3 ));
    InMux I__8296 (
            .O(N__39601),
            .I(N__39598));
    LocalMux I__8295 (
            .O(N__39598),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIOJ9UZ0Z_9 ));
    CascadeMux I__8294 (
            .O(N__39595),
            .I(N__39592));
    InMux I__8293 (
            .O(N__39592),
            .I(N__39589));
    LocalMux I__8292 (
            .O(N__39589),
            .I(N__39586));
    Span4Mux_h I__8291 (
            .O(N__39586),
            .I(N__39583));
    Odrv4 I__8290 (
            .O(N__39583),
            .I(\current_shift_inst.PI_CTRL.integrator_i_5 ));
    InMux I__8289 (
            .O(N__39580),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_4 ));
    InMux I__8288 (
            .O(N__39577),
            .I(N__39574));
    LocalMux I__8287 (
            .O(N__39574),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIA1B41Z0Z_10 ));
    CascadeMux I__8286 (
            .O(N__39571),
            .I(N__39568));
    InMux I__8285 (
            .O(N__39568),
            .I(N__39565));
    LocalMux I__8284 (
            .O(N__39565),
            .I(\current_shift_inst.PI_CTRL.integrator_i_6 ));
    InMux I__8283 (
            .O(N__39562),
            .I(N__39559));
    LocalMux I__8282 (
            .O(N__39559),
            .I(N__39556));
    Odrv12 I__8281 (
            .O(N__39556),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ));
    InMux I__8280 (
            .O(N__39553),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_5 ));
    InMux I__8279 (
            .O(N__39550),
            .I(N__39547));
    LocalMux I__8278 (
            .O(N__39547),
            .I(N__39544));
    Odrv4 I__8277 (
            .O(N__39544),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIL0S01Z0Z_11 ));
    InMux I__8276 (
            .O(N__39541),
            .I(bfn_16_9_0_));
    InMux I__8275 (
            .O(N__39538),
            .I(N__39535));
    LocalMux I__8274 (
            .O(N__39535),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIP5T01Z0Z_12 ));
    InMux I__8273 (
            .O(N__39532),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_7 ));
    InMux I__8272 (
            .O(N__39529),
            .I(N__39526));
    LocalMux I__8271 (
            .O(N__39526),
            .I(N__39523));
    Span4Mux_v I__8270 (
            .O(N__39523),
            .I(N__39520));
    Odrv4 I__8269 (
            .O(N__39520),
            .I(\current_shift_inst.PI_CTRL.error_control_RNITAU01Z0Z_13 ));
    CascadeMux I__8268 (
            .O(N__39517),
            .I(N__39514));
    InMux I__8267 (
            .O(N__39514),
            .I(N__39511));
    LocalMux I__8266 (
            .O(N__39511),
            .I(N__39508));
    Odrv4 I__8265 (
            .O(N__39508),
            .I(\current_shift_inst.PI_CTRL.integrator_i_9 ));
    InMux I__8264 (
            .O(N__39505),
            .I(N__39502));
    LocalMux I__8263 (
            .O(N__39502),
            .I(N__39499));
    Odrv4 I__8262 (
            .O(N__39499),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ));
    InMux I__8261 (
            .O(N__39496),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_8 ));
    CascadeMux I__8260 (
            .O(N__39493),
            .I(N__39488));
    CascadeMux I__8259 (
            .O(N__39492),
            .I(N__39485));
    InMux I__8258 (
            .O(N__39491),
            .I(N__39482));
    InMux I__8257 (
            .O(N__39488),
            .I(N__39479));
    InMux I__8256 (
            .O(N__39485),
            .I(N__39475));
    LocalMux I__8255 (
            .O(N__39482),
            .I(N__39472));
    LocalMux I__8254 (
            .O(N__39479),
            .I(N__39469));
    InMux I__8253 (
            .O(N__39478),
            .I(N__39466));
    LocalMux I__8252 (
            .O(N__39475),
            .I(N__39462));
    Span4Mux_h I__8251 (
            .O(N__39472),
            .I(N__39455));
    Span4Mux_v I__8250 (
            .O(N__39469),
            .I(N__39455));
    LocalMux I__8249 (
            .O(N__39466),
            .I(N__39455));
    InMux I__8248 (
            .O(N__39465),
            .I(N__39452));
    Span4Mux_v I__8247 (
            .O(N__39462),
            .I(N__39449));
    Span4Mux_v I__8246 (
            .O(N__39455),
            .I(N__39446));
    LocalMux I__8245 (
            .O(N__39452),
            .I(N__39443));
    Odrv4 I__8244 (
            .O(N__39449),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv4 I__8243 (
            .O(N__39446),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv4 I__8242 (
            .O(N__39443),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    InMux I__8241 (
            .O(N__39436),
            .I(N__39433));
    LocalMux I__8240 (
            .O(N__39433),
            .I(N__39429));
    InMux I__8239 (
            .O(N__39432),
            .I(N__39426));
    Span4Mux_v I__8238 (
            .O(N__39429),
            .I(N__39422));
    LocalMux I__8237 (
            .O(N__39426),
            .I(N__39419));
    InMux I__8236 (
            .O(N__39425),
            .I(N__39416));
    Span4Mux_h I__8235 (
            .O(N__39422),
            .I(N__39413));
    Span4Mux_h I__8234 (
            .O(N__39419),
            .I(N__39408));
    LocalMux I__8233 (
            .O(N__39416),
            .I(N__39408));
    Odrv4 I__8232 (
            .O(N__39413),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ));
    Odrv4 I__8231 (
            .O(N__39408),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ));
    CascadeMux I__8230 (
            .O(N__39403),
            .I(N__39399));
    InMux I__8229 (
            .O(N__39402),
            .I(N__39396));
    InMux I__8228 (
            .O(N__39399),
            .I(N__39393));
    LocalMux I__8227 (
            .O(N__39396),
            .I(N__39389));
    LocalMux I__8226 (
            .O(N__39393),
            .I(N__39386));
    CascadeMux I__8225 (
            .O(N__39392),
            .I(N__39383));
    Span4Mux_v I__8224 (
            .O(N__39389),
            .I(N__39378));
    Span4Mux_h I__8223 (
            .O(N__39386),
            .I(N__39378));
    InMux I__8222 (
            .O(N__39383),
            .I(N__39374));
    Span4Mux_h I__8221 (
            .O(N__39378),
            .I(N__39371));
    InMux I__8220 (
            .O(N__39377),
            .I(N__39368));
    LocalMux I__8219 (
            .O(N__39374),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    Odrv4 I__8218 (
            .O(N__39371),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    LocalMux I__8217 (
            .O(N__39368),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    CascadeMux I__8216 (
            .O(N__39361),
            .I(N__39357));
    InMux I__8215 (
            .O(N__39360),
            .I(N__39354));
    InMux I__8214 (
            .O(N__39357),
            .I(N__39350));
    LocalMux I__8213 (
            .O(N__39354),
            .I(N__39347));
    InMux I__8212 (
            .O(N__39353),
            .I(N__39344));
    LocalMux I__8211 (
            .O(N__39350),
            .I(N__39338));
    Span4Mux_h I__8210 (
            .O(N__39347),
            .I(N__39338));
    LocalMux I__8209 (
            .O(N__39344),
            .I(N__39335));
    InMux I__8208 (
            .O(N__39343),
            .I(N__39332));
    Span4Mux_h I__8207 (
            .O(N__39338),
            .I(N__39328));
    Span4Mux_h I__8206 (
            .O(N__39335),
            .I(N__39325));
    LocalMux I__8205 (
            .O(N__39332),
            .I(N__39322));
    InMux I__8204 (
            .O(N__39331),
            .I(N__39319));
    Odrv4 I__8203 (
            .O(N__39328),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    Odrv4 I__8202 (
            .O(N__39325),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    Odrv12 I__8201 (
            .O(N__39322),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    LocalMux I__8200 (
            .O(N__39319),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    CascadeMux I__8199 (
            .O(N__39310),
            .I(N__39306));
    InMux I__8198 (
            .O(N__39309),
            .I(N__39303));
    InMux I__8197 (
            .O(N__39306),
            .I(N__39300));
    LocalMux I__8196 (
            .O(N__39303),
            .I(N__39297));
    LocalMux I__8195 (
            .O(N__39300),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_i_26 ));
    Odrv4 I__8194 (
            .O(N__39297),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_i_26 ));
    InMux I__8193 (
            .O(N__39292),
            .I(N__39289));
    LocalMux I__8192 (
            .O(N__39289),
            .I(\current_shift_inst.PI_CTRL.error_control_RNI4Q3UZ0Z_4 ));
    CascadeMux I__8191 (
            .O(N__39286),
            .I(N__39282));
    CascadeMux I__8190 (
            .O(N__39285),
            .I(N__39279));
    InMux I__8189 (
            .O(N__39282),
            .I(N__39276));
    InMux I__8188 (
            .O(N__39279),
            .I(N__39273));
    LocalMux I__8187 (
            .O(N__39276),
            .I(\current_shift_inst.PI_CTRL.integrator_i_0 ));
    LocalMux I__8186 (
            .O(N__39273),
            .I(\current_shift_inst.PI_CTRL.integrator_i_0 ));
    InMux I__8185 (
            .O(N__39268),
            .I(N__39265));
    LocalMux I__8184 (
            .O(N__39265),
            .I(N__39262));
    Odrv4 I__8183 (
            .O(N__39262),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_0 ));
    InMux I__8182 (
            .O(N__39259),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO ));
    InMux I__8181 (
            .O(N__39256),
            .I(N__39253));
    LocalMux I__8180 (
            .O(N__39253),
            .I(\current_shift_inst.PI_CTRL.error_control_RNI8V4UZ0Z_5 ));
    CascadeMux I__8179 (
            .O(N__39250),
            .I(N__39247));
    InMux I__8178 (
            .O(N__39247),
            .I(N__39244));
    LocalMux I__8177 (
            .O(N__39244),
            .I(\current_shift_inst.PI_CTRL.integrator_i_1 ));
    InMux I__8176 (
            .O(N__39241),
            .I(N__39238));
    LocalMux I__8175 (
            .O(N__39238),
            .I(N__39235));
    Span4Mux_h I__8174 (
            .O(N__39235),
            .I(N__39232));
    Span4Mux_h I__8173 (
            .O(N__39232),
            .I(N__39229));
    Odrv4 I__8172 (
            .O(N__39229),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1 ));
    InMux I__8171 (
            .O(N__39226),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_0 ));
    IoInMux I__8170 (
            .O(N__39223),
            .I(N__39220));
    LocalMux I__8169 (
            .O(N__39220),
            .I(N__39217));
    Span4Mux_s1_v I__8168 (
            .O(N__39217),
            .I(N__39214));
    Span4Mux_h I__8167 (
            .O(N__39214),
            .I(N__39211));
    Odrv4 I__8166 (
            .O(N__39211),
            .I(\delay_measurement_inst.delay_tr_timer.N_304_i ));
    InMux I__8165 (
            .O(N__39208),
            .I(N__39203));
    InMux I__8164 (
            .O(N__39207),
            .I(N__39200));
    InMux I__8163 (
            .O(N__39206),
            .I(N__39197));
    LocalMux I__8162 (
            .O(N__39203),
            .I(\delay_measurement_inst.tr_stateZ0Z_0 ));
    LocalMux I__8161 (
            .O(N__39200),
            .I(\delay_measurement_inst.tr_stateZ0Z_0 ));
    LocalMux I__8160 (
            .O(N__39197),
            .I(\delay_measurement_inst.tr_stateZ0Z_0 ));
    InMux I__8159 (
            .O(N__39190),
            .I(N__39182));
    InMux I__8158 (
            .O(N__39189),
            .I(N__39182));
    InMux I__8157 (
            .O(N__39188),
            .I(N__39179));
    InMux I__8156 (
            .O(N__39187),
            .I(N__39176));
    LocalMux I__8155 (
            .O(N__39182),
            .I(delay_tr_d2));
    LocalMux I__8154 (
            .O(N__39179),
            .I(delay_tr_d2));
    LocalMux I__8153 (
            .O(N__39176),
            .I(delay_tr_d2));
    InMux I__8152 (
            .O(N__39169),
            .I(N__39164));
    InMux I__8151 (
            .O(N__39168),
            .I(N__39161));
    InMux I__8150 (
            .O(N__39167),
            .I(N__39158));
    LocalMux I__8149 (
            .O(N__39164),
            .I(\delay_measurement_inst.prev_tr_sigZ0 ));
    LocalMux I__8148 (
            .O(N__39161),
            .I(\delay_measurement_inst.prev_tr_sigZ0 ));
    LocalMux I__8147 (
            .O(N__39158),
            .I(\delay_measurement_inst.prev_tr_sigZ0 ));
    InMux I__8146 (
            .O(N__39151),
            .I(N__39147));
    InMux I__8145 (
            .O(N__39150),
            .I(N__39144));
    LocalMux I__8144 (
            .O(N__39147),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    LocalMux I__8143 (
            .O(N__39144),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    InMux I__8142 (
            .O(N__39139),
            .I(N__39135));
    InMux I__8141 (
            .O(N__39138),
            .I(N__39131));
    LocalMux I__8140 (
            .O(N__39135),
            .I(N__39128));
    InMux I__8139 (
            .O(N__39134),
            .I(N__39125));
    LocalMux I__8138 (
            .O(N__39131),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    Odrv4 I__8137 (
            .O(N__39128),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    LocalMux I__8136 (
            .O(N__39125),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    InMux I__8135 (
            .O(N__39118),
            .I(N__39112));
    InMux I__8134 (
            .O(N__39117),
            .I(N__39107));
    InMux I__8133 (
            .O(N__39116),
            .I(N__39107));
    InMux I__8132 (
            .O(N__39115),
            .I(N__39104));
    LocalMux I__8131 (
            .O(N__39112),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    LocalMux I__8130 (
            .O(N__39107),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    LocalMux I__8129 (
            .O(N__39104),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    InMux I__8128 (
            .O(N__39097),
            .I(N__39094));
    LocalMux I__8127 (
            .O(N__39094),
            .I(N__39091));
    Span4Mux_h I__8126 (
            .O(N__39091),
            .I(N__39088));
    Odrv4 I__8125 (
            .O(N__39088),
            .I(\current_shift_inst.un38_control_input_0_s1_29 ));
    InMux I__8124 (
            .O(N__39085),
            .I(\current_shift_inst.un38_control_input_cry_28_s1 ));
    InMux I__8123 (
            .O(N__39082),
            .I(N__39079));
    LocalMux I__8122 (
            .O(N__39079),
            .I(N__39076));
    Span4Mux_v I__8121 (
            .O(N__39076),
            .I(N__39073));
    Odrv4 I__8120 (
            .O(N__39073),
            .I(\current_shift_inst.un38_control_input_0_s1_30 ));
    InMux I__8119 (
            .O(N__39070),
            .I(\current_shift_inst.un38_control_input_cry_29_s1 ));
    InMux I__8118 (
            .O(N__39067),
            .I(\current_shift_inst.un38_control_input_cry_30_s1 ));
    InMux I__8117 (
            .O(N__39064),
            .I(N__39061));
    LocalMux I__8116 (
            .O(N__39061),
            .I(N__39058));
    Span4Mux_h I__8115 (
            .O(N__39058),
            .I(N__39055));
    Odrv4 I__8114 (
            .O(N__39055),
            .I(\current_shift_inst.un38_control_input_0_s1_31 ));
    InMux I__8113 (
            .O(N__39052),
            .I(N__39049));
    LocalMux I__8112 (
            .O(N__39049),
            .I(N__39044));
    InMux I__8111 (
            .O(N__39048),
            .I(N__39041));
    CascadeMux I__8110 (
            .O(N__39047),
            .I(N__39038));
    Span4Mux_h I__8109 (
            .O(N__39044),
            .I(N__39035));
    LocalMux I__8108 (
            .O(N__39041),
            .I(N__39032));
    InMux I__8107 (
            .O(N__39038),
            .I(N__39029));
    Odrv4 I__8106 (
            .O(N__39035),
            .I(\delay_measurement_inst.elapsed_time_hc_18 ));
    Odrv4 I__8105 (
            .O(N__39032),
            .I(\delay_measurement_inst.elapsed_time_hc_18 ));
    LocalMux I__8104 (
            .O(N__39029),
            .I(\delay_measurement_inst.elapsed_time_hc_18 ));
    InMux I__8103 (
            .O(N__39022),
            .I(N__39019));
    LocalMux I__8102 (
            .O(N__39019),
            .I(N__39014));
    InMux I__8101 (
            .O(N__39018),
            .I(N__39011));
    InMux I__8100 (
            .O(N__39017),
            .I(N__39008));
    Span4Mux_h I__8099 (
            .O(N__39014),
            .I(N__39005));
    LocalMux I__8098 (
            .O(N__39011),
            .I(N__39002));
    LocalMux I__8097 (
            .O(N__39008),
            .I(N__38999));
    Odrv4 I__8096 (
            .O(N__39005),
            .I(\delay_measurement_inst.elapsed_time_hc_17 ));
    Odrv4 I__8095 (
            .O(N__39002),
            .I(\delay_measurement_inst.elapsed_time_hc_17 ));
    Odrv4 I__8094 (
            .O(N__38999),
            .I(\delay_measurement_inst.elapsed_time_hc_17 ));
    InMux I__8093 (
            .O(N__38992),
            .I(N__38988));
    CascadeMux I__8092 (
            .O(N__38991),
            .I(N__38985));
    LocalMux I__8091 (
            .O(N__38988),
            .I(N__38982));
    InMux I__8090 (
            .O(N__38985),
            .I(N__38979));
    Span4Mux_v I__8089 (
            .O(N__38982),
            .I(N__38975));
    LocalMux I__8088 (
            .O(N__38979),
            .I(N__38972));
    InMux I__8087 (
            .O(N__38978),
            .I(N__38969));
    Odrv4 I__8086 (
            .O(N__38975),
            .I(\delay_measurement_inst.elapsed_time_hc_16 ));
    Odrv4 I__8085 (
            .O(N__38972),
            .I(\delay_measurement_inst.elapsed_time_hc_16 ));
    LocalMux I__8084 (
            .O(N__38969),
            .I(\delay_measurement_inst.elapsed_time_hc_16 ));
    CascadeMux I__8083 (
            .O(N__38962),
            .I(N__38957));
    InMux I__8082 (
            .O(N__38961),
            .I(N__38954));
    InMux I__8081 (
            .O(N__38960),
            .I(N__38951));
    InMux I__8080 (
            .O(N__38957),
            .I(N__38948));
    LocalMux I__8079 (
            .O(N__38954),
            .I(N__38945));
    LocalMux I__8078 (
            .O(N__38951),
            .I(N__38940));
    LocalMux I__8077 (
            .O(N__38948),
            .I(N__38940));
    Odrv4 I__8076 (
            .O(N__38945),
            .I(\delay_measurement_inst.elapsed_time_hc_19 ));
    Odrv4 I__8075 (
            .O(N__38940),
            .I(\delay_measurement_inst.elapsed_time_hc_19 ));
    InMux I__8074 (
            .O(N__38935),
            .I(N__38931));
    InMux I__8073 (
            .O(N__38934),
            .I(N__38928));
    LocalMux I__8072 (
            .O(N__38931),
            .I(N__38925));
    LocalMux I__8071 (
            .O(N__38928),
            .I(N__38922));
    Span4Mux_h I__8070 (
            .O(N__38925),
            .I(N__38919));
    Span4Mux_h I__8069 (
            .O(N__38922),
            .I(N__38916));
    Odrv4 I__8068 (
            .O(N__38919),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_1 ));
    Odrv4 I__8067 (
            .O(N__38916),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_1 ));
    InMux I__8066 (
            .O(N__38911),
            .I(N__38908));
    LocalMux I__8065 (
            .O(N__38908),
            .I(N__38905));
    Span4Mux_h I__8064 (
            .O(N__38905),
            .I(N__38901));
    InMux I__8063 (
            .O(N__38904),
            .I(N__38898));
    Span4Mux_v I__8062 (
            .O(N__38901),
            .I(N__38894));
    LocalMux I__8061 (
            .O(N__38898),
            .I(N__38891));
    InMux I__8060 (
            .O(N__38897),
            .I(N__38888));
    Odrv4 I__8059 (
            .O(N__38894),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    Odrv12 I__8058 (
            .O(N__38891),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__8057 (
            .O(N__38888),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    InMux I__8056 (
            .O(N__38881),
            .I(N__38878));
    LocalMux I__8055 (
            .O(N__38878),
            .I(N__38874));
    InMux I__8054 (
            .O(N__38877),
            .I(N__38871));
    Span4Mux_v I__8053 (
            .O(N__38874),
            .I(N__38866));
    LocalMux I__8052 (
            .O(N__38871),
            .I(N__38866));
    Odrv4 I__8051 (
            .O(N__38866),
            .I(\delay_measurement_inst.elapsed_time_hc_1 ));
    InMux I__8050 (
            .O(N__38863),
            .I(N__38860));
    LocalMux I__8049 (
            .O(N__38860),
            .I(N__38856));
    InMux I__8048 (
            .O(N__38859),
            .I(N__38853));
    Span4Mux_v I__8047 (
            .O(N__38856),
            .I(N__38849));
    LocalMux I__8046 (
            .O(N__38853),
            .I(N__38846));
    InMux I__8045 (
            .O(N__38852),
            .I(N__38843));
    Odrv4 I__8044 (
            .O(N__38849),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    Odrv12 I__8043 (
            .O(N__38846),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    LocalMux I__8042 (
            .O(N__38843),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    InMux I__8041 (
            .O(N__38836),
            .I(N__38833));
    LocalMux I__8040 (
            .O(N__38833),
            .I(N__38828));
    InMux I__8039 (
            .O(N__38832),
            .I(N__38825));
    InMux I__8038 (
            .O(N__38831),
            .I(N__38822));
    Span4Mux_v I__8037 (
            .O(N__38828),
            .I(N__38817));
    LocalMux I__8036 (
            .O(N__38825),
            .I(N__38817));
    LocalMux I__8035 (
            .O(N__38822),
            .I(\delay_measurement_inst.elapsed_time_hc_2 ));
    Odrv4 I__8034 (
            .O(N__38817),
            .I(\delay_measurement_inst.elapsed_time_hc_2 ));
    CEMux I__8033 (
            .O(N__38812),
            .I(N__38797));
    CEMux I__8032 (
            .O(N__38811),
            .I(N__38797));
    CEMux I__8031 (
            .O(N__38810),
            .I(N__38797));
    CEMux I__8030 (
            .O(N__38809),
            .I(N__38797));
    CEMux I__8029 (
            .O(N__38808),
            .I(N__38797));
    GlobalMux I__8028 (
            .O(N__38797),
            .I(N__38794));
    gio2CtrlBuf I__8027 (
            .O(N__38794),
            .I(\delay_measurement_inst.delay_hc_timer.N_302_i_g ));
    CascadeMux I__8026 (
            .O(N__38791),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_3_cascade_ ));
    InMux I__8025 (
            .O(N__38788),
            .I(N__38785));
    LocalMux I__8024 (
            .O(N__38785),
            .I(N__38782));
    Odrv4 I__8023 (
            .O(N__38782),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_4 ));
    InMux I__8022 (
            .O(N__38779),
            .I(N__38773));
    InMux I__8021 (
            .O(N__38778),
            .I(N__38770));
    InMux I__8020 (
            .O(N__38777),
            .I(N__38767));
    InMux I__8019 (
            .O(N__38776),
            .I(N__38764));
    LocalMux I__8018 (
            .O(N__38773),
            .I(N__38757));
    LocalMux I__8017 (
            .O(N__38770),
            .I(N__38757));
    LocalMux I__8016 (
            .O(N__38767),
            .I(N__38757));
    LocalMux I__8015 (
            .O(N__38764),
            .I(N__38754));
    Span4Mux_v I__8014 (
            .O(N__38757),
            .I(N__38751));
    Span4Mux_h I__8013 (
            .O(N__38754),
            .I(N__38748));
    Span4Mux_h I__8012 (
            .O(N__38751),
            .I(N__38745));
    Span4Mux_v I__8011 (
            .O(N__38748),
            .I(N__38742));
    Odrv4 I__8010 (
            .O(N__38745),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto30Z0Z_1 ));
    Odrv4 I__8009 (
            .O(N__38742),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto30Z0Z_1 ));
    InMux I__8008 (
            .O(N__38737),
            .I(\current_shift_inst.un38_control_input_cry_19_s1 ));
    InMux I__8007 (
            .O(N__38734),
            .I(N__38731));
    LocalMux I__8006 (
            .O(N__38731),
            .I(N__38728));
    Span4Mux_h I__8005 (
            .O(N__38728),
            .I(N__38725));
    Span4Mux_v I__8004 (
            .O(N__38725),
            .I(N__38722));
    Odrv4 I__8003 (
            .O(N__38722),
            .I(\current_shift_inst.un38_control_input_0_s1_21 ));
    InMux I__8002 (
            .O(N__38719),
            .I(\current_shift_inst.un38_control_input_cry_20_s1 ));
    InMux I__8001 (
            .O(N__38716),
            .I(N__38713));
    LocalMux I__8000 (
            .O(N__38713),
            .I(N__38710));
    Span4Mux_h I__7999 (
            .O(N__38710),
            .I(N__38707));
    Odrv4 I__7998 (
            .O(N__38707),
            .I(\current_shift_inst.un38_control_input_0_s1_22 ));
    InMux I__7997 (
            .O(N__38704),
            .I(\current_shift_inst.un38_control_input_cry_21_s1 ));
    InMux I__7996 (
            .O(N__38701),
            .I(N__38698));
    LocalMux I__7995 (
            .O(N__38698),
            .I(N__38695));
    Span4Mux_h I__7994 (
            .O(N__38695),
            .I(N__38692));
    Span4Mux_v I__7993 (
            .O(N__38692),
            .I(N__38689));
    Odrv4 I__7992 (
            .O(N__38689),
            .I(\current_shift_inst.un38_control_input_0_s1_23 ));
    InMux I__7991 (
            .O(N__38686),
            .I(\current_shift_inst.un38_control_input_cry_22_s1 ));
    InMux I__7990 (
            .O(N__38683),
            .I(N__38680));
    LocalMux I__7989 (
            .O(N__38680),
            .I(N__38677));
    Span4Mux_h I__7988 (
            .O(N__38677),
            .I(N__38674));
    Odrv4 I__7987 (
            .O(N__38674),
            .I(\current_shift_inst.un38_control_input_0_s1_24 ));
    InMux I__7986 (
            .O(N__38671),
            .I(bfn_15_22_0_));
    InMux I__7985 (
            .O(N__38668),
            .I(N__38665));
    LocalMux I__7984 (
            .O(N__38665),
            .I(N__38662));
    Odrv4 I__7983 (
            .O(N__38662),
            .I(\current_shift_inst.un38_control_input_0_s1_25 ));
    InMux I__7982 (
            .O(N__38659),
            .I(\current_shift_inst.un38_control_input_cry_24_s1 ));
    InMux I__7981 (
            .O(N__38656),
            .I(N__38653));
    LocalMux I__7980 (
            .O(N__38653),
            .I(N__38650));
    Odrv4 I__7979 (
            .O(N__38650),
            .I(\current_shift_inst.un38_control_input_0_s1_26 ));
    InMux I__7978 (
            .O(N__38647),
            .I(\current_shift_inst.un38_control_input_cry_25_s1 ));
    CascadeMux I__7977 (
            .O(N__38644),
            .I(N__38641));
    InMux I__7976 (
            .O(N__38641),
            .I(N__38638));
    LocalMux I__7975 (
            .O(N__38638),
            .I(N__38635));
    Odrv4 I__7974 (
            .O(N__38635),
            .I(\current_shift_inst.un38_control_input_0_s1_27 ));
    InMux I__7973 (
            .O(N__38632),
            .I(\current_shift_inst.un38_control_input_cry_26_s1 ));
    InMux I__7972 (
            .O(N__38629),
            .I(N__38626));
    LocalMux I__7971 (
            .O(N__38626),
            .I(N__38623));
    Span4Mux_h I__7970 (
            .O(N__38623),
            .I(N__38620));
    Odrv4 I__7969 (
            .O(N__38620),
            .I(\current_shift_inst.un38_control_input_0_s1_28 ));
    InMux I__7968 (
            .O(N__38617),
            .I(\current_shift_inst.un38_control_input_cry_27_s1 ));
    InMux I__7967 (
            .O(N__38614),
            .I(N__38611));
    LocalMux I__7966 (
            .O(N__38611),
            .I(N__38608));
    Span4Mux_h I__7965 (
            .O(N__38608),
            .I(N__38605));
    Span4Mux_v I__7964 (
            .O(N__38605),
            .I(N__38602));
    Odrv4 I__7963 (
            .O(N__38602),
            .I(\current_shift_inst.un38_control_input_0_s1_12 ));
    InMux I__7962 (
            .O(N__38599),
            .I(\current_shift_inst.un38_control_input_cry_11_s1 ));
    InMux I__7961 (
            .O(N__38596),
            .I(\current_shift_inst.un38_control_input_cry_12_s1 ));
    InMux I__7960 (
            .O(N__38593),
            .I(N__38590));
    LocalMux I__7959 (
            .O(N__38590),
            .I(N__38587));
    Span4Mux_h I__7958 (
            .O(N__38587),
            .I(N__38584));
    Span4Mux_v I__7957 (
            .O(N__38584),
            .I(N__38581));
    Odrv4 I__7956 (
            .O(N__38581),
            .I(\current_shift_inst.un38_control_input_0_s1_14 ));
    InMux I__7955 (
            .O(N__38578),
            .I(\current_shift_inst.un38_control_input_cry_13_s1 ));
    InMux I__7954 (
            .O(N__38575),
            .I(N__38572));
    LocalMux I__7953 (
            .O(N__38572),
            .I(N__38569));
    Span4Mux_h I__7952 (
            .O(N__38569),
            .I(N__38566));
    Span4Mux_v I__7951 (
            .O(N__38566),
            .I(N__38563));
    Odrv4 I__7950 (
            .O(N__38563),
            .I(\current_shift_inst.un38_control_input_0_s1_15 ));
    InMux I__7949 (
            .O(N__38560),
            .I(\current_shift_inst.un38_control_input_cry_14_s1 ));
    InMux I__7948 (
            .O(N__38557),
            .I(N__38554));
    LocalMux I__7947 (
            .O(N__38554),
            .I(N__38551));
    Span4Mux_h I__7946 (
            .O(N__38551),
            .I(N__38548));
    Span4Mux_v I__7945 (
            .O(N__38548),
            .I(N__38545));
    Odrv4 I__7944 (
            .O(N__38545),
            .I(\current_shift_inst.un38_control_input_0_s1_16 ));
    InMux I__7943 (
            .O(N__38542),
            .I(bfn_15_21_0_));
    InMux I__7942 (
            .O(N__38539),
            .I(N__38536));
    LocalMux I__7941 (
            .O(N__38536),
            .I(N__38533));
    Span4Mux_h I__7940 (
            .O(N__38533),
            .I(N__38530));
    Span4Mux_v I__7939 (
            .O(N__38530),
            .I(N__38527));
    Odrv4 I__7938 (
            .O(N__38527),
            .I(\current_shift_inst.un38_control_input_0_s1_17 ));
    InMux I__7937 (
            .O(N__38524),
            .I(\current_shift_inst.un38_control_input_cry_16_s1 ));
    InMux I__7936 (
            .O(N__38521),
            .I(N__38518));
    LocalMux I__7935 (
            .O(N__38518),
            .I(N__38515));
    Span4Mux_v I__7934 (
            .O(N__38515),
            .I(N__38512));
    Span4Mux_v I__7933 (
            .O(N__38512),
            .I(N__38509));
    Odrv4 I__7932 (
            .O(N__38509),
            .I(\current_shift_inst.un38_control_input_0_s1_18 ));
    InMux I__7931 (
            .O(N__38506),
            .I(\current_shift_inst.un38_control_input_cry_17_s1 ));
    InMux I__7930 (
            .O(N__38503),
            .I(N__38500));
    LocalMux I__7929 (
            .O(N__38500),
            .I(N__38497));
    Span4Mux_h I__7928 (
            .O(N__38497),
            .I(N__38494));
    Span4Mux_v I__7927 (
            .O(N__38494),
            .I(N__38491));
    Odrv4 I__7926 (
            .O(N__38491),
            .I(\current_shift_inst.un38_control_input_0_s1_19 ));
    InMux I__7925 (
            .O(N__38488),
            .I(\current_shift_inst.un38_control_input_cry_18_s1 ));
    InMux I__7924 (
            .O(N__38485),
            .I(N__38482));
    LocalMux I__7923 (
            .O(N__38482),
            .I(N__38479));
    Span4Mux_h I__7922 (
            .O(N__38479),
            .I(N__38476));
    Span4Mux_v I__7921 (
            .O(N__38476),
            .I(N__38473));
    Odrv4 I__7920 (
            .O(N__38473),
            .I(\current_shift_inst.un38_control_input_0_s1_20 ));
    InMux I__7919 (
            .O(N__38470),
            .I(N__38467));
    LocalMux I__7918 (
            .O(N__38467),
            .I(\current_shift_inst.un38_control_input_0_s1_6 ));
    InMux I__7917 (
            .O(N__38464),
            .I(\current_shift_inst.un38_control_input_cry_5_s1 ));
    InMux I__7916 (
            .O(N__38461),
            .I(N__38458));
    LocalMux I__7915 (
            .O(N__38458),
            .I(N__38455));
    Odrv4 I__7914 (
            .O(N__38455),
            .I(\current_shift_inst.un38_control_input_0_s1_7 ));
    InMux I__7913 (
            .O(N__38452),
            .I(\current_shift_inst.un38_control_input_cry_6_s1 ));
    InMux I__7912 (
            .O(N__38449),
            .I(N__38446));
    LocalMux I__7911 (
            .O(N__38446),
            .I(N__38443));
    Span4Mux_h I__7910 (
            .O(N__38443),
            .I(N__38440));
    Odrv4 I__7909 (
            .O(N__38440),
            .I(\current_shift_inst.un38_control_input_0_s1_8 ));
    InMux I__7908 (
            .O(N__38437),
            .I(bfn_15_20_0_));
    InMux I__7907 (
            .O(N__38434),
            .I(N__38431));
    LocalMux I__7906 (
            .O(N__38431),
            .I(N__38428));
    Span4Mux_h I__7905 (
            .O(N__38428),
            .I(N__38425));
    Odrv4 I__7904 (
            .O(N__38425),
            .I(\current_shift_inst.un38_control_input_0_s1_9 ));
    InMux I__7903 (
            .O(N__38422),
            .I(\current_shift_inst.un38_control_input_cry_8_s1 ));
    InMux I__7902 (
            .O(N__38419),
            .I(N__38416));
    LocalMux I__7901 (
            .O(N__38416),
            .I(N__38413));
    Span4Mux_h I__7900 (
            .O(N__38413),
            .I(N__38410));
    Span4Mux_v I__7899 (
            .O(N__38410),
            .I(N__38407));
    Odrv4 I__7898 (
            .O(N__38407),
            .I(\current_shift_inst.un38_control_input_0_s1_10 ));
    InMux I__7897 (
            .O(N__38404),
            .I(\current_shift_inst.un38_control_input_cry_9_s1 ));
    InMux I__7896 (
            .O(N__38401),
            .I(\current_shift_inst.un38_control_input_cry_10_s1 ));
    InMux I__7895 (
            .O(N__38398),
            .I(N__38395));
    LocalMux I__7894 (
            .O(N__38395),
            .I(N__38369));
    InMux I__7893 (
            .O(N__38394),
            .I(N__38355));
    InMux I__7892 (
            .O(N__38393),
            .I(N__38355));
    InMux I__7891 (
            .O(N__38392),
            .I(N__38355));
    InMux I__7890 (
            .O(N__38391),
            .I(N__38346));
    InMux I__7889 (
            .O(N__38390),
            .I(N__38346));
    InMux I__7888 (
            .O(N__38389),
            .I(N__38346));
    InMux I__7887 (
            .O(N__38388),
            .I(N__38346));
    CascadeMux I__7886 (
            .O(N__38387),
            .I(N__38343));
    CascadeMux I__7885 (
            .O(N__38386),
            .I(N__38340));
    CascadeMux I__7884 (
            .O(N__38385),
            .I(N__38336));
    CascadeMux I__7883 (
            .O(N__38384),
            .I(N__38333));
    CascadeMux I__7882 (
            .O(N__38383),
            .I(N__38330));
    CascadeMux I__7881 (
            .O(N__38382),
            .I(N__38327));
    CascadeMux I__7880 (
            .O(N__38381),
            .I(N__38323));
    CascadeMux I__7879 (
            .O(N__38380),
            .I(N__38320));
    CascadeMux I__7878 (
            .O(N__38379),
            .I(N__38317));
    CascadeMux I__7877 (
            .O(N__38378),
            .I(N__38314));
    CascadeMux I__7876 (
            .O(N__38377),
            .I(N__38311));
    CascadeMux I__7875 (
            .O(N__38376),
            .I(N__38308));
    CascadeMux I__7874 (
            .O(N__38375),
            .I(N__38305));
    CascadeMux I__7873 (
            .O(N__38374),
            .I(N__38302));
    CascadeMux I__7872 (
            .O(N__38373),
            .I(N__38299));
    CascadeMux I__7871 (
            .O(N__38372),
            .I(N__38296));
    Span4Mux_s2_h I__7870 (
            .O(N__38369),
            .I(N__38276));
    InMux I__7869 (
            .O(N__38368),
            .I(N__38269));
    InMux I__7868 (
            .O(N__38367),
            .I(N__38269));
    InMux I__7867 (
            .O(N__38366),
            .I(N__38269));
    InMux I__7866 (
            .O(N__38365),
            .I(N__38260));
    InMux I__7865 (
            .O(N__38364),
            .I(N__38260));
    InMux I__7864 (
            .O(N__38363),
            .I(N__38260));
    InMux I__7863 (
            .O(N__38362),
            .I(N__38260));
    LocalMux I__7862 (
            .O(N__38355),
            .I(N__38255));
    LocalMux I__7861 (
            .O(N__38346),
            .I(N__38255));
    InMux I__7860 (
            .O(N__38343),
            .I(N__38252));
    InMux I__7859 (
            .O(N__38340),
            .I(N__38247));
    InMux I__7858 (
            .O(N__38339),
            .I(N__38247));
    InMux I__7857 (
            .O(N__38336),
            .I(N__38242));
    InMux I__7856 (
            .O(N__38333),
            .I(N__38242));
    InMux I__7855 (
            .O(N__38330),
            .I(N__38231));
    InMux I__7854 (
            .O(N__38327),
            .I(N__38231));
    InMux I__7853 (
            .O(N__38326),
            .I(N__38231));
    InMux I__7852 (
            .O(N__38323),
            .I(N__38231));
    InMux I__7851 (
            .O(N__38320),
            .I(N__38231));
    InMux I__7850 (
            .O(N__38317),
            .I(N__38222));
    InMux I__7849 (
            .O(N__38314),
            .I(N__38222));
    InMux I__7848 (
            .O(N__38311),
            .I(N__38222));
    InMux I__7847 (
            .O(N__38308),
            .I(N__38222));
    InMux I__7846 (
            .O(N__38305),
            .I(N__38213));
    InMux I__7845 (
            .O(N__38302),
            .I(N__38213));
    InMux I__7844 (
            .O(N__38299),
            .I(N__38213));
    InMux I__7843 (
            .O(N__38296),
            .I(N__38213));
    CascadeMux I__7842 (
            .O(N__38295),
            .I(N__38210));
    CascadeMux I__7841 (
            .O(N__38294),
            .I(N__38207));
    CascadeMux I__7840 (
            .O(N__38293),
            .I(N__38204));
    CascadeMux I__7839 (
            .O(N__38292),
            .I(N__38201));
    CascadeMux I__7838 (
            .O(N__38291),
            .I(N__38197));
    CascadeMux I__7837 (
            .O(N__38290),
            .I(N__38194));
    CascadeMux I__7836 (
            .O(N__38289),
            .I(N__38191));
    InMux I__7835 (
            .O(N__38288),
            .I(N__38188));
    InMux I__7834 (
            .O(N__38287),
            .I(N__38185));
    CascadeMux I__7833 (
            .O(N__38286),
            .I(N__38182));
    CascadeMux I__7832 (
            .O(N__38285),
            .I(N__38179));
    CascadeMux I__7831 (
            .O(N__38284),
            .I(N__38176));
    CascadeMux I__7830 (
            .O(N__38283),
            .I(N__38173));
    CascadeMux I__7829 (
            .O(N__38282),
            .I(N__38170));
    CascadeMux I__7828 (
            .O(N__38281),
            .I(N__38167));
    CascadeMux I__7827 (
            .O(N__38280),
            .I(N__38164));
    InMux I__7826 (
            .O(N__38279),
            .I(N__38159));
    Span4Mux_h I__7825 (
            .O(N__38276),
            .I(N__38156));
    LocalMux I__7824 (
            .O(N__38269),
            .I(N__38151));
    LocalMux I__7823 (
            .O(N__38260),
            .I(N__38151));
    Span4Mux_s3_h I__7822 (
            .O(N__38255),
            .I(N__38148));
    LocalMux I__7821 (
            .O(N__38252),
            .I(N__38143));
    LocalMux I__7820 (
            .O(N__38247),
            .I(N__38143));
    LocalMux I__7819 (
            .O(N__38242),
            .I(N__38134));
    LocalMux I__7818 (
            .O(N__38231),
            .I(N__38134));
    LocalMux I__7817 (
            .O(N__38222),
            .I(N__38134));
    LocalMux I__7816 (
            .O(N__38213),
            .I(N__38134));
    InMux I__7815 (
            .O(N__38210),
            .I(N__38127));
    InMux I__7814 (
            .O(N__38207),
            .I(N__38127));
    InMux I__7813 (
            .O(N__38204),
            .I(N__38127));
    InMux I__7812 (
            .O(N__38201),
            .I(N__38116));
    InMux I__7811 (
            .O(N__38200),
            .I(N__38116));
    InMux I__7810 (
            .O(N__38197),
            .I(N__38116));
    InMux I__7809 (
            .O(N__38194),
            .I(N__38116));
    InMux I__7808 (
            .O(N__38191),
            .I(N__38116));
    LocalMux I__7807 (
            .O(N__38188),
            .I(N__38113));
    LocalMux I__7806 (
            .O(N__38185),
            .I(N__38110));
    InMux I__7805 (
            .O(N__38182),
            .I(N__38103));
    InMux I__7804 (
            .O(N__38179),
            .I(N__38103));
    InMux I__7803 (
            .O(N__38176),
            .I(N__38103));
    InMux I__7802 (
            .O(N__38173),
            .I(N__38094));
    InMux I__7801 (
            .O(N__38170),
            .I(N__38094));
    InMux I__7800 (
            .O(N__38167),
            .I(N__38094));
    InMux I__7799 (
            .O(N__38164),
            .I(N__38094));
    InMux I__7798 (
            .O(N__38163),
            .I(N__38091));
    InMux I__7797 (
            .O(N__38162),
            .I(N__38088));
    LocalMux I__7796 (
            .O(N__38159),
            .I(N__38083));
    Span4Mux_v I__7795 (
            .O(N__38156),
            .I(N__38078));
    Span4Mux_s2_h I__7794 (
            .O(N__38151),
            .I(N__38078));
    Span4Mux_v I__7793 (
            .O(N__38148),
            .I(N__38073));
    Span4Mux_s3_h I__7792 (
            .O(N__38143),
            .I(N__38073));
    Span4Mux_v I__7791 (
            .O(N__38134),
            .I(N__38070));
    LocalMux I__7790 (
            .O(N__38127),
            .I(N__38065));
    LocalMux I__7789 (
            .O(N__38116),
            .I(N__38065));
    Span4Mux_v I__7788 (
            .O(N__38113),
            .I(N__38060));
    Span4Mux_v I__7787 (
            .O(N__38110),
            .I(N__38060));
    LocalMux I__7786 (
            .O(N__38103),
            .I(N__38055));
    LocalMux I__7785 (
            .O(N__38094),
            .I(N__38055));
    LocalMux I__7784 (
            .O(N__38091),
            .I(N__38052));
    LocalMux I__7783 (
            .O(N__38088),
            .I(N__38049));
    InMux I__7782 (
            .O(N__38087),
            .I(N__38046));
    InMux I__7781 (
            .O(N__38086),
            .I(N__38043));
    Span12Mux_s2_h I__7780 (
            .O(N__38083),
            .I(N__38038));
    Sp12to4 I__7779 (
            .O(N__38078),
            .I(N__38038));
    Sp12to4 I__7778 (
            .O(N__38073),
            .I(N__38035));
    Sp12to4 I__7777 (
            .O(N__38070),
            .I(N__38028));
    Span12Mux_s10_h I__7776 (
            .O(N__38065),
            .I(N__38028));
    Sp12to4 I__7775 (
            .O(N__38060),
            .I(N__38028));
    Span12Mux_v I__7774 (
            .O(N__38055),
            .I(N__38023));
    Span12Mux_s10_h I__7773 (
            .O(N__38052),
            .I(N__38023));
    Span4Mux_s3_h I__7772 (
            .O(N__38049),
            .I(N__38020));
    LocalMux I__7771 (
            .O(N__38046),
            .I(N__38015));
    LocalMux I__7770 (
            .O(N__38043),
            .I(N__38015));
    Span12Mux_v I__7769 (
            .O(N__38038),
            .I(N__38012));
    Span12Mux_v I__7768 (
            .O(N__38035),
            .I(N__38001));
    Span12Mux_h I__7767 (
            .O(N__38028),
            .I(N__38001));
    Span12Mux_h I__7766 (
            .O(N__38023),
            .I(N__38001));
    Sp12to4 I__7765 (
            .O(N__38020),
            .I(N__38001));
    Span12Mux_s3_h I__7764 (
            .O(N__38015),
            .I(N__38001));
    Odrv12 I__7763 (
            .O(N__38012),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__7762 (
            .O(N__38001),
            .I(CONSTANT_ONE_NET));
    InMux I__7761 (
            .O(N__37996),
            .I(\current_shift_inst.un10_control_input_cry_30 ));
    InMux I__7760 (
            .O(N__37993),
            .I(N__37989));
    InMux I__7759 (
            .O(N__37992),
            .I(N__37986));
    LocalMux I__7758 (
            .O(N__37989),
            .I(N__37983));
    LocalMux I__7757 (
            .O(N__37986),
            .I(N__37978));
    Span4Mux_h I__7756 (
            .O(N__37983),
            .I(N__37978));
    Odrv4 I__7755 (
            .O(N__37978),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    CascadeMux I__7754 (
            .O(N__37975),
            .I(N__37971));
    CascadeMux I__7753 (
            .O(N__37974),
            .I(N__37968));
    InMux I__7752 (
            .O(N__37971),
            .I(N__37965));
    InMux I__7751 (
            .O(N__37968),
            .I(N__37962));
    LocalMux I__7750 (
            .O(N__37965),
            .I(N__37959));
    LocalMux I__7749 (
            .O(N__37962),
            .I(N__37956));
    Odrv4 I__7748 (
            .O(N__37959),
            .I(\current_shift_inst.un38_control_input_5_0 ));
    Odrv12 I__7747 (
            .O(N__37956),
            .I(\current_shift_inst.un38_control_input_5_0 ));
    InMux I__7746 (
            .O(N__37951),
            .I(N__37948));
    LocalMux I__7745 (
            .O(N__37948),
            .I(N__37945));
    Span4Mux_h I__7744 (
            .O(N__37945),
            .I(N__37942));
    Odrv4 I__7743 (
            .O(N__37942),
            .I(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ));
    InMux I__7742 (
            .O(N__37939),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ));
    CascadeMux I__7741 (
            .O(N__37936),
            .I(N__37928));
    CascadeMux I__7740 (
            .O(N__37935),
            .I(N__37923));
    InMux I__7739 (
            .O(N__37934),
            .I(N__37916));
    InMux I__7738 (
            .O(N__37933),
            .I(N__37916));
    InMux I__7737 (
            .O(N__37932),
            .I(N__37916));
    CascadeMux I__7736 (
            .O(N__37931),
            .I(N__37913));
    InMux I__7735 (
            .O(N__37928),
            .I(N__37905));
    InMux I__7734 (
            .O(N__37927),
            .I(N__37900));
    InMux I__7733 (
            .O(N__37926),
            .I(N__37900));
    InMux I__7732 (
            .O(N__37923),
            .I(N__37897));
    LocalMux I__7731 (
            .O(N__37916),
            .I(N__37894));
    InMux I__7730 (
            .O(N__37913),
            .I(N__37881));
    InMux I__7729 (
            .O(N__37912),
            .I(N__37881));
    InMux I__7728 (
            .O(N__37911),
            .I(N__37881));
    InMux I__7727 (
            .O(N__37910),
            .I(N__37881));
    InMux I__7726 (
            .O(N__37909),
            .I(N__37881));
    InMux I__7725 (
            .O(N__37908),
            .I(N__37881));
    LocalMux I__7724 (
            .O(N__37905),
            .I(N__37878));
    LocalMux I__7723 (
            .O(N__37900),
            .I(N__37873));
    LocalMux I__7722 (
            .O(N__37897),
            .I(N__37873));
    Span4Mux_h I__7721 (
            .O(N__37894),
            .I(N__37870));
    LocalMux I__7720 (
            .O(N__37881),
            .I(N__37867));
    Span4Mux_h I__7719 (
            .O(N__37878),
            .I(N__37864));
    Span4Mux_h I__7718 (
            .O(N__37873),
            .I(N__37861));
    Odrv4 I__7717 (
            .O(N__37870),
            .I(\delay_measurement_inst.elapsed_time_tr_31 ));
    Odrv12 I__7716 (
            .O(N__37867),
            .I(\delay_measurement_inst.elapsed_time_tr_31 ));
    Odrv4 I__7715 (
            .O(N__37864),
            .I(\delay_measurement_inst.elapsed_time_tr_31 ));
    Odrv4 I__7714 (
            .O(N__37861),
            .I(\delay_measurement_inst.elapsed_time_tr_31 ));
    CascadeMux I__7713 (
            .O(N__37852),
            .I(N__37849));
    InMux I__7712 (
            .O(N__37849),
            .I(N__37846));
    LocalMux I__7711 (
            .O(N__37846),
            .I(N__37840));
    InMux I__7710 (
            .O(N__37845),
            .I(N__37837));
    InMux I__7709 (
            .O(N__37844),
            .I(N__37832));
    InMux I__7708 (
            .O(N__37843),
            .I(N__37832));
    Span4Mux_h I__7707 (
            .O(N__37840),
            .I(N__37827));
    LocalMux I__7706 (
            .O(N__37837),
            .I(N__37827));
    LocalMux I__7705 (
            .O(N__37832),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    Odrv4 I__7704 (
            .O(N__37827),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    InMux I__7703 (
            .O(N__37822),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ));
    InMux I__7702 (
            .O(N__37819),
            .I(N__37816));
    LocalMux I__7701 (
            .O(N__37816),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    InMux I__7700 (
            .O(N__37813),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ));
    InMux I__7699 (
            .O(N__37810),
            .I(N__37807));
    LocalMux I__7698 (
            .O(N__37807),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    InMux I__7697 (
            .O(N__37804),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ));
    InMux I__7696 (
            .O(N__37801),
            .I(N__37798));
    LocalMux I__7695 (
            .O(N__37798),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    InMux I__7694 (
            .O(N__37795),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__7693 (
            .O(N__37792),
            .I(N__37789));
    InMux I__7692 (
            .O(N__37789),
            .I(N__37786));
    LocalMux I__7691 (
            .O(N__37786),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    InMux I__7690 (
            .O(N__37783),
            .I(bfn_15_14_0_));
    InMux I__7689 (
            .O(N__37780),
            .I(N__37777));
    LocalMux I__7688 (
            .O(N__37777),
            .I(N__37774));
    Odrv12 I__7687 (
            .O(N__37774),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    InMux I__7686 (
            .O(N__37771),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__7685 (
            .O(N__37768),
            .I(N__37765));
    LocalMux I__7684 (
            .O(N__37765),
            .I(N__37762));
    Odrv4 I__7683 (
            .O(N__37762),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    InMux I__7682 (
            .O(N__37759),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ));
    CascadeMux I__7681 (
            .O(N__37756),
            .I(N__37753));
    InMux I__7680 (
            .O(N__37753),
            .I(N__37750));
    LocalMux I__7679 (
            .O(N__37750),
            .I(N__37747));
    Span4Mux_v I__7678 (
            .O(N__37747),
            .I(N__37744));
    Odrv4 I__7677 (
            .O(N__37744),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30 ));
    InMux I__7676 (
            .O(N__37741),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__7675 (
            .O(N__37738),
            .I(N__37733));
    InMux I__7674 (
            .O(N__37737),
            .I(N__37728));
    InMux I__7673 (
            .O(N__37736),
            .I(N__37725));
    LocalMux I__7672 (
            .O(N__37733),
            .I(N__37722));
    InMux I__7671 (
            .O(N__37732),
            .I(N__37717));
    InMux I__7670 (
            .O(N__37731),
            .I(N__37717));
    LocalMux I__7669 (
            .O(N__37728),
            .I(N__37712));
    LocalMux I__7668 (
            .O(N__37725),
            .I(N__37712));
    Span4Mux_v I__7667 (
            .O(N__37722),
            .I(N__37705));
    LocalMux I__7666 (
            .O(N__37717),
            .I(N__37705));
    Span4Mux_v I__7665 (
            .O(N__37712),
            .I(N__37705));
    Odrv4 I__7664 (
            .O(N__37705),
            .I(\delay_measurement_inst.delay_tr_reg3lto14 ));
    InMux I__7663 (
            .O(N__37702),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ));
    CascadeMux I__7662 (
            .O(N__37699),
            .I(N__37696));
    InMux I__7661 (
            .O(N__37696),
            .I(N__37687));
    InMux I__7660 (
            .O(N__37695),
            .I(N__37687));
    CascadeMux I__7659 (
            .O(N__37694),
            .I(N__37683));
    InMux I__7658 (
            .O(N__37693),
            .I(N__37680));
    InMux I__7657 (
            .O(N__37692),
            .I(N__37677));
    LocalMux I__7656 (
            .O(N__37687),
            .I(N__37674));
    InMux I__7655 (
            .O(N__37686),
            .I(N__37669));
    InMux I__7654 (
            .O(N__37683),
            .I(N__37669));
    LocalMux I__7653 (
            .O(N__37680),
            .I(N__37660));
    LocalMux I__7652 (
            .O(N__37677),
            .I(N__37660));
    Span4Mux_v I__7651 (
            .O(N__37674),
            .I(N__37660));
    LocalMux I__7650 (
            .O(N__37669),
            .I(N__37660));
    Span4Mux_v I__7649 (
            .O(N__37660),
            .I(N__37657));
    Odrv4 I__7648 (
            .O(N__37657),
            .I(\delay_measurement_inst.delay_tr_reg3lto15 ));
    InMux I__7647 (
            .O(N__37654),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ));
    InMux I__7646 (
            .O(N__37651),
            .I(N__37648));
    LocalMux I__7645 (
            .O(N__37648),
            .I(N__37643));
    InMux I__7644 (
            .O(N__37647),
            .I(N__37640));
    InMux I__7643 (
            .O(N__37646),
            .I(N__37637));
    Span4Mux_v I__7642 (
            .O(N__37643),
            .I(N__37634));
    LocalMux I__7641 (
            .O(N__37640),
            .I(N__37629));
    LocalMux I__7640 (
            .O(N__37637),
            .I(N__37629));
    Span4Mux_h I__7639 (
            .O(N__37634),
            .I(N__37626));
    Span4Mux_v I__7638 (
            .O(N__37629),
            .I(N__37623));
    Odrv4 I__7637 (
            .O(N__37626),
            .I(\delay_measurement_inst.elapsed_time_tr_16 ));
    Odrv4 I__7636 (
            .O(N__37623),
            .I(\delay_measurement_inst.elapsed_time_tr_16 ));
    InMux I__7635 (
            .O(N__37618),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__7634 (
            .O(N__37615),
            .I(N__37611));
    InMux I__7633 (
            .O(N__37614),
            .I(N__37607));
    InMux I__7632 (
            .O(N__37611),
            .I(N__37604));
    InMux I__7631 (
            .O(N__37610),
            .I(N__37601));
    LocalMux I__7630 (
            .O(N__37607),
            .I(N__37598));
    LocalMux I__7629 (
            .O(N__37604),
            .I(N__37595));
    LocalMux I__7628 (
            .O(N__37601),
            .I(N__37592));
    Span4Mux_v I__7627 (
            .O(N__37598),
            .I(N__37589));
    Span4Mux_h I__7626 (
            .O(N__37595),
            .I(N__37586));
    Span4Mux_h I__7625 (
            .O(N__37592),
            .I(N__37583));
    Odrv4 I__7624 (
            .O(N__37589),
            .I(\delay_measurement_inst.elapsed_time_tr_17 ));
    Odrv4 I__7623 (
            .O(N__37586),
            .I(\delay_measurement_inst.elapsed_time_tr_17 ));
    Odrv4 I__7622 (
            .O(N__37583),
            .I(\delay_measurement_inst.elapsed_time_tr_17 ));
    InMux I__7621 (
            .O(N__37576),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ));
    InMux I__7620 (
            .O(N__37573),
            .I(N__37568));
    InMux I__7619 (
            .O(N__37572),
            .I(N__37565));
    InMux I__7618 (
            .O(N__37571),
            .I(N__37562));
    LocalMux I__7617 (
            .O(N__37568),
            .I(N__37559));
    LocalMux I__7616 (
            .O(N__37565),
            .I(N__37556));
    LocalMux I__7615 (
            .O(N__37562),
            .I(N__37553));
    Span4Mux_v I__7614 (
            .O(N__37559),
            .I(N__37550));
    Span4Mux_h I__7613 (
            .O(N__37556),
            .I(N__37547));
    Span4Mux_h I__7612 (
            .O(N__37553),
            .I(N__37544));
    Odrv4 I__7611 (
            .O(N__37550),
            .I(\delay_measurement_inst.elapsed_time_tr_18 ));
    Odrv4 I__7610 (
            .O(N__37547),
            .I(\delay_measurement_inst.elapsed_time_tr_18 ));
    Odrv4 I__7609 (
            .O(N__37544),
            .I(\delay_measurement_inst.elapsed_time_tr_18 ));
    InMux I__7608 (
            .O(N__37537),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ));
    InMux I__7607 (
            .O(N__37534),
            .I(N__37529));
    InMux I__7606 (
            .O(N__37533),
            .I(N__37526));
    CascadeMux I__7605 (
            .O(N__37532),
            .I(N__37523));
    LocalMux I__7604 (
            .O(N__37529),
            .I(N__37520));
    LocalMux I__7603 (
            .O(N__37526),
            .I(N__37517));
    InMux I__7602 (
            .O(N__37523),
            .I(N__37514));
    Span4Mux_v I__7601 (
            .O(N__37520),
            .I(N__37511));
    Span4Mux_h I__7600 (
            .O(N__37517),
            .I(N__37508));
    LocalMux I__7599 (
            .O(N__37514),
            .I(N__37505));
    Odrv4 I__7598 (
            .O(N__37511),
            .I(\delay_measurement_inst.elapsed_time_tr_19 ));
    Odrv4 I__7597 (
            .O(N__37508),
            .I(\delay_measurement_inst.elapsed_time_tr_19 ));
    Odrv12 I__7596 (
            .O(N__37505),
            .I(\delay_measurement_inst.elapsed_time_tr_19 ));
    InMux I__7595 (
            .O(N__37498),
            .I(bfn_15_13_0_));
    InMux I__7594 (
            .O(N__37495),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ));
    InMux I__7593 (
            .O(N__37492),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__7592 (
            .O(N__37489),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ));
    InMux I__7591 (
            .O(N__37486),
            .I(N__37475));
    InMux I__7590 (
            .O(N__37485),
            .I(N__37475));
    InMux I__7589 (
            .O(N__37484),
            .I(N__37465));
    InMux I__7588 (
            .O(N__37483),
            .I(N__37465));
    InMux I__7587 (
            .O(N__37482),
            .I(N__37465));
    InMux I__7586 (
            .O(N__37481),
            .I(N__37465));
    InMux I__7585 (
            .O(N__37480),
            .I(N__37462));
    LocalMux I__7584 (
            .O(N__37475),
            .I(N__37459));
    InMux I__7583 (
            .O(N__37474),
            .I(N__37456));
    LocalMux I__7582 (
            .O(N__37465),
            .I(N__37451));
    LocalMux I__7581 (
            .O(N__37462),
            .I(N__37451));
    Span4Mux_v I__7580 (
            .O(N__37459),
            .I(N__37446));
    LocalMux I__7579 (
            .O(N__37456),
            .I(N__37446));
    Span4Mux_v I__7578 (
            .O(N__37451),
            .I(N__37443));
    Span4Mux_h I__7577 (
            .O(N__37446),
            .I(N__37440));
    Odrv4 I__7576 (
            .O(N__37443),
            .I(\delay_measurement_inst.delay_tr_reg3lto6 ));
    Odrv4 I__7575 (
            .O(N__37440),
            .I(\delay_measurement_inst.delay_tr_reg3lto6 ));
    InMux I__7574 (
            .O(N__37435),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ));
    InMux I__7573 (
            .O(N__37432),
            .I(N__37428));
    InMux I__7572 (
            .O(N__37431),
            .I(N__37425));
    LocalMux I__7571 (
            .O(N__37428),
            .I(N__37422));
    LocalMux I__7570 (
            .O(N__37425),
            .I(N__37419));
    Span4Mux_v I__7569 (
            .O(N__37422),
            .I(N__37416));
    Span4Mux_v I__7568 (
            .O(N__37419),
            .I(N__37413));
    Odrv4 I__7567 (
            .O(N__37416),
            .I(\delay_measurement_inst.elapsed_time_tr_7 ));
    Odrv4 I__7566 (
            .O(N__37413),
            .I(\delay_measurement_inst.elapsed_time_tr_7 ));
    InMux I__7565 (
            .O(N__37408),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ));
    InMux I__7564 (
            .O(N__37405),
            .I(N__37401));
    InMux I__7563 (
            .O(N__37404),
            .I(N__37398));
    LocalMux I__7562 (
            .O(N__37401),
            .I(N__37395));
    LocalMux I__7561 (
            .O(N__37398),
            .I(N__37392));
    Span4Mux_v I__7560 (
            .O(N__37395),
            .I(N__37389));
    Odrv12 I__7559 (
            .O(N__37392),
            .I(\delay_measurement_inst.elapsed_time_tr_8 ));
    Odrv4 I__7558 (
            .O(N__37389),
            .I(\delay_measurement_inst.elapsed_time_tr_8 ));
    InMux I__7557 (
            .O(N__37384),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__7556 (
            .O(N__37381),
            .I(N__37377));
    InMux I__7555 (
            .O(N__37380),
            .I(N__37372));
    InMux I__7554 (
            .O(N__37377),
            .I(N__37372));
    LocalMux I__7553 (
            .O(N__37372),
            .I(N__37366));
    InMux I__7552 (
            .O(N__37371),
            .I(N__37363));
    InMux I__7551 (
            .O(N__37370),
            .I(N__37360));
    InMux I__7550 (
            .O(N__37369),
            .I(N__37357));
    Span4Mux_h I__7549 (
            .O(N__37366),
            .I(N__37354));
    LocalMux I__7548 (
            .O(N__37363),
            .I(N__37349));
    LocalMux I__7547 (
            .O(N__37360),
            .I(N__37349));
    LocalMux I__7546 (
            .O(N__37357),
            .I(N__37346));
    Span4Mux_h I__7545 (
            .O(N__37354),
            .I(N__37343));
    Span4Mux_h I__7544 (
            .O(N__37349),
            .I(N__37340));
    Span4Mux_h I__7543 (
            .O(N__37346),
            .I(N__37337));
    Odrv4 I__7542 (
            .O(N__37343),
            .I(\delay_measurement_inst.delay_tr_reg3lto9 ));
    Odrv4 I__7541 (
            .O(N__37340),
            .I(\delay_measurement_inst.delay_tr_reg3lto9 ));
    Odrv4 I__7540 (
            .O(N__37337),
            .I(\delay_measurement_inst.delay_tr_reg3lto9 ));
    InMux I__7539 (
            .O(N__37330),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ));
    InMux I__7538 (
            .O(N__37327),
            .I(N__37324));
    LocalMux I__7537 (
            .O(N__37324),
            .I(N__37320));
    InMux I__7536 (
            .O(N__37323),
            .I(N__37317));
    Span4Mux_v I__7535 (
            .O(N__37320),
            .I(N__37312));
    LocalMux I__7534 (
            .O(N__37317),
            .I(N__37312));
    Span4Mux_h I__7533 (
            .O(N__37312),
            .I(N__37309));
    Odrv4 I__7532 (
            .O(N__37309),
            .I(\delay_measurement_inst.elapsed_time_tr_10 ));
    InMux I__7531 (
            .O(N__37306),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ));
    InMux I__7530 (
            .O(N__37303),
            .I(N__37300));
    LocalMux I__7529 (
            .O(N__37300),
            .I(N__37296));
    InMux I__7528 (
            .O(N__37299),
            .I(N__37293));
    Span12Mux_v I__7527 (
            .O(N__37296),
            .I(N__37288));
    LocalMux I__7526 (
            .O(N__37293),
            .I(N__37288));
    Odrv12 I__7525 (
            .O(N__37288),
            .I(\delay_measurement_inst.elapsed_time_tr_11 ));
    InMux I__7524 (
            .O(N__37285),
            .I(bfn_15_12_0_));
    InMux I__7523 (
            .O(N__37282),
            .I(N__37279));
    LocalMux I__7522 (
            .O(N__37279),
            .I(N__37275));
    InMux I__7521 (
            .O(N__37278),
            .I(N__37272));
    Span4Mux_h I__7520 (
            .O(N__37275),
            .I(N__37269));
    LocalMux I__7519 (
            .O(N__37272),
            .I(N__37266));
    Odrv4 I__7518 (
            .O(N__37269),
            .I(\delay_measurement_inst.elapsed_time_tr_12 ));
    Odrv12 I__7517 (
            .O(N__37266),
            .I(\delay_measurement_inst.elapsed_time_tr_12 ));
    InMux I__7516 (
            .O(N__37261),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ));
    InMux I__7515 (
            .O(N__37258),
            .I(N__37254));
    CascadeMux I__7514 (
            .O(N__37257),
            .I(N__37251));
    LocalMux I__7513 (
            .O(N__37254),
            .I(N__37248));
    InMux I__7512 (
            .O(N__37251),
            .I(N__37245));
    Span4Mux_v I__7511 (
            .O(N__37248),
            .I(N__37240));
    LocalMux I__7510 (
            .O(N__37245),
            .I(N__37240));
    Odrv4 I__7509 (
            .O(N__37240),
            .I(\delay_measurement_inst.elapsed_time_tr_13 ));
    InMux I__7508 (
            .O(N__37237),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ));
    InMux I__7507 (
            .O(N__37234),
            .I(N__37229));
    InMux I__7506 (
            .O(N__37233),
            .I(N__37226));
    InMux I__7505 (
            .O(N__37232),
            .I(N__37223));
    LocalMux I__7504 (
            .O(N__37229),
            .I(N__37220));
    LocalMux I__7503 (
            .O(N__37226),
            .I(N__37217));
    LocalMux I__7502 (
            .O(N__37223),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ));
    Odrv4 I__7501 (
            .O(N__37220),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ));
    Odrv4 I__7500 (
            .O(N__37217),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ));
    InMux I__7499 (
            .O(N__37210),
            .I(N__37207));
    LocalMux I__7498 (
            .O(N__37207),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO ));
    InMux I__7497 (
            .O(N__37204),
            .I(N__37201));
    LocalMux I__7496 (
            .O(N__37201),
            .I(N__37196));
    InMux I__7495 (
            .O(N__37200),
            .I(N__37193));
    InMux I__7494 (
            .O(N__37199),
            .I(N__37190));
    Sp12to4 I__7493 (
            .O(N__37196),
            .I(N__37185));
    LocalMux I__7492 (
            .O(N__37193),
            .I(N__37185));
    LocalMux I__7491 (
            .O(N__37190),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ));
    Odrv12 I__7490 (
            .O(N__37185),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ));
    InMux I__7489 (
            .O(N__37180),
            .I(N__37177));
    LocalMux I__7488 (
            .O(N__37177),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO ));
    InMux I__7487 (
            .O(N__37174),
            .I(N__37169));
    InMux I__7486 (
            .O(N__37173),
            .I(N__37166));
    InMux I__7485 (
            .O(N__37172),
            .I(N__37163));
    LocalMux I__7484 (
            .O(N__37169),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ));
    LocalMux I__7483 (
            .O(N__37166),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ));
    LocalMux I__7482 (
            .O(N__37163),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ));
    CascadeMux I__7481 (
            .O(N__37156),
            .I(N__37153));
    InMux I__7480 (
            .O(N__37153),
            .I(N__37150));
    LocalMux I__7479 (
            .O(N__37150),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO ));
    InMux I__7478 (
            .O(N__37147),
            .I(N__37143));
    InMux I__7477 (
            .O(N__37146),
            .I(N__37140));
    LocalMux I__7476 (
            .O(N__37143),
            .I(N__37137));
    LocalMux I__7475 (
            .O(N__37140),
            .I(N__37134));
    Span4Mux_h I__7474 (
            .O(N__37137),
            .I(N__37128));
    Span4Mux_h I__7473 (
            .O(N__37134),
            .I(N__37128));
    InMux I__7472 (
            .O(N__37133),
            .I(N__37125));
    Odrv4 I__7471 (
            .O(N__37128),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_20 ));
    LocalMux I__7470 (
            .O(N__37125),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_20 ));
    CascadeMux I__7469 (
            .O(N__37120),
            .I(N__37117));
    InMux I__7468 (
            .O(N__37117),
            .I(N__37112));
    InMux I__7467 (
            .O(N__37116),
            .I(N__37109));
    InMux I__7466 (
            .O(N__37115),
            .I(N__37106));
    LocalMux I__7465 (
            .O(N__37112),
            .I(N__37103));
    LocalMux I__7464 (
            .O(N__37109),
            .I(N__37100));
    LocalMux I__7463 (
            .O(N__37106),
            .I(N__37095));
    Span4Mux_h I__7462 (
            .O(N__37103),
            .I(N__37090));
    Span4Mux_h I__7461 (
            .O(N__37100),
            .I(N__37090));
    InMux I__7460 (
            .O(N__37099),
            .I(N__37085));
    InMux I__7459 (
            .O(N__37098),
            .I(N__37085));
    Span4Mux_h I__7458 (
            .O(N__37095),
            .I(N__37082));
    Odrv4 I__7457 (
            .O(N__37090),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    LocalMux I__7456 (
            .O(N__37085),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    Odrv4 I__7455 (
            .O(N__37082),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    InMux I__7454 (
            .O(N__37075),
            .I(N__37072));
    LocalMux I__7453 (
            .O(N__37072),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_20 ));
    InMux I__7452 (
            .O(N__37069),
            .I(N__37066));
    LocalMux I__7451 (
            .O(N__37066),
            .I(N__37061));
    InMux I__7450 (
            .O(N__37065),
            .I(N__37058));
    InMux I__7449 (
            .O(N__37064),
            .I(N__37055));
    Sp12to4 I__7448 (
            .O(N__37061),
            .I(N__37050));
    LocalMux I__7447 (
            .O(N__37058),
            .I(N__37050));
    LocalMux I__7446 (
            .O(N__37055),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ));
    Odrv12 I__7445 (
            .O(N__37050),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ));
    InMux I__7444 (
            .O(N__37045),
            .I(N__37042));
    LocalMux I__7443 (
            .O(N__37042),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO ));
    CascadeMux I__7442 (
            .O(N__37039),
            .I(N__37036));
    InMux I__7441 (
            .O(N__37036),
            .I(N__37032));
    InMux I__7440 (
            .O(N__37035),
            .I(N__37028));
    LocalMux I__7439 (
            .O(N__37032),
            .I(N__37025));
    InMux I__7438 (
            .O(N__37031),
            .I(N__37022));
    LocalMux I__7437 (
            .O(N__37028),
            .I(N__37019));
    Span4Mux_v I__7436 (
            .O(N__37025),
            .I(N__37016));
    LocalMux I__7435 (
            .O(N__37022),
            .I(N__37013));
    Span4Mux_v I__7434 (
            .O(N__37019),
            .I(N__37010));
    Span4Mux_h I__7433 (
            .O(N__37016),
            .I(N__37007));
    Span4Mux_v I__7432 (
            .O(N__37013),
            .I(N__37004));
    Span4Mux_h I__7431 (
            .O(N__37010),
            .I(N__37001));
    Odrv4 I__7430 (
            .O(N__37007),
            .I(\delay_measurement_inst.elapsed_time_tr_3 ));
    Odrv4 I__7429 (
            .O(N__37004),
            .I(\delay_measurement_inst.elapsed_time_tr_3 ));
    Odrv4 I__7428 (
            .O(N__37001),
            .I(\delay_measurement_inst.elapsed_time_tr_3 ));
    InMux I__7427 (
            .O(N__36994),
            .I(N__36990));
    InMux I__7426 (
            .O(N__36993),
            .I(N__36987));
    LocalMux I__7425 (
            .O(N__36990),
            .I(N__36982));
    LocalMux I__7424 (
            .O(N__36987),
            .I(N__36982));
    Span4Mux_h I__7423 (
            .O(N__36982),
            .I(N__36979));
    Odrv4 I__7422 (
            .O(N__36979),
            .I(\delay_measurement_inst.elapsed_time_tr_4 ));
    InMux I__7421 (
            .O(N__36976),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ));
    InMux I__7420 (
            .O(N__36973),
            .I(N__36969));
    InMux I__7419 (
            .O(N__36972),
            .I(N__36966));
    LocalMux I__7418 (
            .O(N__36969),
            .I(N__36961));
    LocalMux I__7417 (
            .O(N__36966),
            .I(N__36961));
    Span4Mux_h I__7416 (
            .O(N__36961),
            .I(N__36958));
    Odrv4 I__7415 (
            .O(N__36958),
            .I(\delay_measurement_inst.elapsed_time_tr_5 ));
    InMux I__7414 (
            .O(N__36955),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ));
    InMux I__7413 (
            .O(N__36952),
            .I(N__36947));
    InMux I__7412 (
            .O(N__36951),
            .I(N__36942));
    InMux I__7411 (
            .O(N__36950),
            .I(N__36942));
    LocalMux I__7410 (
            .O(N__36947),
            .I(N__36939));
    LocalMux I__7409 (
            .O(N__36942),
            .I(N__36936));
    Span4Mux_h I__7408 (
            .O(N__36939),
            .I(N__36931));
    Span4Mux_h I__7407 (
            .O(N__36936),
            .I(N__36931));
    Odrv4 I__7406 (
            .O(N__36931),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_19 ));
    CascadeMux I__7405 (
            .O(N__36928),
            .I(N__36924));
    CascadeMux I__7404 (
            .O(N__36927),
            .I(N__36921));
    InMux I__7403 (
            .O(N__36924),
            .I(N__36918));
    InMux I__7402 (
            .O(N__36921),
            .I(N__36915));
    LocalMux I__7401 (
            .O(N__36918),
            .I(N__36912));
    LocalMux I__7400 (
            .O(N__36915),
            .I(N__36908));
    Span4Mux_v I__7399 (
            .O(N__36912),
            .I(N__36903));
    InMux I__7398 (
            .O(N__36911),
            .I(N__36900));
    Span4Mux_v I__7397 (
            .O(N__36908),
            .I(N__36897));
    InMux I__7396 (
            .O(N__36907),
            .I(N__36894));
    InMux I__7395 (
            .O(N__36906),
            .I(N__36891));
    Span4Mux_h I__7394 (
            .O(N__36903),
            .I(N__36886));
    LocalMux I__7393 (
            .O(N__36900),
            .I(N__36886));
    Odrv4 I__7392 (
            .O(N__36897),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    LocalMux I__7391 (
            .O(N__36894),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    LocalMux I__7390 (
            .O(N__36891),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    Odrv4 I__7389 (
            .O(N__36886),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    InMux I__7388 (
            .O(N__36877),
            .I(N__36874));
    LocalMux I__7387 (
            .O(N__36874),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_19 ));
    CascadeMux I__7386 (
            .O(N__36871),
            .I(N__36868));
    InMux I__7385 (
            .O(N__36868),
            .I(N__36865));
    LocalMux I__7384 (
            .O(N__36865),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_15 ));
    InMux I__7383 (
            .O(N__36862),
            .I(N__36858));
    InMux I__7382 (
            .O(N__36861),
            .I(N__36855));
    LocalMux I__7381 (
            .O(N__36858),
            .I(N__36851));
    LocalMux I__7380 (
            .O(N__36855),
            .I(N__36848));
    InMux I__7379 (
            .O(N__36854),
            .I(N__36845));
    Span4Mux_h I__7378 (
            .O(N__36851),
            .I(N__36840));
    Span4Mux_h I__7377 (
            .O(N__36848),
            .I(N__36840));
    LocalMux I__7376 (
            .O(N__36845),
            .I(N__36837));
    Odrv4 I__7375 (
            .O(N__36840),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_15 ));
    Odrv4 I__7374 (
            .O(N__36837),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_15 ));
    CascadeMux I__7373 (
            .O(N__36832),
            .I(N__36828));
    InMux I__7372 (
            .O(N__36831),
            .I(N__36824));
    InMux I__7371 (
            .O(N__36828),
            .I(N__36821));
    InMux I__7370 (
            .O(N__36827),
            .I(N__36816));
    LocalMux I__7369 (
            .O(N__36824),
            .I(N__36813));
    LocalMux I__7368 (
            .O(N__36821),
            .I(N__36810));
    InMux I__7367 (
            .O(N__36820),
            .I(N__36807));
    CascadeMux I__7366 (
            .O(N__36819),
            .I(N__36804));
    LocalMux I__7365 (
            .O(N__36816),
            .I(N__36801));
    Span4Mux_v I__7364 (
            .O(N__36813),
            .I(N__36796));
    Span4Mux_h I__7363 (
            .O(N__36810),
            .I(N__36796));
    LocalMux I__7362 (
            .O(N__36807),
            .I(N__36793));
    InMux I__7361 (
            .O(N__36804),
            .I(N__36790));
    Span4Mux_h I__7360 (
            .O(N__36801),
            .I(N__36787));
    Odrv4 I__7359 (
            .O(N__36796),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    Odrv12 I__7358 (
            .O(N__36793),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    LocalMux I__7357 (
            .O(N__36790),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    Odrv4 I__7356 (
            .O(N__36787),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    InMux I__7355 (
            .O(N__36778),
            .I(N__36775));
    LocalMux I__7354 (
            .O(N__36775),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_16 ));
    InMux I__7353 (
            .O(N__36772),
            .I(N__36768));
    InMux I__7352 (
            .O(N__36771),
            .I(N__36765));
    LocalMux I__7351 (
            .O(N__36768),
            .I(N__36761));
    LocalMux I__7350 (
            .O(N__36765),
            .I(N__36758));
    InMux I__7349 (
            .O(N__36764),
            .I(N__36755));
    Span4Mux_h I__7348 (
            .O(N__36761),
            .I(N__36752));
    Span4Mux_h I__7347 (
            .O(N__36758),
            .I(N__36749));
    LocalMux I__7346 (
            .O(N__36755),
            .I(N__36746));
    Odrv4 I__7345 (
            .O(N__36752),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_16 ));
    Odrv4 I__7344 (
            .O(N__36749),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_16 ));
    Odrv4 I__7343 (
            .O(N__36746),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_16 ));
    InMux I__7342 (
            .O(N__36739),
            .I(N__36735));
    InMux I__7341 (
            .O(N__36738),
            .I(N__36732));
    LocalMux I__7340 (
            .O(N__36735),
            .I(N__36729));
    LocalMux I__7339 (
            .O(N__36732),
            .I(N__36726));
    Span4Mux_h I__7338 (
            .O(N__36729),
            .I(N__36722));
    Span4Mux_h I__7337 (
            .O(N__36726),
            .I(N__36719));
    InMux I__7336 (
            .O(N__36725),
            .I(N__36716));
    Odrv4 I__7335 (
            .O(N__36722),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_23 ));
    Odrv4 I__7334 (
            .O(N__36719),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_23 ));
    LocalMux I__7333 (
            .O(N__36716),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_23 ));
    InMux I__7332 (
            .O(N__36709),
            .I(N__36706));
    LocalMux I__7331 (
            .O(N__36706),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_23 ));
    InMux I__7330 (
            .O(N__36703),
            .I(N__36699));
    InMux I__7329 (
            .O(N__36702),
            .I(N__36696));
    LocalMux I__7328 (
            .O(N__36699),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ));
    LocalMux I__7327 (
            .O(N__36696),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ));
    CascadeMux I__7326 (
            .O(N__36691),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_27_cascade_ ));
    InMux I__7325 (
            .O(N__36688),
            .I(N__36685));
    LocalMux I__7324 (
            .O(N__36685),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO ));
    InMux I__7323 (
            .O(N__36682),
            .I(N__36679));
    LocalMux I__7322 (
            .O(N__36679),
            .I(N__36674));
    InMux I__7321 (
            .O(N__36678),
            .I(N__36671));
    InMux I__7320 (
            .O(N__36677),
            .I(N__36668));
    Span4Mux_h I__7319 (
            .O(N__36674),
            .I(N__36665));
    LocalMux I__7318 (
            .O(N__36671),
            .I(N__36660));
    LocalMux I__7317 (
            .O(N__36668),
            .I(N__36660));
    Odrv4 I__7316 (
            .O(N__36665),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    Odrv4 I__7315 (
            .O(N__36660),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    InMux I__7314 (
            .O(N__36655),
            .I(N__36652));
    LocalMux I__7313 (
            .O(N__36652),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_7 ));
    CascadeMux I__7312 (
            .O(N__36649),
            .I(N__36646));
    InMux I__7311 (
            .O(N__36646),
            .I(N__36643));
    LocalMux I__7310 (
            .O(N__36643),
            .I(N__36639));
    InMux I__7309 (
            .O(N__36642),
            .I(N__36635));
    Span4Mux_h I__7308 (
            .O(N__36639),
            .I(N__36632));
    InMux I__7307 (
            .O(N__36638),
            .I(N__36629));
    LocalMux I__7306 (
            .O(N__36635),
            .I(N__36626));
    Span4Mux_h I__7305 (
            .O(N__36632),
            .I(N__36621));
    LocalMux I__7304 (
            .O(N__36629),
            .I(N__36621));
    Odrv12 I__7303 (
            .O(N__36626),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    Odrv4 I__7302 (
            .O(N__36621),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    InMux I__7301 (
            .O(N__36616),
            .I(N__36613));
    LocalMux I__7300 (
            .O(N__36613),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_9 ));
    InMux I__7299 (
            .O(N__36610),
            .I(N__36606));
    InMux I__7298 (
            .O(N__36609),
            .I(N__36603));
    LocalMux I__7297 (
            .O(N__36606),
            .I(N__36599));
    LocalMux I__7296 (
            .O(N__36603),
            .I(N__36596));
    InMux I__7295 (
            .O(N__36602),
            .I(N__36593));
    Span4Mux_h I__7294 (
            .O(N__36599),
            .I(N__36590));
    Span4Mux_h I__7293 (
            .O(N__36596),
            .I(N__36585));
    LocalMux I__7292 (
            .O(N__36593),
            .I(N__36585));
    Odrv4 I__7291 (
            .O(N__36590),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    Odrv4 I__7290 (
            .O(N__36585),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    InMux I__7289 (
            .O(N__36580),
            .I(N__36577));
    LocalMux I__7288 (
            .O(N__36577),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_10 ));
    CascadeMux I__7287 (
            .O(N__36574),
            .I(N__36571));
    InMux I__7286 (
            .O(N__36571),
            .I(N__36567));
    InMux I__7285 (
            .O(N__36570),
            .I(N__36564));
    LocalMux I__7284 (
            .O(N__36567),
            .I(N__36561));
    LocalMux I__7283 (
            .O(N__36564),
            .I(N__36557));
    Span4Mux_v I__7282 (
            .O(N__36561),
            .I(N__36554));
    InMux I__7281 (
            .O(N__36560),
            .I(N__36551));
    Span4Mux_v I__7280 (
            .O(N__36557),
            .I(N__36546));
    Span4Mux_v I__7279 (
            .O(N__36554),
            .I(N__36546));
    LocalMux I__7278 (
            .O(N__36551),
            .I(N__36543));
    Odrv4 I__7277 (
            .O(N__36546),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    Odrv4 I__7276 (
            .O(N__36543),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    InMux I__7275 (
            .O(N__36538),
            .I(N__36535));
    LocalMux I__7274 (
            .O(N__36535),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_12 ));
    CascadeMux I__7273 (
            .O(N__36532),
            .I(N__36527));
    InMux I__7272 (
            .O(N__36531),
            .I(N__36524));
    InMux I__7271 (
            .O(N__36530),
            .I(N__36521));
    InMux I__7270 (
            .O(N__36527),
            .I(N__36518));
    LocalMux I__7269 (
            .O(N__36524),
            .I(N__36514));
    LocalMux I__7268 (
            .O(N__36521),
            .I(N__36511));
    LocalMux I__7267 (
            .O(N__36518),
            .I(N__36508));
    InMux I__7266 (
            .O(N__36517),
            .I(N__36505));
    Span4Mux_v I__7265 (
            .O(N__36514),
            .I(N__36502));
    Span4Mux_v I__7264 (
            .O(N__36511),
            .I(N__36499));
    Span4Mux_h I__7263 (
            .O(N__36508),
            .I(N__36492));
    LocalMux I__7262 (
            .O(N__36505),
            .I(N__36492));
    Span4Mux_h I__7261 (
            .O(N__36502),
            .I(N__36492));
    Odrv4 I__7260 (
            .O(N__36499),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv4 I__7259 (
            .O(N__36492),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    InMux I__7258 (
            .O(N__36487),
            .I(N__36483));
    InMux I__7257 (
            .O(N__36486),
            .I(N__36480));
    LocalMux I__7256 (
            .O(N__36483),
            .I(N__36476));
    LocalMux I__7255 (
            .O(N__36480),
            .I(N__36473));
    InMux I__7254 (
            .O(N__36479),
            .I(N__36470));
    Span4Mux_h I__7253 (
            .O(N__36476),
            .I(N__36465));
    Span4Mux_v I__7252 (
            .O(N__36473),
            .I(N__36465));
    LocalMux I__7251 (
            .O(N__36470),
            .I(N__36462));
    Odrv4 I__7250 (
            .O(N__36465),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    Odrv4 I__7249 (
            .O(N__36462),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    InMux I__7248 (
            .O(N__36457),
            .I(N__36454));
    LocalMux I__7247 (
            .O(N__36454),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_11 ));
    InMux I__7246 (
            .O(N__36451),
            .I(N__36447));
    InMux I__7245 (
            .O(N__36450),
            .I(N__36444));
    LocalMux I__7244 (
            .O(N__36447),
            .I(N__36441));
    LocalMux I__7243 (
            .O(N__36444),
            .I(N__36438));
    Span4Mux_h I__7242 (
            .O(N__36441),
            .I(N__36434));
    Span4Mux_h I__7241 (
            .O(N__36438),
            .I(N__36431));
    InMux I__7240 (
            .O(N__36437),
            .I(N__36428));
    Odrv4 I__7239 (
            .O(N__36434),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_22 ));
    Odrv4 I__7238 (
            .O(N__36431),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_22 ));
    LocalMux I__7237 (
            .O(N__36428),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_22 ));
    InMux I__7236 (
            .O(N__36421),
            .I(N__36418));
    LocalMux I__7235 (
            .O(N__36418),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_22 ));
    CEMux I__7234 (
            .O(N__36415),
            .I(N__36412));
    LocalMux I__7233 (
            .O(N__36412),
            .I(N__36406));
    CEMux I__7232 (
            .O(N__36411),
            .I(N__36403));
    CEMux I__7231 (
            .O(N__36410),
            .I(N__36400));
    CEMux I__7230 (
            .O(N__36409),
            .I(N__36396));
    Span4Mux_h I__7229 (
            .O(N__36406),
            .I(N__36392));
    LocalMux I__7228 (
            .O(N__36403),
            .I(N__36389));
    LocalMux I__7227 (
            .O(N__36400),
            .I(N__36386));
    CEMux I__7226 (
            .O(N__36399),
            .I(N__36383));
    LocalMux I__7225 (
            .O(N__36396),
            .I(N__36380));
    IoInMux I__7224 (
            .O(N__36395),
            .I(N__36377));
    Sp12to4 I__7223 (
            .O(N__36392),
            .I(N__36374));
    Span4Mux_v I__7222 (
            .O(N__36389),
            .I(N__36371));
    Span4Mux_h I__7221 (
            .O(N__36386),
            .I(N__36366));
    LocalMux I__7220 (
            .O(N__36383),
            .I(N__36366));
    Span4Mux_v I__7219 (
            .O(N__36380),
            .I(N__36363));
    LocalMux I__7218 (
            .O(N__36377),
            .I(N__36360));
    Span12Mux_v I__7217 (
            .O(N__36374),
            .I(N__36357));
    Sp12to4 I__7216 (
            .O(N__36371),
            .I(N__36354));
    Span4Mux_v I__7215 (
            .O(N__36366),
            .I(N__36351));
    Span4Mux_v I__7214 (
            .O(N__36363),
            .I(N__36348));
    Span4Mux_s2_v I__7213 (
            .O(N__36360),
            .I(N__36345));
    Span12Mux_v I__7212 (
            .O(N__36357),
            .I(N__36342));
    Span12Mux_v I__7211 (
            .O(N__36354),
            .I(N__36339));
    Span4Mux_v I__7210 (
            .O(N__36351),
            .I(N__36336));
    Span4Mux_v I__7209 (
            .O(N__36348),
            .I(N__36331));
    Span4Mux_h I__7208 (
            .O(N__36345),
            .I(N__36331));
    Odrv12 I__7207 (
            .O(N__36342),
            .I(red_c_i));
    Odrv12 I__7206 (
            .O(N__36339),
            .I(red_c_i));
    Odrv4 I__7205 (
            .O(N__36336),
            .I(red_c_i));
    Odrv4 I__7204 (
            .O(N__36331),
            .I(red_c_i));
    InMux I__7203 (
            .O(N__36322),
            .I(N__36318));
    InMux I__7202 (
            .O(N__36321),
            .I(N__36315));
    LocalMux I__7201 (
            .O(N__36318),
            .I(N__36312));
    LocalMux I__7200 (
            .O(N__36315),
            .I(N__36308));
    Span4Mux_h I__7199 (
            .O(N__36312),
            .I(N__36305));
    InMux I__7198 (
            .O(N__36311),
            .I(N__36302));
    Span4Mux_h I__7197 (
            .O(N__36308),
            .I(N__36299));
    Span4Mux_v I__7196 (
            .O(N__36305),
            .I(N__36296));
    LocalMux I__7195 (
            .O(N__36302),
            .I(N__36293));
    Odrv4 I__7194 (
            .O(N__36299),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_13 ));
    Odrv4 I__7193 (
            .O(N__36296),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_13 ));
    Odrv4 I__7192 (
            .O(N__36293),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_13 ));
    InMux I__7191 (
            .O(N__36286),
            .I(N__36283));
    LocalMux I__7190 (
            .O(N__36283),
            .I(N__36280));
    Odrv4 I__7189 (
            .O(N__36280),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_13 ));
    InMux I__7188 (
            .O(N__36277),
            .I(N__36273));
    InMux I__7187 (
            .O(N__36276),
            .I(N__36270));
    LocalMux I__7186 (
            .O(N__36273),
            .I(N__36266));
    LocalMux I__7185 (
            .O(N__36270),
            .I(N__36263));
    InMux I__7184 (
            .O(N__36269),
            .I(N__36260));
    Span4Mux_h I__7183 (
            .O(N__36266),
            .I(N__36257));
    Span4Mux_h I__7182 (
            .O(N__36263),
            .I(N__36252));
    LocalMux I__7181 (
            .O(N__36260),
            .I(N__36252));
    Odrv4 I__7180 (
            .O(N__36257),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    Odrv4 I__7179 (
            .O(N__36252),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    InMux I__7178 (
            .O(N__36247),
            .I(N__36244));
    LocalMux I__7177 (
            .O(N__36244),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_6 ));
    InMux I__7176 (
            .O(N__36241),
            .I(N__36237));
    InMux I__7175 (
            .O(N__36240),
            .I(N__36234));
    LocalMux I__7174 (
            .O(N__36237),
            .I(N__36230));
    LocalMux I__7173 (
            .O(N__36234),
            .I(N__36227));
    InMux I__7172 (
            .O(N__36233),
            .I(N__36224));
    Span4Mux_v I__7171 (
            .O(N__36230),
            .I(N__36219));
    Span4Mux_v I__7170 (
            .O(N__36227),
            .I(N__36219));
    LocalMux I__7169 (
            .O(N__36224),
            .I(N__36216));
    Odrv4 I__7168 (
            .O(N__36219),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    Odrv4 I__7167 (
            .O(N__36216),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    InMux I__7166 (
            .O(N__36211),
            .I(N__36208));
    LocalMux I__7165 (
            .O(N__36208),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_5 ));
    InMux I__7164 (
            .O(N__36205),
            .I(N__36201));
    InMux I__7163 (
            .O(N__36204),
            .I(N__36198));
    LocalMux I__7162 (
            .O(N__36201),
            .I(N__36194));
    LocalMux I__7161 (
            .O(N__36198),
            .I(N__36191));
    InMux I__7160 (
            .O(N__36197),
            .I(N__36188));
    Span4Mux_v I__7159 (
            .O(N__36194),
            .I(N__36183));
    Span4Mux_v I__7158 (
            .O(N__36191),
            .I(N__36183));
    LocalMux I__7157 (
            .O(N__36188),
            .I(N__36180));
    Odrv4 I__7156 (
            .O(N__36183),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_4 ));
    Odrv4 I__7155 (
            .O(N__36180),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_4 ));
    InMux I__7154 (
            .O(N__36175),
            .I(N__36172));
    LocalMux I__7153 (
            .O(N__36172),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_4 ));
    InMux I__7152 (
            .O(N__36169),
            .I(N__36165));
    InMux I__7151 (
            .O(N__36168),
            .I(N__36162));
    LocalMux I__7150 (
            .O(N__36165),
            .I(N__36158));
    LocalMux I__7149 (
            .O(N__36162),
            .I(N__36155));
    InMux I__7148 (
            .O(N__36161),
            .I(N__36152));
    Span4Mux_h I__7147 (
            .O(N__36158),
            .I(N__36149));
    Span4Mux_h I__7146 (
            .O(N__36155),
            .I(N__36144));
    LocalMux I__7145 (
            .O(N__36152),
            .I(N__36144));
    Odrv4 I__7144 (
            .O(N__36149),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    Odrv4 I__7143 (
            .O(N__36144),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    InMux I__7142 (
            .O(N__36139),
            .I(N__36136));
    LocalMux I__7141 (
            .O(N__36136),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_8 ));
    InMux I__7140 (
            .O(N__36133),
            .I(N__36127));
    InMux I__7139 (
            .O(N__36132),
            .I(N__36127));
    LocalMux I__7138 (
            .O(N__36127),
            .I(N__36123));
    InMux I__7137 (
            .O(N__36126),
            .I(N__36120));
    Span4Mux_v I__7136 (
            .O(N__36123),
            .I(N__36117));
    LocalMux I__7135 (
            .O(N__36120),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    Odrv4 I__7134 (
            .O(N__36117),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    CascadeMux I__7133 (
            .O(N__36112),
            .I(N__36109));
    InMux I__7132 (
            .O(N__36109),
            .I(N__36106));
    LocalMux I__7131 (
            .O(N__36106),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    InMux I__7130 (
            .O(N__36103),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__7129 (
            .O(N__36100),
            .I(N__36096));
    InMux I__7128 (
            .O(N__36099),
            .I(N__36093));
    InMux I__7127 (
            .O(N__36096),
            .I(N__36090));
    LocalMux I__7126 (
            .O(N__36093),
            .I(N__36084));
    LocalMux I__7125 (
            .O(N__36090),
            .I(N__36084));
    InMux I__7124 (
            .O(N__36089),
            .I(N__36081));
    Span4Mux_v I__7123 (
            .O(N__36084),
            .I(N__36078));
    LocalMux I__7122 (
            .O(N__36081),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    Odrv4 I__7121 (
            .O(N__36078),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    InMux I__7120 (
            .O(N__36073),
            .I(N__36070));
    LocalMux I__7119 (
            .O(N__36070),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    InMux I__7118 (
            .O(N__36067),
            .I(bfn_14_29_0_));
    InMux I__7117 (
            .O(N__36064),
            .I(N__36060));
    CascadeMux I__7116 (
            .O(N__36063),
            .I(N__36057));
    LocalMux I__7115 (
            .O(N__36060),
            .I(N__36054));
    InMux I__7114 (
            .O(N__36057),
            .I(N__36051));
    Span4Mux_s2_v I__7113 (
            .O(N__36054),
            .I(N__36045));
    LocalMux I__7112 (
            .O(N__36051),
            .I(N__36045));
    InMux I__7111 (
            .O(N__36050),
            .I(N__36042));
    Span4Mux_v I__7110 (
            .O(N__36045),
            .I(N__36039));
    LocalMux I__7109 (
            .O(N__36042),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    Odrv4 I__7108 (
            .O(N__36039),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    InMux I__7107 (
            .O(N__36034),
            .I(N__36031));
    LocalMux I__7106 (
            .O(N__36031),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    InMux I__7105 (
            .O(N__36028),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ));
    CascadeMux I__7104 (
            .O(N__36025),
            .I(N__36021));
    InMux I__7103 (
            .O(N__36024),
            .I(N__36017));
    InMux I__7102 (
            .O(N__36021),
            .I(N__36014));
    InMux I__7101 (
            .O(N__36020),
            .I(N__36011));
    LocalMux I__7100 (
            .O(N__36017),
            .I(N__36006));
    LocalMux I__7099 (
            .O(N__36014),
            .I(N__36006));
    LocalMux I__7098 (
            .O(N__36011),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    Odrv12 I__7097 (
            .O(N__36006),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    CascadeMux I__7096 (
            .O(N__36001),
            .I(N__35998));
    InMux I__7095 (
            .O(N__35998),
            .I(N__35995));
    LocalMux I__7094 (
            .O(N__35995),
            .I(N__35991));
    InMux I__7093 (
            .O(N__35994),
            .I(N__35988));
    Span4Mux_s3_v I__7092 (
            .O(N__35991),
            .I(N__35985));
    LocalMux I__7091 (
            .O(N__35988),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    Odrv4 I__7090 (
            .O(N__35985),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    InMux I__7089 (
            .O(N__35980),
            .I(N__35977));
    LocalMux I__7088 (
            .O(N__35977),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    InMux I__7087 (
            .O(N__35974),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ));
    CascadeMux I__7086 (
            .O(N__35971),
            .I(N__35967));
    InMux I__7085 (
            .O(N__35970),
            .I(N__35963));
    InMux I__7084 (
            .O(N__35967),
            .I(N__35960));
    InMux I__7083 (
            .O(N__35966),
            .I(N__35957));
    LocalMux I__7082 (
            .O(N__35963),
            .I(N__35952));
    LocalMux I__7081 (
            .O(N__35960),
            .I(N__35952));
    LocalMux I__7080 (
            .O(N__35957),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    Odrv12 I__7079 (
            .O(N__35952),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    CascadeMux I__7078 (
            .O(N__35947),
            .I(N__35944));
    InMux I__7077 (
            .O(N__35944),
            .I(N__35940));
    InMux I__7076 (
            .O(N__35943),
            .I(N__35937));
    LocalMux I__7075 (
            .O(N__35940),
            .I(N__35934));
    LocalMux I__7074 (
            .O(N__35937),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    Odrv12 I__7073 (
            .O(N__35934),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    CascadeMux I__7072 (
            .O(N__35929),
            .I(N__35926));
    InMux I__7071 (
            .O(N__35926),
            .I(N__35923));
    LocalMux I__7070 (
            .O(N__35923),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    InMux I__7069 (
            .O(N__35920),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__7068 (
            .O(N__35917),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ));
    InMux I__7067 (
            .O(N__35914),
            .I(N__35911));
    LocalMux I__7066 (
            .O(N__35911),
            .I(N__35907));
    InMux I__7065 (
            .O(N__35910),
            .I(N__35904));
    Odrv4 I__7064 (
            .O(N__35907),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    LocalMux I__7063 (
            .O(N__35904),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    InMux I__7062 (
            .O(N__35899),
            .I(N__35896));
    LocalMux I__7061 (
            .O(N__35896),
            .I(N__35893));
    Odrv12 I__7060 (
            .O(N__35893),
            .I(delay_tr_input_c));
    InMux I__7059 (
            .O(N__35890),
            .I(N__35887));
    LocalMux I__7058 (
            .O(N__35887),
            .I(delay_tr_d1));
    InMux I__7057 (
            .O(N__35884),
            .I(N__35878));
    InMux I__7056 (
            .O(N__35883),
            .I(N__35878));
    LocalMux I__7055 (
            .O(N__35878),
            .I(N__35874));
    InMux I__7054 (
            .O(N__35877),
            .I(N__35871));
    Span4Mux_v I__7053 (
            .O(N__35874),
            .I(N__35868));
    LocalMux I__7052 (
            .O(N__35871),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    Odrv4 I__7051 (
            .O(N__35868),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    InMux I__7050 (
            .O(N__35863),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ));
    InMux I__7049 (
            .O(N__35860),
            .I(N__35856));
    CascadeMux I__7048 (
            .O(N__35859),
            .I(N__35853));
    LocalMux I__7047 (
            .O(N__35856),
            .I(N__35850));
    InMux I__7046 (
            .O(N__35853),
            .I(N__35847));
    Span4Mux_s3_v I__7045 (
            .O(N__35850),
            .I(N__35841));
    LocalMux I__7044 (
            .O(N__35847),
            .I(N__35841));
    InMux I__7043 (
            .O(N__35846),
            .I(N__35838));
    Span4Mux_v I__7042 (
            .O(N__35841),
            .I(N__35835));
    LocalMux I__7041 (
            .O(N__35838),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    Odrv4 I__7040 (
            .O(N__35835),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    InMux I__7039 (
            .O(N__35830),
            .I(bfn_14_28_0_));
    InMux I__7038 (
            .O(N__35827),
            .I(N__35823));
    CascadeMux I__7037 (
            .O(N__35826),
            .I(N__35820));
    LocalMux I__7036 (
            .O(N__35823),
            .I(N__35817));
    InMux I__7035 (
            .O(N__35820),
            .I(N__35814));
    Span4Mux_s3_v I__7034 (
            .O(N__35817),
            .I(N__35808));
    LocalMux I__7033 (
            .O(N__35814),
            .I(N__35808));
    InMux I__7032 (
            .O(N__35813),
            .I(N__35805));
    Span4Mux_v I__7031 (
            .O(N__35808),
            .I(N__35802));
    LocalMux I__7030 (
            .O(N__35805),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    Odrv4 I__7029 (
            .O(N__35802),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    CascadeMux I__7028 (
            .O(N__35797),
            .I(N__35793));
    InMux I__7027 (
            .O(N__35796),
            .I(N__35790));
    InMux I__7026 (
            .O(N__35793),
            .I(N__35787));
    LocalMux I__7025 (
            .O(N__35790),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    LocalMux I__7024 (
            .O(N__35787),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    InMux I__7023 (
            .O(N__35782),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ));
    CascadeMux I__7022 (
            .O(N__35779),
            .I(N__35775));
    InMux I__7021 (
            .O(N__35778),
            .I(N__35771));
    InMux I__7020 (
            .O(N__35775),
            .I(N__35768));
    InMux I__7019 (
            .O(N__35774),
            .I(N__35765));
    LocalMux I__7018 (
            .O(N__35771),
            .I(N__35760));
    LocalMux I__7017 (
            .O(N__35768),
            .I(N__35760));
    LocalMux I__7016 (
            .O(N__35765),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    Odrv12 I__7015 (
            .O(N__35760),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    InMux I__7014 (
            .O(N__35755),
            .I(N__35749));
    InMux I__7013 (
            .O(N__35754),
            .I(N__35749));
    LocalMux I__7012 (
            .O(N__35749),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    InMux I__7011 (
            .O(N__35746),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ));
    CascadeMux I__7010 (
            .O(N__35743),
            .I(N__35739));
    InMux I__7009 (
            .O(N__35742),
            .I(N__35735));
    InMux I__7008 (
            .O(N__35739),
            .I(N__35732));
    InMux I__7007 (
            .O(N__35738),
            .I(N__35729));
    LocalMux I__7006 (
            .O(N__35735),
            .I(N__35724));
    LocalMux I__7005 (
            .O(N__35732),
            .I(N__35724));
    LocalMux I__7004 (
            .O(N__35729),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    Odrv12 I__7003 (
            .O(N__35724),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    InMux I__7002 (
            .O(N__35719),
            .I(N__35713));
    InMux I__7001 (
            .O(N__35718),
            .I(N__35713));
    LocalMux I__7000 (
            .O(N__35713),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    InMux I__6999 (
            .O(N__35710),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__6998 (
            .O(N__35707),
            .I(N__35703));
    CascadeMux I__6997 (
            .O(N__35706),
            .I(N__35700));
    InMux I__6996 (
            .O(N__35703),
            .I(N__35695));
    InMux I__6995 (
            .O(N__35700),
            .I(N__35695));
    LocalMux I__6994 (
            .O(N__35695),
            .I(N__35691));
    InMux I__6993 (
            .O(N__35694),
            .I(N__35688));
    Span4Mux_v I__6992 (
            .O(N__35691),
            .I(N__35685));
    LocalMux I__6991 (
            .O(N__35688),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    Odrv4 I__6990 (
            .O(N__35685),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    InMux I__6989 (
            .O(N__35680),
            .I(N__35677));
    LocalMux I__6988 (
            .O(N__35677),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    InMux I__6987 (
            .O(N__35674),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ));
    CascadeMux I__6986 (
            .O(N__35671),
            .I(N__35667));
    CascadeMux I__6985 (
            .O(N__35670),
            .I(N__35664));
    InMux I__6984 (
            .O(N__35667),
            .I(N__35658));
    InMux I__6983 (
            .O(N__35664),
            .I(N__35658));
    InMux I__6982 (
            .O(N__35663),
            .I(N__35655));
    LocalMux I__6981 (
            .O(N__35658),
            .I(N__35652));
    LocalMux I__6980 (
            .O(N__35655),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    Odrv12 I__6979 (
            .O(N__35652),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    InMux I__6978 (
            .O(N__35647),
            .I(N__35644));
    LocalMux I__6977 (
            .O(N__35644),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    InMux I__6976 (
            .O(N__35641),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ));
    InMux I__6975 (
            .O(N__35638),
            .I(N__35632));
    InMux I__6974 (
            .O(N__35637),
            .I(N__35632));
    LocalMux I__6973 (
            .O(N__35632),
            .I(N__35628));
    InMux I__6972 (
            .O(N__35631),
            .I(N__35625));
    Span4Mux_v I__6971 (
            .O(N__35628),
            .I(N__35622));
    LocalMux I__6970 (
            .O(N__35625),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    Odrv4 I__6969 (
            .O(N__35622),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    InMux I__6968 (
            .O(N__35617),
            .I(N__35614));
    LocalMux I__6967 (
            .O(N__35614),
            .I(N__35611));
    Odrv4 I__6966 (
            .O(N__35611),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    InMux I__6965 (
            .O(N__35608),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__6964 (
            .O(N__35605),
            .I(N__35601));
    CascadeMux I__6963 (
            .O(N__35604),
            .I(N__35598));
    InMux I__6962 (
            .O(N__35601),
            .I(N__35593));
    InMux I__6961 (
            .O(N__35598),
            .I(N__35593));
    LocalMux I__6960 (
            .O(N__35593),
            .I(N__35589));
    InMux I__6959 (
            .O(N__35592),
            .I(N__35586));
    Span4Mux_v I__6958 (
            .O(N__35589),
            .I(N__35583));
    LocalMux I__6957 (
            .O(N__35586),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    Odrv4 I__6956 (
            .O(N__35583),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    InMux I__6955 (
            .O(N__35578),
            .I(N__35574));
    InMux I__6954 (
            .O(N__35577),
            .I(N__35571));
    LocalMux I__6953 (
            .O(N__35574),
            .I(N__35568));
    LocalMux I__6952 (
            .O(N__35571),
            .I(N__35565));
    Span4Mux_h I__6951 (
            .O(N__35568),
            .I(N__35561));
    Span4Mux_h I__6950 (
            .O(N__35565),
            .I(N__35558));
    InMux I__6949 (
            .O(N__35564),
            .I(N__35555));
    Odrv4 I__6948 (
            .O(N__35561),
            .I(\delay_measurement_inst.elapsed_time_hc_10 ));
    Odrv4 I__6947 (
            .O(N__35558),
            .I(\delay_measurement_inst.elapsed_time_hc_10 ));
    LocalMux I__6946 (
            .O(N__35555),
            .I(\delay_measurement_inst.elapsed_time_hc_10 ));
    InMux I__6945 (
            .O(N__35548),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__6944 (
            .O(N__35545),
            .I(N__35541));
    InMux I__6943 (
            .O(N__35544),
            .I(N__35537));
    InMux I__6942 (
            .O(N__35541),
            .I(N__35534));
    InMux I__6941 (
            .O(N__35540),
            .I(N__35531));
    LocalMux I__6940 (
            .O(N__35537),
            .I(N__35526));
    LocalMux I__6939 (
            .O(N__35534),
            .I(N__35526));
    LocalMux I__6938 (
            .O(N__35531),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    Odrv12 I__6937 (
            .O(N__35526),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    InMux I__6936 (
            .O(N__35521),
            .I(N__35518));
    LocalMux I__6935 (
            .O(N__35518),
            .I(N__35513));
    InMux I__6934 (
            .O(N__35517),
            .I(N__35510));
    InMux I__6933 (
            .O(N__35516),
            .I(N__35507));
    Span4Mux_v I__6932 (
            .O(N__35513),
            .I(N__35502));
    LocalMux I__6931 (
            .O(N__35510),
            .I(N__35502));
    LocalMux I__6930 (
            .O(N__35507),
            .I(\delay_measurement_inst.elapsed_time_hc_11 ));
    Odrv4 I__6929 (
            .O(N__35502),
            .I(\delay_measurement_inst.elapsed_time_hc_11 ));
    InMux I__6928 (
            .O(N__35497),
            .I(bfn_14_27_0_));
    InMux I__6927 (
            .O(N__35494),
            .I(N__35491));
    LocalMux I__6926 (
            .O(N__35491),
            .I(N__35487));
    InMux I__6925 (
            .O(N__35490),
            .I(N__35484));
    Span4Mux_v I__6924 (
            .O(N__35487),
            .I(N__35478));
    LocalMux I__6923 (
            .O(N__35484),
            .I(N__35478));
    InMux I__6922 (
            .O(N__35483),
            .I(N__35475));
    Span4Mux_v I__6921 (
            .O(N__35478),
            .I(N__35472));
    LocalMux I__6920 (
            .O(N__35475),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    Odrv4 I__6919 (
            .O(N__35472),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    InMux I__6918 (
            .O(N__35467),
            .I(N__35463));
    InMux I__6917 (
            .O(N__35466),
            .I(N__35460));
    LocalMux I__6916 (
            .O(N__35463),
            .I(N__35456));
    LocalMux I__6915 (
            .O(N__35460),
            .I(N__35453));
    InMux I__6914 (
            .O(N__35459),
            .I(N__35450));
    Span4Mux_v I__6913 (
            .O(N__35456),
            .I(N__35445));
    Span4Mux_h I__6912 (
            .O(N__35453),
            .I(N__35445));
    LocalMux I__6911 (
            .O(N__35450),
            .I(\delay_measurement_inst.elapsed_time_hc_12 ));
    Odrv4 I__6910 (
            .O(N__35445),
            .I(\delay_measurement_inst.elapsed_time_hc_12 ));
    InMux I__6909 (
            .O(N__35440),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__6908 (
            .O(N__35437),
            .I(N__35433));
    InMux I__6907 (
            .O(N__35436),
            .I(N__35429));
    InMux I__6906 (
            .O(N__35433),
            .I(N__35426));
    InMux I__6905 (
            .O(N__35432),
            .I(N__35423));
    LocalMux I__6904 (
            .O(N__35429),
            .I(N__35418));
    LocalMux I__6903 (
            .O(N__35426),
            .I(N__35418));
    LocalMux I__6902 (
            .O(N__35423),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    Odrv12 I__6901 (
            .O(N__35418),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    InMux I__6900 (
            .O(N__35413),
            .I(N__35409));
    CascadeMux I__6899 (
            .O(N__35412),
            .I(N__35406));
    LocalMux I__6898 (
            .O(N__35409),
            .I(N__35403));
    InMux I__6897 (
            .O(N__35406),
            .I(N__35399));
    Span4Mux_h I__6896 (
            .O(N__35403),
            .I(N__35396));
    InMux I__6895 (
            .O(N__35402),
            .I(N__35393));
    LocalMux I__6894 (
            .O(N__35399),
            .I(N__35390));
    Odrv4 I__6893 (
            .O(N__35396),
            .I(\delay_measurement_inst.elapsed_time_hc_13 ));
    LocalMux I__6892 (
            .O(N__35393),
            .I(\delay_measurement_inst.elapsed_time_hc_13 ));
    Odrv4 I__6891 (
            .O(N__35390),
            .I(\delay_measurement_inst.elapsed_time_hc_13 ));
    InMux I__6890 (
            .O(N__35383),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ));
    CascadeMux I__6889 (
            .O(N__35380),
            .I(N__35376));
    InMux I__6888 (
            .O(N__35379),
            .I(N__35372));
    InMux I__6887 (
            .O(N__35376),
            .I(N__35369));
    InMux I__6886 (
            .O(N__35375),
            .I(N__35366));
    LocalMux I__6885 (
            .O(N__35372),
            .I(N__35361));
    LocalMux I__6884 (
            .O(N__35369),
            .I(N__35361));
    LocalMux I__6883 (
            .O(N__35366),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    Odrv12 I__6882 (
            .O(N__35361),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    InMux I__6881 (
            .O(N__35356),
            .I(N__35353));
    LocalMux I__6880 (
            .O(N__35353),
            .I(N__35350));
    Span4Mux_h I__6879 (
            .O(N__35350),
            .I(N__35344));
    InMux I__6878 (
            .O(N__35349),
            .I(N__35339));
    InMux I__6877 (
            .O(N__35348),
            .I(N__35339));
    InMux I__6876 (
            .O(N__35347),
            .I(N__35336));
    Odrv4 I__6875 (
            .O(N__35344),
            .I(\delay_measurement_inst.delay_hc_reg3lto14 ));
    LocalMux I__6874 (
            .O(N__35339),
            .I(\delay_measurement_inst.delay_hc_reg3lto14 ));
    LocalMux I__6873 (
            .O(N__35336),
            .I(\delay_measurement_inst.delay_hc_reg3lto14 ));
    InMux I__6872 (
            .O(N__35329),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ));
    CascadeMux I__6871 (
            .O(N__35326),
            .I(N__35322));
    CascadeMux I__6870 (
            .O(N__35325),
            .I(N__35319));
    InMux I__6869 (
            .O(N__35322),
            .I(N__35314));
    InMux I__6868 (
            .O(N__35319),
            .I(N__35314));
    LocalMux I__6867 (
            .O(N__35314),
            .I(N__35310));
    InMux I__6866 (
            .O(N__35313),
            .I(N__35307));
    Span4Mux_v I__6865 (
            .O(N__35310),
            .I(N__35304));
    LocalMux I__6864 (
            .O(N__35307),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    Odrv4 I__6863 (
            .O(N__35304),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    InMux I__6862 (
            .O(N__35299),
            .I(N__35295));
    CascadeMux I__6861 (
            .O(N__35298),
            .I(N__35290));
    LocalMux I__6860 (
            .O(N__35295),
            .I(N__35287));
    InMux I__6859 (
            .O(N__35294),
            .I(N__35284));
    InMux I__6858 (
            .O(N__35293),
            .I(N__35279));
    InMux I__6857 (
            .O(N__35290),
            .I(N__35279));
    Odrv4 I__6856 (
            .O(N__35287),
            .I(\delay_measurement_inst.delay_hc_reg3lto15 ));
    LocalMux I__6855 (
            .O(N__35284),
            .I(\delay_measurement_inst.delay_hc_reg3lto15 ));
    LocalMux I__6854 (
            .O(N__35279),
            .I(\delay_measurement_inst.delay_hc_reg3lto15 ));
    InMux I__6853 (
            .O(N__35272),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ));
    CascadeMux I__6852 (
            .O(N__35269),
            .I(N__35265));
    CascadeMux I__6851 (
            .O(N__35268),
            .I(N__35262));
    InMux I__6850 (
            .O(N__35265),
            .I(N__35256));
    InMux I__6849 (
            .O(N__35262),
            .I(N__35256));
    InMux I__6848 (
            .O(N__35261),
            .I(N__35253));
    LocalMux I__6847 (
            .O(N__35256),
            .I(N__35250));
    LocalMux I__6846 (
            .O(N__35253),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    Odrv12 I__6845 (
            .O(N__35250),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    InMux I__6844 (
            .O(N__35245),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ));
    InMux I__6843 (
            .O(N__35242),
            .I(N__35236));
    InMux I__6842 (
            .O(N__35241),
            .I(N__35236));
    LocalMux I__6841 (
            .O(N__35236),
            .I(N__35232));
    InMux I__6840 (
            .O(N__35235),
            .I(N__35229));
    Span4Mux_v I__6839 (
            .O(N__35232),
            .I(N__35226));
    LocalMux I__6838 (
            .O(N__35229),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    Odrv4 I__6837 (
            .O(N__35226),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    InMux I__6836 (
            .O(N__35221),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ));
    CascadeMux I__6835 (
            .O(N__35218),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6_cascade_ ));
    InMux I__6834 (
            .O(N__35215),
            .I(N__35212));
    LocalMux I__6833 (
            .O(N__35212),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_10 ));
    InMux I__6832 (
            .O(N__35209),
            .I(N__35206));
    LocalMux I__6831 (
            .O(N__35206),
            .I(N__35203));
    Span4Mux_h I__6830 (
            .O(N__35203),
            .I(N__35198));
    InMux I__6829 (
            .O(N__35202),
            .I(N__35195));
    InMux I__6828 (
            .O(N__35201),
            .I(N__35192));
    Odrv4 I__6827 (
            .O(N__35198),
            .I(\delay_measurement_inst.elapsed_time_hc_3 ));
    LocalMux I__6826 (
            .O(N__35195),
            .I(\delay_measurement_inst.elapsed_time_hc_3 ));
    LocalMux I__6825 (
            .O(N__35192),
            .I(\delay_measurement_inst.elapsed_time_hc_3 ));
    InMux I__6824 (
            .O(N__35185),
            .I(N__35180));
    InMux I__6823 (
            .O(N__35184),
            .I(N__35175));
    InMux I__6822 (
            .O(N__35183),
            .I(N__35175));
    LocalMux I__6821 (
            .O(N__35180),
            .I(\delay_measurement_inst.elapsed_time_hc_4 ));
    LocalMux I__6820 (
            .O(N__35175),
            .I(\delay_measurement_inst.elapsed_time_hc_4 ));
    InMux I__6819 (
            .O(N__35170),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ));
    CascadeMux I__6818 (
            .O(N__35167),
            .I(N__35163));
    InMux I__6817 (
            .O(N__35166),
            .I(N__35159));
    InMux I__6816 (
            .O(N__35163),
            .I(N__35156));
    InMux I__6815 (
            .O(N__35162),
            .I(N__35153));
    LocalMux I__6814 (
            .O(N__35159),
            .I(N__35148));
    LocalMux I__6813 (
            .O(N__35156),
            .I(N__35148));
    LocalMux I__6812 (
            .O(N__35153),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    Odrv12 I__6811 (
            .O(N__35148),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    InMux I__6810 (
            .O(N__35143),
            .I(N__35140));
    LocalMux I__6809 (
            .O(N__35140),
            .I(N__35137));
    Span4Mux_h I__6808 (
            .O(N__35137),
            .I(N__35132));
    InMux I__6807 (
            .O(N__35136),
            .I(N__35127));
    InMux I__6806 (
            .O(N__35135),
            .I(N__35127));
    Odrv4 I__6805 (
            .O(N__35132),
            .I(\delay_measurement_inst.elapsed_time_hc_5 ));
    LocalMux I__6804 (
            .O(N__35127),
            .I(\delay_measurement_inst.elapsed_time_hc_5 ));
    InMux I__6803 (
            .O(N__35122),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__6802 (
            .O(N__35119),
            .I(N__35115));
    InMux I__6801 (
            .O(N__35118),
            .I(N__35111));
    InMux I__6800 (
            .O(N__35115),
            .I(N__35108));
    InMux I__6799 (
            .O(N__35114),
            .I(N__35105));
    LocalMux I__6798 (
            .O(N__35111),
            .I(N__35100));
    LocalMux I__6797 (
            .O(N__35108),
            .I(N__35100));
    LocalMux I__6796 (
            .O(N__35105),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    Odrv12 I__6795 (
            .O(N__35100),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    InMux I__6794 (
            .O(N__35095),
            .I(N__35092));
    LocalMux I__6793 (
            .O(N__35092),
            .I(N__35086));
    InMux I__6792 (
            .O(N__35091),
            .I(N__35079));
    InMux I__6791 (
            .O(N__35090),
            .I(N__35079));
    InMux I__6790 (
            .O(N__35089),
            .I(N__35079));
    Odrv4 I__6789 (
            .O(N__35086),
            .I(\delay_measurement_inst.delay_hc_reg3lto6 ));
    LocalMux I__6788 (
            .O(N__35079),
            .I(\delay_measurement_inst.delay_hc_reg3lto6 ));
    InMux I__6787 (
            .O(N__35074),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ));
    CascadeMux I__6786 (
            .O(N__35071),
            .I(N__35067));
    CascadeMux I__6785 (
            .O(N__35070),
            .I(N__35064));
    InMux I__6784 (
            .O(N__35067),
            .I(N__35059));
    InMux I__6783 (
            .O(N__35064),
            .I(N__35059));
    LocalMux I__6782 (
            .O(N__35059),
            .I(N__35055));
    InMux I__6781 (
            .O(N__35058),
            .I(N__35052));
    Span4Mux_v I__6780 (
            .O(N__35055),
            .I(N__35049));
    LocalMux I__6779 (
            .O(N__35052),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    Odrv4 I__6778 (
            .O(N__35049),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    InMux I__6777 (
            .O(N__35044),
            .I(N__35041));
    LocalMux I__6776 (
            .O(N__35041),
            .I(N__35035));
    InMux I__6775 (
            .O(N__35040),
            .I(N__35032));
    InMux I__6774 (
            .O(N__35039),
            .I(N__35029));
    InMux I__6773 (
            .O(N__35038),
            .I(N__35026));
    Odrv4 I__6772 (
            .O(N__35035),
            .I(\delay_measurement_inst.elapsed_time_hc_7 ));
    LocalMux I__6771 (
            .O(N__35032),
            .I(\delay_measurement_inst.elapsed_time_hc_7 ));
    LocalMux I__6770 (
            .O(N__35029),
            .I(\delay_measurement_inst.elapsed_time_hc_7 ));
    LocalMux I__6769 (
            .O(N__35026),
            .I(\delay_measurement_inst.elapsed_time_hc_7 ));
    InMux I__6768 (
            .O(N__35017),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__6767 (
            .O(N__35014),
            .I(N__35010));
    InMux I__6766 (
            .O(N__35013),
            .I(N__35007));
    InMux I__6765 (
            .O(N__35010),
            .I(N__35004));
    LocalMux I__6764 (
            .O(N__35007),
            .I(N__34998));
    LocalMux I__6763 (
            .O(N__35004),
            .I(N__34998));
    InMux I__6762 (
            .O(N__35003),
            .I(N__34995));
    Span4Mux_v I__6761 (
            .O(N__34998),
            .I(N__34992));
    LocalMux I__6760 (
            .O(N__34995),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    Odrv4 I__6759 (
            .O(N__34992),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    CascadeMux I__6758 (
            .O(N__34987),
            .I(N__34983));
    CascadeMux I__6757 (
            .O(N__34986),
            .I(N__34979));
    InMux I__6756 (
            .O(N__34983),
            .I(N__34976));
    CascadeMux I__6755 (
            .O(N__34982),
            .I(N__34973));
    InMux I__6754 (
            .O(N__34979),
            .I(N__34969));
    LocalMux I__6753 (
            .O(N__34976),
            .I(N__34966));
    InMux I__6752 (
            .O(N__34973),
            .I(N__34963));
    InMux I__6751 (
            .O(N__34972),
            .I(N__34960));
    LocalMux I__6750 (
            .O(N__34969),
            .I(N__34957));
    Odrv4 I__6749 (
            .O(N__34966),
            .I(\delay_measurement_inst.elapsed_time_hc_8 ));
    LocalMux I__6748 (
            .O(N__34963),
            .I(\delay_measurement_inst.elapsed_time_hc_8 ));
    LocalMux I__6747 (
            .O(N__34960),
            .I(\delay_measurement_inst.elapsed_time_hc_8 ));
    Odrv4 I__6746 (
            .O(N__34957),
            .I(\delay_measurement_inst.elapsed_time_hc_8 ));
    InMux I__6745 (
            .O(N__34948),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ));
    InMux I__6744 (
            .O(N__34945),
            .I(N__34939));
    InMux I__6743 (
            .O(N__34944),
            .I(N__34939));
    LocalMux I__6742 (
            .O(N__34939),
            .I(N__34935));
    InMux I__6741 (
            .O(N__34938),
            .I(N__34932));
    Span4Mux_v I__6740 (
            .O(N__34935),
            .I(N__34929));
    LocalMux I__6739 (
            .O(N__34932),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    Odrv4 I__6738 (
            .O(N__34929),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    InMux I__6737 (
            .O(N__34924),
            .I(N__34921));
    LocalMux I__6736 (
            .O(N__34921),
            .I(N__34917));
    CascadeMux I__6735 (
            .O(N__34920),
            .I(N__34913));
    Span4Mux_h I__6734 (
            .O(N__34917),
            .I(N__34909));
    InMux I__6733 (
            .O(N__34916),
            .I(N__34906));
    InMux I__6732 (
            .O(N__34913),
            .I(N__34901));
    InMux I__6731 (
            .O(N__34912),
            .I(N__34901));
    Odrv4 I__6730 (
            .O(N__34909),
            .I(\delay_measurement_inst.delay_hc_reg3lto9 ));
    LocalMux I__6729 (
            .O(N__34906),
            .I(\delay_measurement_inst.delay_hc_reg3lto9 ));
    LocalMux I__6728 (
            .O(N__34901),
            .I(\delay_measurement_inst.delay_hc_reg3lto9 ));
    InMux I__6727 (
            .O(N__34894),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ));
    InMux I__6726 (
            .O(N__34891),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ));
    InMux I__6725 (
            .O(N__34888),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ));
    InMux I__6724 (
            .O(N__34885),
            .I(bfn_14_24_0_));
    InMux I__6723 (
            .O(N__34882),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ));
    InMux I__6722 (
            .O(N__34879),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ));
    InMux I__6721 (
            .O(N__34876),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ));
    InMux I__6720 (
            .O(N__34873),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ));
    InMux I__6719 (
            .O(N__34870),
            .I(N__34840));
    InMux I__6718 (
            .O(N__34869),
            .I(N__34840));
    InMux I__6717 (
            .O(N__34868),
            .I(N__34840));
    InMux I__6716 (
            .O(N__34867),
            .I(N__34840));
    InMux I__6715 (
            .O(N__34866),
            .I(N__34831));
    InMux I__6714 (
            .O(N__34865),
            .I(N__34831));
    InMux I__6713 (
            .O(N__34864),
            .I(N__34831));
    InMux I__6712 (
            .O(N__34863),
            .I(N__34831));
    InMux I__6711 (
            .O(N__34862),
            .I(N__34826));
    InMux I__6710 (
            .O(N__34861),
            .I(N__34826));
    InMux I__6709 (
            .O(N__34860),
            .I(N__34809));
    InMux I__6708 (
            .O(N__34859),
            .I(N__34809));
    InMux I__6707 (
            .O(N__34858),
            .I(N__34809));
    InMux I__6706 (
            .O(N__34857),
            .I(N__34809));
    InMux I__6705 (
            .O(N__34856),
            .I(N__34800));
    InMux I__6704 (
            .O(N__34855),
            .I(N__34800));
    InMux I__6703 (
            .O(N__34854),
            .I(N__34800));
    InMux I__6702 (
            .O(N__34853),
            .I(N__34800));
    InMux I__6701 (
            .O(N__34852),
            .I(N__34791));
    InMux I__6700 (
            .O(N__34851),
            .I(N__34791));
    InMux I__6699 (
            .O(N__34850),
            .I(N__34791));
    InMux I__6698 (
            .O(N__34849),
            .I(N__34791));
    LocalMux I__6697 (
            .O(N__34840),
            .I(N__34784));
    LocalMux I__6696 (
            .O(N__34831),
            .I(N__34784));
    LocalMux I__6695 (
            .O(N__34826),
            .I(N__34784));
    InMux I__6694 (
            .O(N__34825),
            .I(N__34775));
    InMux I__6693 (
            .O(N__34824),
            .I(N__34775));
    InMux I__6692 (
            .O(N__34823),
            .I(N__34775));
    InMux I__6691 (
            .O(N__34822),
            .I(N__34775));
    InMux I__6690 (
            .O(N__34821),
            .I(N__34766));
    InMux I__6689 (
            .O(N__34820),
            .I(N__34766));
    InMux I__6688 (
            .O(N__34819),
            .I(N__34766));
    InMux I__6687 (
            .O(N__34818),
            .I(N__34766));
    LocalMux I__6686 (
            .O(N__34809),
            .I(N__34759));
    LocalMux I__6685 (
            .O(N__34800),
            .I(N__34759));
    LocalMux I__6684 (
            .O(N__34791),
            .I(N__34759));
    Span4Mux_v I__6683 (
            .O(N__34784),
            .I(N__34756));
    LocalMux I__6682 (
            .O(N__34775),
            .I(N__34747));
    LocalMux I__6681 (
            .O(N__34766),
            .I(N__34747));
    Span4Mux_v I__6680 (
            .O(N__34759),
            .I(N__34747));
    Span4Mux_h I__6679 (
            .O(N__34756),
            .I(N__34747));
    Odrv4 I__6678 (
            .O(N__34747),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    InMux I__6677 (
            .O(N__34744),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ));
    CEMux I__6676 (
            .O(N__34741),
            .I(N__34736));
    CEMux I__6675 (
            .O(N__34740),
            .I(N__34733));
    CEMux I__6674 (
            .O(N__34739),
            .I(N__34730));
    LocalMux I__6673 (
            .O(N__34736),
            .I(N__34727));
    LocalMux I__6672 (
            .O(N__34733),
            .I(N__34721));
    LocalMux I__6671 (
            .O(N__34730),
            .I(N__34721));
    Span4Mux_v I__6670 (
            .O(N__34727),
            .I(N__34718));
    CEMux I__6669 (
            .O(N__34726),
            .I(N__34715));
    Span4Mux_v I__6668 (
            .O(N__34721),
            .I(N__34712));
    Span4Mux_h I__6667 (
            .O(N__34718),
            .I(N__34707));
    LocalMux I__6666 (
            .O(N__34715),
            .I(N__34707));
    Span4Mux_h I__6665 (
            .O(N__34712),
            .I(N__34702));
    Span4Mux_h I__6664 (
            .O(N__34707),
            .I(N__34702));
    Span4Mux_v I__6663 (
            .O(N__34702),
            .I(N__34699));
    Span4Mux_v I__6662 (
            .O(N__34699),
            .I(N__34696));
    Odrv4 I__6661 (
            .O(N__34696),
            .I(\delay_measurement_inst.delay_hc_timer.N_303_i ));
    InMux I__6660 (
            .O(N__34693),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ));
    InMux I__6659 (
            .O(N__34690),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ));
    InMux I__6658 (
            .O(N__34687),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ));
    InMux I__6657 (
            .O(N__34684),
            .I(bfn_14_23_0_));
    InMux I__6656 (
            .O(N__34681),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ));
    InMux I__6655 (
            .O(N__34678),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ));
    InMux I__6654 (
            .O(N__34675),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ));
    InMux I__6653 (
            .O(N__34672),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ));
    InMux I__6652 (
            .O(N__34669),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ));
    InMux I__6651 (
            .O(N__34666),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ));
    InMux I__6650 (
            .O(N__34663),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ));
    InMux I__6649 (
            .O(N__34660),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ));
    InMux I__6648 (
            .O(N__34657),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ));
    InMux I__6647 (
            .O(N__34654),
            .I(bfn_14_22_0_));
    InMux I__6646 (
            .O(N__34651),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ));
    InMux I__6645 (
            .O(N__34648),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ));
    InMux I__6644 (
            .O(N__34645),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ));
    InMux I__6643 (
            .O(N__34642),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ));
    InMux I__6642 (
            .O(N__34639),
            .I(N__34636));
    LocalMux I__6641 (
            .O(N__34636),
            .I(\current_shift_inst.un38_control_input_0_s0_25 ));
    InMux I__6640 (
            .O(N__34633),
            .I(N__34630));
    LocalMux I__6639 (
            .O(N__34630),
            .I(N__34627));
    Odrv4 I__6638 (
            .O(N__34627),
            .I(\current_shift_inst.control_input_1_axb_19 ));
    InMux I__6637 (
            .O(N__34624),
            .I(N__34621));
    LocalMux I__6636 (
            .O(N__34621),
            .I(\current_shift_inst.un38_control_input_0_s0_30 ));
    InMux I__6635 (
            .O(N__34618),
            .I(N__34615));
    LocalMux I__6634 (
            .O(N__34615),
            .I(\current_shift_inst.control_input_1_axb_24 ));
    InMux I__6633 (
            .O(N__34612),
            .I(N__34609));
    LocalMux I__6632 (
            .O(N__34609),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ));
    InMux I__6631 (
            .O(N__34606),
            .I(N__34603));
    LocalMux I__6630 (
            .O(N__34603),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ));
    InMux I__6629 (
            .O(N__34600),
            .I(N__34597));
    LocalMux I__6628 (
            .O(N__34597),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ));
    InMux I__6627 (
            .O(N__34594),
            .I(bfn_14_21_0_));
    InMux I__6626 (
            .O(N__34591),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ));
    InMux I__6625 (
            .O(N__34588),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ));
    InMux I__6624 (
            .O(N__34585),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ));
    InMux I__6623 (
            .O(N__34582),
            .I(N__34579));
    LocalMux I__6622 (
            .O(N__34579),
            .I(N__34576));
    Odrv4 I__6621 (
            .O(N__34576),
            .I(\current_shift_inst.un38_control_input_0_s0_22 ));
    InMux I__6620 (
            .O(N__34573),
            .I(N__34570));
    LocalMux I__6619 (
            .O(N__34570),
            .I(\current_shift_inst.control_input_1_axb_16 ));
    InMux I__6618 (
            .O(N__34567),
            .I(N__34564));
    LocalMux I__6617 (
            .O(N__34564),
            .I(N__34561));
    Span4Mux_h I__6616 (
            .O(N__34561),
            .I(N__34558));
    Odrv4 I__6615 (
            .O(N__34558),
            .I(\current_shift_inst.un38_control_input_0_s0_29 ));
    InMux I__6614 (
            .O(N__34555),
            .I(N__34552));
    LocalMux I__6613 (
            .O(N__34552),
            .I(\current_shift_inst.control_input_1_axb_23 ));
    InMux I__6612 (
            .O(N__34549),
            .I(N__34546));
    LocalMux I__6611 (
            .O(N__34546),
            .I(N__34543));
    Odrv4 I__6610 (
            .O(N__34543),
            .I(\current_shift_inst.un38_control_input_0_s0_7 ));
    InMux I__6609 (
            .O(N__34540),
            .I(N__34537));
    LocalMux I__6608 (
            .O(N__34537),
            .I(N__34534));
    Odrv12 I__6607 (
            .O(N__34534),
            .I(\current_shift_inst.control_input_1_axb_1 ));
    InMux I__6606 (
            .O(N__34531),
            .I(N__34528));
    LocalMux I__6605 (
            .O(N__34528),
            .I(N__34525));
    Odrv4 I__6604 (
            .O(N__34525),
            .I(\current_shift_inst.un38_control_input_0_s0_27 ));
    InMux I__6603 (
            .O(N__34522),
            .I(N__34519));
    LocalMux I__6602 (
            .O(N__34519),
            .I(N__34516));
    Odrv4 I__6601 (
            .O(N__34516),
            .I(\current_shift_inst.control_input_1_axb_21 ));
    InMux I__6600 (
            .O(N__34513),
            .I(N__34510));
    LocalMux I__6599 (
            .O(N__34510),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13 ));
    CascadeMux I__6598 (
            .O(N__34507),
            .I(N__34504));
    InMux I__6597 (
            .O(N__34504),
            .I(N__34501));
    LocalMux I__6596 (
            .O(N__34501),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI25021_0_19 ));
    InMux I__6595 (
            .O(N__34498),
            .I(N__34495));
    LocalMux I__6594 (
            .O(N__34495),
            .I(\current_shift_inst.un38_control_input_0_s0_24 ));
    InMux I__6593 (
            .O(N__34492),
            .I(N__34489));
    LocalMux I__6592 (
            .O(N__34489),
            .I(N__34486));
    Odrv4 I__6591 (
            .O(N__34486),
            .I(\current_shift_inst.control_input_1_axb_18 ));
    InMux I__6590 (
            .O(N__34483),
            .I(N__34480));
    LocalMux I__6589 (
            .O(N__34480),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ));
    InMux I__6588 (
            .O(N__34477),
            .I(N__34474));
    LocalMux I__6587 (
            .O(N__34474),
            .I(\current_shift_inst.un38_control_input_0_s0_26 ));
    InMux I__6586 (
            .O(N__34471),
            .I(N__34468));
    LocalMux I__6585 (
            .O(N__34468),
            .I(N__34465));
    Odrv4 I__6584 (
            .O(N__34465),
            .I(\current_shift_inst.control_input_1_axb_20 ));
    InMux I__6583 (
            .O(N__34462),
            .I(N__34459));
    LocalMux I__6582 (
            .O(N__34459),
            .I(N__34456));
    Span4Mux_v I__6581 (
            .O(N__34456),
            .I(N__34453));
    Span4Mux_h I__6580 (
            .O(N__34453),
            .I(N__34450));
    Odrv4 I__6579 (
            .O(N__34450),
            .I(\current_shift_inst.control_inputZ0Z_21 ));
    InMux I__6578 (
            .O(N__34447),
            .I(\current_shift_inst.control_input_1_cry_20 ));
    InMux I__6577 (
            .O(N__34444),
            .I(N__34441));
    LocalMux I__6576 (
            .O(N__34441),
            .I(N__34438));
    Span4Mux_h I__6575 (
            .O(N__34438),
            .I(N__34435));
    Odrv4 I__6574 (
            .O(N__34435),
            .I(\current_shift_inst.control_inputZ0Z_22 ));
    InMux I__6573 (
            .O(N__34432),
            .I(\current_shift_inst.control_input_1_cry_21 ));
    InMux I__6572 (
            .O(N__34429),
            .I(N__34426));
    LocalMux I__6571 (
            .O(N__34426),
            .I(N__34423));
    Odrv12 I__6570 (
            .O(N__34423),
            .I(\current_shift_inst.control_inputZ0Z_23 ));
    InMux I__6569 (
            .O(N__34420),
            .I(\current_shift_inst.control_input_1_cry_22 ));
    InMux I__6568 (
            .O(N__34417),
            .I(N__34414));
    LocalMux I__6567 (
            .O(N__34414),
            .I(N__34411));
    Span4Mux_v I__6566 (
            .O(N__34411),
            .I(N__34408));
    Odrv4 I__6565 (
            .O(N__34408),
            .I(\current_shift_inst.control_inputZ0Z_24 ));
    InMux I__6564 (
            .O(N__34405),
            .I(bfn_14_18_0_));
    InMux I__6563 (
            .O(N__34402),
            .I(N__34399));
    LocalMux I__6562 (
            .O(N__34399),
            .I(N__34396));
    Span4Mux_h I__6561 (
            .O(N__34396),
            .I(N__34393));
    Odrv4 I__6560 (
            .O(N__34393),
            .I(\current_shift_inst.control_input_1_axb_25 ));
    InMux I__6559 (
            .O(N__34390),
            .I(\current_shift_inst.control_input_1_cry_24 ));
    InMux I__6558 (
            .O(N__34387),
            .I(N__34381));
    InMux I__6557 (
            .O(N__34386),
            .I(N__34381));
    LocalMux I__6556 (
            .O(N__34381),
            .I(N__34378));
    Span4Mux_v I__6555 (
            .O(N__34378),
            .I(N__34375));
    Odrv4 I__6554 (
            .O(N__34375),
            .I(\current_shift_inst.control_inputZ0Z_25 ));
    InMux I__6553 (
            .O(N__34372),
            .I(N__34369));
    LocalMux I__6552 (
            .O(N__34369),
            .I(N__34366));
    Odrv4 I__6551 (
            .O(N__34366),
            .I(\current_shift_inst.un38_control_input_0_s0_28 ));
    InMux I__6550 (
            .O(N__34363),
            .I(N__34360));
    LocalMux I__6549 (
            .O(N__34360),
            .I(\current_shift_inst.control_input_1_axb_22 ));
    CascadeMux I__6548 (
            .O(N__34357),
            .I(N__34353));
    InMux I__6547 (
            .O(N__34356),
            .I(N__34350));
    InMux I__6546 (
            .O(N__34353),
            .I(N__34347));
    LocalMux I__6545 (
            .O(N__34350),
            .I(N__34342));
    LocalMux I__6544 (
            .O(N__34347),
            .I(N__34342));
    Odrv4 I__6543 (
            .O(N__34342),
            .I(\current_shift_inst.N_1355_i ));
    InMux I__6542 (
            .O(N__34339),
            .I(N__34336));
    LocalMux I__6541 (
            .O(N__34336),
            .I(\current_shift_inst.un38_control_input_0_s0_6 ));
    InMux I__6540 (
            .O(N__34333),
            .I(N__34330));
    LocalMux I__6539 (
            .O(N__34330),
            .I(N__34327));
    Odrv4 I__6538 (
            .O(N__34327),
            .I(\current_shift_inst.control_input_1_axb_0 ));
    InMux I__6537 (
            .O(N__34324),
            .I(N__34321));
    LocalMux I__6536 (
            .O(N__34321),
            .I(N__34318));
    Odrv4 I__6535 (
            .O(N__34318),
            .I(\current_shift_inst.control_input_1_axb_13 ));
    InMux I__6534 (
            .O(N__34315),
            .I(N__34312));
    LocalMux I__6533 (
            .O(N__34312),
            .I(N__34309));
    Odrv12 I__6532 (
            .O(N__34309),
            .I(\current_shift_inst.control_inputZ0Z_13 ));
    InMux I__6531 (
            .O(N__34306),
            .I(\current_shift_inst.control_input_1_cry_12 ));
    InMux I__6530 (
            .O(N__34303),
            .I(N__34300));
    LocalMux I__6529 (
            .O(N__34300),
            .I(\current_shift_inst.control_input_1_axb_14 ));
    InMux I__6528 (
            .O(N__34297),
            .I(N__34294));
    LocalMux I__6527 (
            .O(N__34294),
            .I(N__34291));
    Odrv12 I__6526 (
            .O(N__34291),
            .I(\current_shift_inst.control_inputZ0Z_14 ));
    InMux I__6525 (
            .O(N__34288),
            .I(\current_shift_inst.control_input_1_cry_13 ));
    InMux I__6524 (
            .O(N__34285),
            .I(N__34282));
    LocalMux I__6523 (
            .O(N__34282),
            .I(\current_shift_inst.control_input_1_axb_15 ));
    InMux I__6522 (
            .O(N__34279),
            .I(N__34276));
    LocalMux I__6521 (
            .O(N__34276),
            .I(N__34273));
    Odrv12 I__6520 (
            .O(N__34273),
            .I(\current_shift_inst.control_inputZ0Z_15 ));
    InMux I__6519 (
            .O(N__34270),
            .I(\current_shift_inst.control_input_1_cry_14 ));
    InMux I__6518 (
            .O(N__34267),
            .I(N__34264));
    LocalMux I__6517 (
            .O(N__34264),
            .I(N__34261));
    Odrv12 I__6516 (
            .O(N__34261),
            .I(\current_shift_inst.control_inputZ0Z_16 ));
    InMux I__6515 (
            .O(N__34258),
            .I(bfn_14_17_0_));
    InMux I__6514 (
            .O(N__34255),
            .I(N__34252));
    LocalMux I__6513 (
            .O(N__34252),
            .I(\current_shift_inst.control_input_1_axb_17 ));
    InMux I__6512 (
            .O(N__34249),
            .I(N__34246));
    LocalMux I__6511 (
            .O(N__34246),
            .I(N__34243));
    Span12Mux_v I__6510 (
            .O(N__34243),
            .I(N__34240));
    Odrv12 I__6509 (
            .O(N__34240),
            .I(\current_shift_inst.control_inputZ0Z_17 ));
    InMux I__6508 (
            .O(N__34237),
            .I(\current_shift_inst.control_input_1_cry_16 ));
    InMux I__6507 (
            .O(N__34234),
            .I(N__34231));
    LocalMux I__6506 (
            .O(N__34231),
            .I(N__34228));
    Odrv12 I__6505 (
            .O(N__34228),
            .I(\current_shift_inst.control_inputZ0Z_18 ));
    InMux I__6504 (
            .O(N__34225),
            .I(\current_shift_inst.control_input_1_cry_17 ));
    InMux I__6503 (
            .O(N__34222),
            .I(N__34219));
    LocalMux I__6502 (
            .O(N__34219),
            .I(N__34216));
    Odrv12 I__6501 (
            .O(N__34216),
            .I(\current_shift_inst.control_inputZ0Z_19 ));
    InMux I__6500 (
            .O(N__34213),
            .I(\current_shift_inst.control_input_1_cry_18 ));
    InMux I__6499 (
            .O(N__34210),
            .I(N__34207));
    LocalMux I__6498 (
            .O(N__34207),
            .I(N__34204));
    Odrv12 I__6497 (
            .O(N__34204),
            .I(\current_shift_inst.control_inputZ0Z_20 ));
    InMux I__6496 (
            .O(N__34201),
            .I(\current_shift_inst.control_input_1_cry_19 ));
    InMux I__6495 (
            .O(N__34198),
            .I(N__34195));
    LocalMux I__6494 (
            .O(N__34195),
            .I(N__34192));
    Odrv4 I__6493 (
            .O(N__34192),
            .I(\current_shift_inst.control_inputZ0Z_5 ));
    InMux I__6492 (
            .O(N__34189),
            .I(\current_shift_inst.control_input_1_cry_4 ));
    InMux I__6491 (
            .O(N__34186),
            .I(N__34183));
    LocalMux I__6490 (
            .O(N__34183),
            .I(\current_shift_inst.control_input_1_axb_6 ));
    InMux I__6489 (
            .O(N__34180),
            .I(N__34177));
    LocalMux I__6488 (
            .O(N__34177),
            .I(\current_shift_inst.control_inputZ0Z_6 ));
    InMux I__6487 (
            .O(N__34174),
            .I(\current_shift_inst.control_input_1_cry_5 ));
    InMux I__6486 (
            .O(N__34171),
            .I(N__34168));
    LocalMux I__6485 (
            .O(N__34168),
            .I(N__34165));
    Odrv12 I__6484 (
            .O(N__34165),
            .I(\current_shift_inst.control_inputZ0Z_7 ));
    InMux I__6483 (
            .O(N__34162),
            .I(\current_shift_inst.control_input_1_cry_6 ));
    InMux I__6482 (
            .O(N__34159),
            .I(N__34156));
    LocalMux I__6481 (
            .O(N__34156),
            .I(\current_shift_inst.control_input_1_axb_8 ));
    InMux I__6480 (
            .O(N__34153),
            .I(N__34150));
    LocalMux I__6479 (
            .O(N__34150),
            .I(N__34147));
    Odrv12 I__6478 (
            .O(N__34147),
            .I(\current_shift_inst.control_inputZ0Z_8 ));
    InMux I__6477 (
            .O(N__34144),
            .I(bfn_14_16_0_));
    InMux I__6476 (
            .O(N__34141),
            .I(N__34138));
    LocalMux I__6475 (
            .O(N__34138),
            .I(\current_shift_inst.control_input_1_axb_9 ));
    InMux I__6474 (
            .O(N__34135),
            .I(N__34132));
    LocalMux I__6473 (
            .O(N__34132),
            .I(N__34129));
    Span4Mux_h I__6472 (
            .O(N__34129),
            .I(N__34126));
    Span4Mux_v I__6471 (
            .O(N__34126),
            .I(N__34123));
    Odrv4 I__6470 (
            .O(N__34123),
            .I(\current_shift_inst.control_inputZ0Z_9 ));
    InMux I__6469 (
            .O(N__34120),
            .I(\current_shift_inst.control_input_1_cry_8 ));
    InMux I__6468 (
            .O(N__34117),
            .I(N__34114));
    LocalMux I__6467 (
            .O(N__34114),
            .I(N__34111));
    Odrv4 I__6466 (
            .O(N__34111),
            .I(\current_shift_inst.control_input_1_axb_10 ));
    InMux I__6465 (
            .O(N__34108),
            .I(N__34105));
    LocalMux I__6464 (
            .O(N__34105),
            .I(N__34102));
    Odrv12 I__6463 (
            .O(N__34102),
            .I(\current_shift_inst.control_inputZ0Z_10 ));
    InMux I__6462 (
            .O(N__34099),
            .I(\current_shift_inst.control_input_1_cry_9 ));
    InMux I__6461 (
            .O(N__34096),
            .I(N__34093));
    LocalMux I__6460 (
            .O(N__34093),
            .I(\current_shift_inst.control_input_1_axb_11 ));
    InMux I__6459 (
            .O(N__34090),
            .I(N__34087));
    LocalMux I__6458 (
            .O(N__34087),
            .I(N__34084));
    Odrv12 I__6457 (
            .O(N__34084),
            .I(\current_shift_inst.control_inputZ0Z_11 ));
    InMux I__6456 (
            .O(N__34081),
            .I(\current_shift_inst.control_input_1_cry_10 ));
    InMux I__6455 (
            .O(N__34078),
            .I(N__34075));
    LocalMux I__6454 (
            .O(N__34075),
            .I(\current_shift_inst.control_input_1_axb_12 ));
    InMux I__6453 (
            .O(N__34072),
            .I(N__34069));
    LocalMux I__6452 (
            .O(N__34069),
            .I(N__34066));
    Odrv4 I__6451 (
            .O(N__34066),
            .I(\current_shift_inst.control_inputZ0Z_12 ));
    InMux I__6450 (
            .O(N__34063),
            .I(\current_shift_inst.control_input_1_cry_11 ));
    InMux I__6449 (
            .O(N__34060),
            .I(N__34057));
    LocalMux I__6448 (
            .O(N__34057),
            .I(N__34054));
    Span4Mux_h I__6447 (
            .O(N__34054),
            .I(N__34051));
    Odrv4 I__6446 (
            .O(N__34051),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15 ));
    InMux I__6445 (
            .O(N__34048),
            .I(N__34035));
    InMux I__6444 (
            .O(N__34047),
            .I(N__34035));
    InMux I__6443 (
            .O(N__34046),
            .I(N__34035));
    InMux I__6442 (
            .O(N__34045),
            .I(N__34030));
    InMux I__6441 (
            .O(N__34044),
            .I(N__34030));
    CascadeMux I__6440 (
            .O(N__34043),
            .I(N__34027));
    InMux I__6439 (
            .O(N__34042),
            .I(N__34022));
    LocalMux I__6438 (
            .O(N__34035),
            .I(N__34016));
    LocalMux I__6437 (
            .O(N__34030),
            .I(N__34016));
    InMux I__6436 (
            .O(N__34027),
            .I(N__34013));
    InMux I__6435 (
            .O(N__34026),
            .I(N__34010));
    InMux I__6434 (
            .O(N__34025),
            .I(N__34007));
    LocalMux I__6433 (
            .O(N__34022),
            .I(N__34004));
    InMux I__6432 (
            .O(N__34021),
            .I(N__34001));
    Span4Mux_h I__6431 (
            .O(N__34016),
            .I(N__33996));
    LocalMux I__6430 (
            .O(N__34013),
            .I(N__33996));
    LocalMux I__6429 (
            .O(N__34010),
            .I(measured_delay_tr_15));
    LocalMux I__6428 (
            .O(N__34007),
            .I(measured_delay_tr_15));
    Odrv4 I__6427 (
            .O(N__34004),
            .I(measured_delay_tr_15));
    LocalMux I__6426 (
            .O(N__34001),
            .I(measured_delay_tr_15));
    Odrv4 I__6425 (
            .O(N__33996),
            .I(measured_delay_tr_15));
    InMux I__6424 (
            .O(N__33985),
            .I(N__33980));
    InMux I__6423 (
            .O(N__33984),
            .I(N__33975));
    InMux I__6422 (
            .O(N__33983),
            .I(N__33975));
    LocalMux I__6421 (
            .O(N__33980),
            .I(N__33972));
    LocalMux I__6420 (
            .O(N__33975),
            .I(N__33969));
    Span4Mux_h I__6419 (
            .O(N__33972),
            .I(N__33963));
    Span4Mux_h I__6418 (
            .O(N__33969),
            .I(N__33960));
    InMux I__6417 (
            .O(N__33968),
            .I(N__33957));
    InMux I__6416 (
            .O(N__33967),
            .I(N__33952));
    InMux I__6415 (
            .O(N__33966),
            .I(N__33952));
    Odrv4 I__6414 (
            .O(N__33963),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15 ));
    Odrv4 I__6413 (
            .O(N__33960),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15 ));
    LocalMux I__6412 (
            .O(N__33957),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15 ));
    LocalMux I__6411 (
            .O(N__33952),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15 ));
    CascadeMux I__6410 (
            .O(N__33943),
            .I(N__33940));
    InMux I__6409 (
            .O(N__33940),
            .I(N__33937));
    LocalMux I__6408 (
            .O(N__33937),
            .I(N__33934));
    Span4Mux_h I__6407 (
            .O(N__33934),
            .I(N__33931));
    Odrv4 I__6406 (
            .O(N__33931),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ));
    CEMux I__6405 (
            .O(N__33928),
            .I(N__33922));
    CEMux I__6404 (
            .O(N__33927),
            .I(N__33918));
    CEMux I__6403 (
            .O(N__33926),
            .I(N__33914));
    CEMux I__6402 (
            .O(N__33925),
            .I(N__33911));
    LocalMux I__6401 (
            .O(N__33922),
            .I(N__33908));
    CEMux I__6400 (
            .O(N__33921),
            .I(N__33905));
    LocalMux I__6399 (
            .O(N__33918),
            .I(N__33902));
    CEMux I__6398 (
            .O(N__33917),
            .I(N__33899));
    LocalMux I__6397 (
            .O(N__33914),
            .I(N__33896));
    LocalMux I__6396 (
            .O(N__33911),
            .I(N__33893));
    Span4Mux_v I__6395 (
            .O(N__33908),
            .I(N__33890));
    LocalMux I__6394 (
            .O(N__33905),
            .I(N__33887));
    Span4Mux_h I__6393 (
            .O(N__33902),
            .I(N__33884));
    LocalMux I__6392 (
            .O(N__33899),
            .I(N__33879));
    Span4Mux_h I__6391 (
            .O(N__33896),
            .I(N__33879));
    Span4Mux_h I__6390 (
            .O(N__33893),
            .I(N__33876));
    Span4Mux_h I__6389 (
            .O(N__33890),
            .I(N__33871));
    Span4Mux_h I__6388 (
            .O(N__33887),
            .I(N__33871));
    Odrv4 I__6387 (
            .O(N__33884),
            .I(\phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv4 I__6386 (
            .O(N__33879),
            .I(\phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv4 I__6385 (
            .O(N__33876),
            .I(\phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv4 I__6384 (
            .O(N__33871),
            .I(\phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa ));
    InMux I__6383 (
            .O(N__33862),
            .I(N__33859));
    LocalMux I__6382 (
            .O(N__33859),
            .I(N__33856));
    Span4Mux_h I__6381 (
            .O(N__33856),
            .I(N__33853));
    Odrv4 I__6380 (
            .O(N__33853),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ));
    InMux I__6379 (
            .O(N__33850),
            .I(N__33847));
    LocalMux I__6378 (
            .O(N__33847),
            .I(N__33844));
    Span4Mux_h I__6377 (
            .O(N__33844),
            .I(N__33841));
    Odrv4 I__6376 (
            .O(N__33841),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23 ));
    InMux I__6375 (
            .O(N__33838),
            .I(N__33835));
    LocalMux I__6374 (
            .O(N__33835),
            .I(N__33831));
    InMux I__6373 (
            .O(N__33834),
            .I(N__33828));
    Span4Mux_v I__6372 (
            .O(N__33831),
            .I(N__33823));
    LocalMux I__6371 (
            .O(N__33828),
            .I(N__33823));
    Span4Mux_v I__6370 (
            .O(N__33823),
            .I(N__33820));
    Odrv4 I__6369 (
            .O(N__33820),
            .I(\current_shift_inst.control_inputZ0Z_0 ));
    InMux I__6368 (
            .O(N__33817),
            .I(N__33814));
    LocalMux I__6367 (
            .O(N__33814),
            .I(N__33811));
    Odrv4 I__6366 (
            .O(N__33811),
            .I(\current_shift_inst.control_inputZ0Z_1 ));
    InMux I__6365 (
            .O(N__33808),
            .I(\current_shift_inst.control_input_1_cry_0 ));
    InMux I__6364 (
            .O(N__33805),
            .I(N__33802));
    LocalMux I__6363 (
            .O(N__33802),
            .I(\current_shift_inst.control_input_1_axb_2 ));
    InMux I__6362 (
            .O(N__33799),
            .I(N__33796));
    LocalMux I__6361 (
            .O(N__33796),
            .I(\current_shift_inst.control_inputZ0Z_2 ));
    InMux I__6360 (
            .O(N__33793),
            .I(\current_shift_inst.control_input_1_cry_1 ));
    InMux I__6359 (
            .O(N__33790),
            .I(N__33787));
    LocalMux I__6358 (
            .O(N__33787),
            .I(\current_shift_inst.control_input_1_axb_3 ));
    InMux I__6357 (
            .O(N__33784),
            .I(N__33781));
    LocalMux I__6356 (
            .O(N__33781),
            .I(N__33778));
    Odrv4 I__6355 (
            .O(N__33778),
            .I(\current_shift_inst.control_inputZ0Z_3 ));
    InMux I__6354 (
            .O(N__33775),
            .I(\current_shift_inst.control_input_1_cry_2 ));
    InMux I__6353 (
            .O(N__33772),
            .I(N__33769));
    LocalMux I__6352 (
            .O(N__33769),
            .I(\current_shift_inst.control_input_1_axb_4 ));
    InMux I__6351 (
            .O(N__33766),
            .I(N__33763));
    LocalMux I__6350 (
            .O(N__33763),
            .I(N__33760));
    Span4Mux_v I__6349 (
            .O(N__33760),
            .I(N__33757));
    Span4Mux_h I__6348 (
            .O(N__33757),
            .I(N__33754));
    Odrv4 I__6347 (
            .O(N__33754),
            .I(\current_shift_inst.control_inputZ0Z_4 ));
    InMux I__6346 (
            .O(N__33751),
            .I(\current_shift_inst.control_input_1_cry_3 ));
    InMux I__6345 (
            .O(N__33748),
            .I(N__33745));
    LocalMux I__6344 (
            .O(N__33745),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ));
    InMux I__6343 (
            .O(N__33742),
            .I(N__33739));
    LocalMux I__6342 (
            .O(N__33739),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ));
    CascadeMux I__6341 (
            .O(N__33736),
            .I(N__33733));
    InMux I__6340 (
            .O(N__33733),
            .I(N__33730));
    LocalMux I__6339 (
            .O(N__33730),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18 ));
    CascadeMux I__6338 (
            .O(N__33727),
            .I(N__33724));
    InMux I__6337 (
            .O(N__33724),
            .I(N__33721));
    LocalMux I__6336 (
            .O(N__33721),
            .I(N__33718));
    Odrv4 I__6335 (
            .O(N__33718),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ));
    InMux I__6334 (
            .O(N__33715),
            .I(N__33712));
    LocalMux I__6333 (
            .O(N__33712),
            .I(N__33709));
    Odrv4 I__6332 (
            .O(N__33709),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14 ));
    InMux I__6331 (
            .O(N__33706),
            .I(N__33703));
    LocalMux I__6330 (
            .O(N__33703),
            .I(N__33700));
    Odrv4 I__6329 (
            .O(N__33700),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ));
    InMux I__6328 (
            .O(N__33697),
            .I(N__33694));
    LocalMux I__6327 (
            .O(N__33694),
            .I(N__33691));
    Odrv4 I__6326 (
            .O(N__33691),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ));
    InMux I__6325 (
            .O(N__33688),
            .I(N__33685));
    LocalMux I__6324 (
            .O(N__33685),
            .I(N__33682));
    Span4Mux_h I__6323 (
            .O(N__33682),
            .I(N__33679));
    Odrv4 I__6322 (
            .O(N__33679),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19 ));
    InMux I__6321 (
            .O(N__33676),
            .I(N__33673));
    LocalMux I__6320 (
            .O(N__33673),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19 ));
    InMux I__6319 (
            .O(N__33670),
            .I(N__33667));
    LocalMux I__6318 (
            .O(N__33667),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ));
    InMux I__6317 (
            .O(N__33664),
            .I(N__33661));
    LocalMux I__6316 (
            .O(N__33661),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ));
    InMux I__6315 (
            .O(N__33658),
            .I(N__33655));
    LocalMux I__6314 (
            .O(N__33655),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16 ));
    InMux I__6313 (
            .O(N__33652),
            .I(N__33649));
    LocalMux I__6312 (
            .O(N__33649),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ));
    InMux I__6311 (
            .O(N__33646),
            .I(N__33643));
    LocalMux I__6310 (
            .O(N__33643),
            .I(N__33640));
    Odrv12 I__6309 (
            .O(N__33640),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ));
    InMux I__6308 (
            .O(N__33637),
            .I(N__33634));
    LocalMux I__6307 (
            .O(N__33634),
            .I(N__33631));
    Odrv4 I__6306 (
            .O(N__33631),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ));
    InMux I__6305 (
            .O(N__33628),
            .I(N__33625));
    LocalMux I__6304 (
            .O(N__33625),
            .I(N__33622));
    Odrv4 I__6303 (
            .O(N__33622),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ));
    InMux I__6302 (
            .O(N__33619),
            .I(N__33616));
    LocalMux I__6301 (
            .O(N__33616),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20 ));
    InMux I__6300 (
            .O(N__33613),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27 ));
    InMux I__6299 (
            .O(N__33610),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28 ));
    InMux I__6298 (
            .O(N__33607),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29 ));
    InMux I__6297 (
            .O(N__33604),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_31 ));
    InMux I__6296 (
            .O(N__33601),
            .I(N__33598));
    LocalMux I__6295 (
            .O(N__33598),
            .I(N__33595));
    Odrv4 I__6294 (
            .O(N__33595),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ));
    InMux I__6293 (
            .O(N__33592),
            .I(N__33589));
    LocalMux I__6292 (
            .O(N__33589),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ));
    InMux I__6291 (
            .O(N__33586),
            .I(N__33583));
    LocalMux I__6290 (
            .O(N__33583),
            .I(N__33580));
    Odrv4 I__6289 (
            .O(N__33580),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ));
    InMux I__6288 (
            .O(N__33577),
            .I(N__33574));
    LocalMux I__6287 (
            .O(N__33574),
            .I(N__33571));
    Odrv4 I__6286 (
            .O(N__33571),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ));
    InMux I__6285 (
            .O(N__33568),
            .I(N__33565));
    LocalMux I__6284 (
            .O(N__33565),
            .I(N__33562));
    Odrv4 I__6283 (
            .O(N__33562),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ));
    InMux I__6282 (
            .O(N__33559),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18 ));
    InMux I__6281 (
            .O(N__33556),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19 ));
    InMux I__6280 (
            .O(N__33553),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20 ));
    InMux I__6279 (
            .O(N__33550),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21 ));
    InMux I__6278 (
            .O(N__33547),
            .I(N__33544));
    LocalMux I__6277 (
            .O(N__33544),
            .I(N__33541));
    Span4Mux_h I__6276 (
            .O(N__33541),
            .I(N__33538));
    Odrv4 I__6275 (
            .O(N__33538),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ));
    InMux I__6274 (
            .O(N__33535),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22 ));
    InMux I__6273 (
            .O(N__33532),
            .I(bfn_14_10_0_));
    InMux I__6272 (
            .O(N__33529),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24 ));
    InMux I__6271 (
            .O(N__33526),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25 ));
    InMux I__6270 (
            .O(N__33523),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26 ));
    InMux I__6269 (
            .O(N__33520),
            .I(N__33517));
    LocalMux I__6268 (
            .O(N__33517),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_10 ));
    InMux I__6267 (
            .O(N__33514),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_9 ));
    InMux I__6266 (
            .O(N__33511),
            .I(N__33508));
    LocalMux I__6265 (
            .O(N__33508),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_11 ));
    InMux I__6264 (
            .O(N__33505),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_10 ));
    InMux I__6263 (
            .O(N__33502),
            .I(N__33499));
    LocalMux I__6262 (
            .O(N__33499),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_12 ));
    InMux I__6261 (
            .O(N__33496),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11 ));
    InMux I__6260 (
            .O(N__33493),
            .I(N__33490));
    LocalMux I__6259 (
            .O(N__33490),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_13 ));
    InMux I__6258 (
            .O(N__33487),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12 ));
    InMux I__6257 (
            .O(N__33484),
            .I(N__33481));
    LocalMux I__6256 (
            .O(N__33481),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ));
    InMux I__6255 (
            .O(N__33478),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13 ));
    InMux I__6254 (
            .O(N__33475),
            .I(N__33472));
    LocalMux I__6253 (
            .O(N__33472),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_15 ));
    InMux I__6252 (
            .O(N__33469),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14 ));
    InMux I__6251 (
            .O(N__33466),
            .I(N__33463));
    LocalMux I__6250 (
            .O(N__33463),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ));
    InMux I__6249 (
            .O(N__33460),
            .I(bfn_14_9_0_));
    InMux I__6248 (
            .O(N__33457),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16 ));
    InMux I__6247 (
            .O(N__33454),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17 ));
    InMux I__6246 (
            .O(N__33451),
            .I(N__33447));
    InMux I__6245 (
            .O(N__33450),
            .I(N__33444));
    LocalMux I__6244 (
            .O(N__33447),
            .I(N__33441));
    LocalMux I__6243 (
            .O(N__33444),
            .I(N__33438));
    Span4Mux_v I__6242 (
            .O(N__33441),
            .I(N__33435));
    Span4Mux_h I__6241 (
            .O(N__33438),
            .I(N__33432));
    Odrv4 I__6240 (
            .O(N__33435),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_2 ));
    Odrv4 I__6239 (
            .O(N__33432),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_2 ));
    InMux I__6238 (
            .O(N__33427),
            .I(N__33424));
    LocalMux I__6237 (
            .O(N__33424),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_2 ));
    InMux I__6236 (
            .O(N__33421),
            .I(N__33417));
    InMux I__6235 (
            .O(N__33420),
            .I(N__33414));
    LocalMux I__6234 (
            .O(N__33417),
            .I(N__33411));
    LocalMux I__6233 (
            .O(N__33414),
            .I(N__33408));
    Odrv4 I__6232 (
            .O(N__33411),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_3 ));
    Odrv4 I__6231 (
            .O(N__33408),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_3 ));
    InMux I__6230 (
            .O(N__33403),
            .I(N__33400));
    LocalMux I__6229 (
            .O(N__33400),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_3 ));
    InMux I__6228 (
            .O(N__33397),
            .I(N__33394));
    LocalMux I__6227 (
            .O(N__33394),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_4 ));
    InMux I__6226 (
            .O(N__33391),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_3 ));
    CascadeMux I__6225 (
            .O(N__33388),
            .I(N__33385));
    InMux I__6224 (
            .O(N__33385),
            .I(N__33382));
    LocalMux I__6223 (
            .O(N__33382),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_5 ));
    InMux I__6222 (
            .O(N__33379),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_4 ));
    InMux I__6221 (
            .O(N__33376),
            .I(N__33373));
    LocalMux I__6220 (
            .O(N__33373),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_6 ));
    InMux I__6219 (
            .O(N__33370),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_5 ));
    InMux I__6218 (
            .O(N__33367),
            .I(N__33364));
    LocalMux I__6217 (
            .O(N__33364),
            .I(N__33361));
    Odrv4 I__6216 (
            .O(N__33361),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_7 ));
    InMux I__6215 (
            .O(N__33358),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_6 ));
    InMux I__6214 (
            .O(N__33355),
            .I(N__33352));
    LocalMux I__6213 (
            .O(N__33352),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_8 ));
    InMux I__6212 (
            .O(N__33349),
            .I(bfn_14_8_0_));
    InMux I__6211 (
            .O(N__33346),
            .I(N__33343));
    LocalMux I__6210 (
            .O(N__33343),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_9 ));
    InMux I__6209 (
            .O(N__33340),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_8 ));
    InMux I__6208 (
            .O(N__33337),
            .I(N__33334));
    LocalMux I__6207 (
            .O(N__33334),
            .I(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1 ));
    CascadeMux I__6206 (
            .O(N__33331),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8_cascade_ ));
    InMux I__6205 (
            .O(N__33328),
            .I(N__33325));
    LocalMux I__6204 (
            .O(N__33325),
            .I(N__33322));
    Odrv4 I__6203 (
            .O(N__33322),
            .I(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_3 ));
    InMux I__6202 (
            .O(N__33319),
            .I(N__33313));
    InMux I__6201 (
            .O(N__33318),
            .I(N__33310));
    InMux I__6200 (
            .O(N__33317),
            .I(N__33307));
    InMux I__6199 (
            .O(N__33316),
            .I(N__33304));
    LocalMux I__6198 (
            .O(N__33313),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__6197 (
            .O(N__33310),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__6196 (
            .O(N__33307),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__6195 (
            .O(N__33304),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    IoInMux I__6194 (
            .O(N__33295),
            .I(N__33292));
    LocalMux I__6193 (
            .O(N__33292),
            .I(N__33289));
    Odrv4 I__6192 (
            .O(N__33289),
            .I(\current_shift_inst.timer_s1.N_180_i ));
    InMux I__6191 (
            .O(N__33286),
            .I(N__33280));
    InMux I__6190 (
            .O(N__33285),
            .I(N__33280));
    LocalMux I__6189 (
            .O(N__33280),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9 ));
    InMux I__6188 (
            .O(N__33277),
            .I(N__33274));
    LocalMux I__6187 (
            .O(N__33274),
            .I(N__33271));
    Sp12to4 I__6186 (
            .O(N__33271),
            .I(N__33268));
    Odrv12 I__6185 (
            .O(N__33268),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17 ));
    InMux I__6184 (
            .O(N__33265),
            .I(N__33262));
    LocalMux I__6183 (
            .O(N__33262),
            .I(N__33259));
    Span4Mux_h I__6182 (
            .O(N__33259),
            .I(N__33255));
    InMux I__6181 (
            .O(N__33258),
            .I(N__33252));
    Odrv4 I__6180 (
            .O(N__33255),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_0 ));
    LocalMux I__6179 (
            .O(N__33252),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_0 ));
    InMux I__6178 (
            .O(N__33247),
            .I(N__33244));
    LocalMux I__6177 (
            .O(N__33244),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_0 ));
    InMux I__6176 (
            .O(N__33241),
            .I(N__33238));
    LocalMux I__6175 (
            .O(N__33238),
            .I(N__33234));
    InMux I__6174 (
            .O(N__33237),
            .I(N__33231));
    Span4Mux_h I__6173 (
            .O(N__33234),
            .I(N__33228));
    LocalMux I__6172 (
            .O(N__33231),
            .I(N__33225));
    Odrv4 I__6171 (
            .O(N__33228),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_1 ));
    Odrv4 I__6170 (
            .O(N__33225),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_1 ));
    InMux I__6169 (
            .O(N__33220),
            .I(N__33217));
    LocalMux I__6168 (
            .O(N__33217),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_1 ));
    InMux I__6167 (
            .O(N__33214),
            .I(N__33211));
    LocalMux I__6166 (
            .O(N__33211),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9 ));
    InMux I__6165 (
            .O(N__33208),
            .I(N__33205));
    LocalMux I__6164 (
            .O(N__33205),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt8 ));
    CascadeMux I__6163 (
            .O(N__33202),
            .I(N__33199));
    InMux I__6162 (
            .O(N__33199),
            .I(N__33195));
    InMux I__6161 (
            .O(N__33198),
            .I(N__33192));
    LocalMux I__6160 (
            .O(N__33195),
            .I(N__33189));
    LocalMux I__6159 (
            .O(N__33192),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1 ));
    Odrv4 I__6158 (
            .O(N__33189),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1 ));
    CascadeMux I__6157 (
            .O(N__33184),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt13_cascade_ ));
    CascadeMux I__6156 (
            .O(N__33181),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt19_0_cascade_ ));
    InMux I__6155 (
            .O(N__33178),
            .I(N__33172));
    InMux I__6154 (
            .O(N__33177),
            .I(N__33169));
    InMux I__6153 (
            .O(N__33176),
            .I(N__33166));
    InMux I__6152 (
            .O(N__33175),
            .I(N__33163));
    LocalMux I__6151 (
            .O(N__33172),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    LocalMux I__6150 (
            .O(N__33169),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    LocalMux I__6149 (
            .O(N__33166),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    LocalMux I__6148 (
            .O(N__33163),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    CascadeMux I__6147 (
            .O(N__33154),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2_cascade_ ));
    InMux I__6146 (
            .O(N__33151),
            .I(N__33148));
    LocalMux I__6145 (
            .O(N__33148),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_2 ));
    InMux I__6144 (
            .O(N__33145),
            .I(N__33142));
    LocalMux I__6143 (
            .O(N__33142),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8 ));
    CascadeMux I__6142 (
            .O(N__33139),
            .I(N__33136));
    InMux I__6141 (
            .O(N__33136),
            .I(N__33131));
    CascadeMux I__6140 (
            .O(N__33135),
            .I(N__33128));
    CascadeMux I__6139 (
            .O(N__33134),
            .I(N__33125));
    LocalMux I__6138 (
            .O(N__33131),
            .I(N__33122));
    InMux I__6137 (
            .O(N__33128),
            .I(N__33119));
    InMux I__6136 (
            .O(N__33125),
            .I(N__33116));
    Span4Mux_v I__6135 (
            .O(N__33122),
            .I(N__33113));
    LocalMux I__6134 (
            .O(N__33119),
            .I(N__33110));
    LocalMux I__6133 (
            .O(N__33116),
            .I(measured_delay_hc_19));
    Odrv4 I__6132 (
            .O(N__33113),
            .I(measured_delay_hc_19));
    Odrv12 I__6131 (
            .O(N__33110),
            .I(measured_delay_hc_19));
    CascadeMux I__6130 (
            .O(N__33103),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto5_2_cascade_ ));
    CascadeMux I__6129 (
            .O(N__33100),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8_cascade_ ));
    CascadeMux I__6128 (
            .O(N__33097),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclt31_0_cascade_ ));
    InMux I__6127 (
            .O(N__33094),
            .I(N__33091));
    LocalMux I__6126 (
            .O(N__33091),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_7 ));
    InMux I__6125 (
            .O(N__33088),
            .I(N__33085));
    LocalMux I__6124 (
            .O(N__33085),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt13_0 ));
    InMux I__6123 (
            .O(N__33082),
            .I(N__33079));
    LocalMux I__6122 (
            .O(N__33079),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt19 ));
    InMux I__6121 (
            .O(N__33076),
            .I(N__33072));
    InMux I__6120 (
            .O(N__33075),
            .I(N__33069));
    LocalMux I__6119 (
            .O(N__33072),
            .I(N__33062));
    LocalMux I__6118 (
            .O(N__33069),
            .I(N__33062));
    InMux I__6117 (
            .O(N__33068),
            .I(N__33059));
    InMux I__6116 (
            .O(N__33067),
            .I(N__33056));
    Span4Mux_v I__6115 (
            .O(N__33062),
            .I(N__33053));
    LocalMux I__6114 (
            .O(N__33059),
            .I(N__33050));
    LocalMux I__6113 (
            .O(N__33056),
            .I(measured_delay_hc_0));
    Odrv4 I__6112 (
            .O(N__33053),
            .I(measured_delay_hc_0));
    Odrv4 I__6111 (
            .O(N__33050),
            .I(measured_delay_hc_0));
    InMux I__6110 (
            .O(N__33043),
            .I(N__33038));
    InMux I__6109 (
            .O(N__33042),
            .I(N__33033));
    InMux I__6108 (
            .O(N__33041),
            .I(N__33033));
    LocalMux I__6107 (
            .O(N__33038),
            .I(measured_delay_hc_20));
    LocalMux I__6106 (
            .O(N__33033),
            .I(measured_delay_hc_20));
    CascadeMux I__6105 (
            .O(N__33028),
            .I(N__33022));
    InMux I__6104 (
            .O(N__33027),
            .I(N__33018));
    InMux I__6103 (
            .O(N__33026),
            .I(N__33015));
    InMux I__6102 (
            .O(N__33025),
            .I(N__33010));
    InMux I__6101 (
            .O(N__33022),
            .I(N__33010));
    CascadeMux I__6100 (
            .O(N__33021),
            .I(N__33007));
    LocalMux I__6099 (
            .O(N__33018),
            .I(N__33004));
    LocalMux I__6098 (
            .O(N__33015),
            .I(N__32999));
    LocalMux I__6097 (
            .O(N__33010),
            .I(N__32999));
    InMux I__6096 (
            .O(N__33007),
            .I(N__32996));
    Span4Mux_h I__6095 (
            .O(N__33004),
            .I(N__32993));
    Span4Mux_h I__6094 (
            .O(N__32999),
            .I(N__32990));
    LocalMux I__6093 (
            .O(N__32996),
            .I(measured_delay_hc_16));
    Odrv4 I__6092 (
            .O(N__32993),
            .I(measured_delay_hc_16));
    Odrv4 I__6091 (
            .O(N__32990),
            .I(measured_delay_hc_16));
    InMux I__6090 (
            .O(N__32983),
            .I(N__32978));
    InMux I__6089 (
            .O(N__32982),
            .I(N__32975));
    CascadeMux I__6088 (
            .O(N__32981),
            .I(N__32971));
    LocalMux I__6087 (
            .O(N__32978),
            .I(N__32966));
    LocalMux I__6086 (
            .O(N__32975),
            .I(N__32966));
    InMux I__6085 (
            .O(N__32974),
            .I(N__32963));
    InMux I__6084 (
            .O(N__32971),
            .I(N__32960));
    Span4Mux_h I__6083 (
            .O(N__32966),
            .I(N__32957));
    LocalMux I__6082 (
            .O(N__32963),
            .I(N__32954));
    LocalMux I__6081 (
            .O(N__32960),
            .I(measured_delay_hc_1));
    Odrv4 I__6080 (
            .O(N__32957),
            .I(measured_delay_hc_1));
    Odrv4 I__6079 (
            .O(N__32954),
            .I(measured_delay_hc_1));
    InMux I__6078 (
            .O(N__32947),
            .I(N__32943));
    InMux I__6077 (
            .O(N__32946),
            .I(N__32940));
    LocalMux I__6076 (
            .O(N__32943),
            .I(N__32935));
    LocalMux I__6075 (
            .O(N__32940),
            .I(N__32932));
    InMux I__6074 (
            .O(N__32939),
            .I(N__32929));
    InMux I__6073 (
            .O(N__32938),
            .I(N__32926));
    Span4Mux_h I__6072 (
            .O(N__32935),
            .I(N__32923));
    Span4Mux_v I__6071 (
            .O(N__32932),
            .I(N__32918));
    LocalMux I__6070 (
            .O(N__32929),
            .I(N__32918));
    LocalMux I__6069 (
            .O(N__32926),
            .I(measured_delay_hc_8));
    Odrv4 I__6068 (
            .O(N__32923),
            .I(measured_delay_hc_8));
    Odrv4 I__6067 (
            .O(N__32918),
            .I(measured_delay_hc_8));
    InMux I__6066 (
            .O(N__32911),
            .I(N__32904));
    InMux I__6065 (
            .O(N__32910),
            .I(N__32904));
    InMux I__6064 (
            .O(N__32909),
            .I(N__32901));
    LocalMux I__6063 (
            .O(N__32904),
            .I(N__32898));
    LocalMux I__6062 (
            .O(N__32901),
            .I(measured_delay_hc_21));
    Odrv4 I__6061 (
            .O(N__32898),
            .I(measured_delay_hc_21));
    InMux I__6060 (
            .O(N__32893),
            .I(N__32886));
    InMux I__6059 (
            .O(N__32892),
            .I(N__32883));
    InMux I__6058 (
            .O(N__32891),
            .I(N__32880));
    InMux I__6057 (
            .O(N__32890),
            .I(N__32877));
    CascadeMux I__6056 (
            .O(N__32889),
            .I(N__32874));
    LocalMux I__6055 (
            .O(N__32886),
            .I(N__32871));
    LocalMux I__6054 (
            .O(N__32883),
            .I(N__32868));
    LocalMux I__6053 (
            .O(N__32880),
            .I(N__32865));
    LocalMux I__6052 (
            .O(N__32877),
            .I(N__32862));
    InMux I__6051 (
            .O(N__32874),
            .I(N__32859));
    Span4Mux_h I__6050 (
            .O(N__32871),
            .I(N__32856));
    Span4Mux_v I__6049 (
            .O(N__32868),
            .I(N__32851));
    Span4Mux_v I__6048 (
            .O(N__32865),
            .I(N__32851));
    Span4Mux_h I__6047 (
            .O(N__32862),
            .I(N__32848));
    LocalMux I__6046 (
            .O(N__32859),
            .I(measured_delay_hc_15));
    Odrv4 I__6045 (
            .O(N__32856),
            .I(measured_delay_hc_15));
    Odrv4 I__6044 (
            .O(N__32851),
            .I(measured_delay_hc_15));
    Odrv4 I__6043 (
            .O(N__32848),
            .I(measured_delay_hc_15));
    InMux I__6042 (
            .O(N__32839),
            .I(N__32836));
    LocalMux I__6041 (
            .O(N__32836),
            .I(N__32831));
    InMux I__6040 (
            .O(N__32835),
            .I(N__32828));
    InMux I__6039 (
            .O(N__32834),
            .I(N__32824));
    Span4Mux_h I__6038 (
            .O(N__32831),
            .I(N__32818));
    LocalMux I__6037 (
            .O(N__32828),
            .I(N__32818));
    InMux I__6036 (
            .O(N__32827),
            .I(N__32815));
    LocalMux I__6035 (
            .O(N__32824),
            .I(N__32812));
    InMux I__6034 (
            .O(N__32823),
            .I(N__32809));
    Span4Mux_v I__6033 (
            .O(N__32818),
            .I(N__32802));
    LocalMux I__6032 (
            .O(N__32815),
            .I(N__32802));
    Span4Mux_h I__6031 (
            .O(N__32812),
            .I(N__32802));
    LocalMux I__6030 (
            .O(N__32809),
            .I(measured_delay_hc_4));
    Odrv4 I__6029 (
            .O(N__32802),
            .I(measured_delay_hc_4));
    CascadeMux I__6028 (
            .O(N__32797),
            .I(N__32793));
    CascadeMux I__6027 (
            .O(N__32796),
            .I(N__32790));
    InMux I__6026 (
            .O(N__32793),
            .I(N__32787));
    InMux I__6025 (
            .O(N__32790),
            .I(N__32784));
    LocalMux I__6024 (
            .O(N__32787),
            .I(N__32779));
    LocalMux I__6023 (
            .O(N__32784),
            .I(N__32779));
    Span4Mux_h I__6022 (
            .O(N__32779),
            .I(N__32774));
    InMux I__6021 (
            .O(N__32778),
            .I(N__32771));
    InMux I__6020 (
            .O(N__32777),
            .I(N__32768));
    Sp12to4 I__6019 (
            .O(N__32774),
            .I(N__32763));
    LocalMux I__6018 (
            .O(N__32771),
            .I(N__32763));
    LocalMux I__6017 (
            .O(N__32768),
            .I(measured_delay_hc_2));
    Odrv12 I__6016 (
            .O(N__32763),
            .I(measured_delay_hc_2));
    InMux I__6015 (
            .O(N__32758),
            .I(\current_shift_inst.un38_control_input_cry_26_s0 ));
    InMux I__6014 (
            .O(N__32755),
            .I(\current_shift_inst.un38_control_input_cry_27_s0 ));
    InMux I__6013 (
            .O(N__32752),
            .I(\current_shift_inst.un38_control_input_cry_28_s0 ));
    InMux I__6012 (
            .O(N__32749),
            .I(\current_shift_inst.un38_control_input_cry_29_s0 ));
    InMux I__6011 (
            .O(N__32746),
            .I(\current_shift_inst.un38_control_input_cry_30_s0 ));
    InMux I__6010 (
            .O(N__32743),
            .I(N__32737));
    InMux I__6009 (
            .O(N__32742),
            .I(N__32737));
    LocalMux I__6008 (
            .O(N__32737),
            .I(N__32734));
    Odrv4 I__6007 (
            .O(N__32734),
            .I(\phase_controller_inst1.stoper_hc.un2_startlt3 ));
    InMux I__6006 (
            .O(N__32731),
            .I(N__32727));
    InMux I__6005 (
            .O(N__32730),
            .I(N__32724));
    LocalMux I__6004 (
            .O(N__32727),
            .I(N__32721));
    LocalMux I__6003 (
            .O(N__32724),
            .I(N__32718));
    Span4Mux_h I__6002 (
            .O(N__32721),
            .I(N__32714));
    Span4Mux_h I__6001 (
            .O(N__32718),
            .I(N__32711));
    InMux I__6000 (
            .O(N__32717),
            .I(N__32708));
    Odrv4 I__5999 (
            .O(N__32714),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1 ));
    Odrv4 I__5998 (
            .O(N__32711),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1 ));
    LocalMux I__5997 (
            .O(N__32708),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1 ));
    InMux I__5996 (
            .O(N__32701),
            .I(N__32698));
    LocalMux I__5995 (
            .O(N__32698),
            .I(N__32695));
    Odrv4 I__5994 (
            .O(N__32695),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_6 ));
    CascadeMux I__5993 (
            .O(N__32692),
            .I(N__32687));
    InMux I__5992 (
            .O(N__32691),
            .I(N__32684));
    InMux I__5991 (
            .O(N__32690),
            .I(N__32679));
    InMux I__5990 (
            .O(N__32687),
            .I(N__32679));
    LocalMux I__5989 (
            .O(N__32684),
            .I(measured_delay_hc_22));
    LocalMux I__5988 (
            .O(N__32679),
            .I(measured_delay_hc_22));
    InMux I__5987 (
            .O(N__32674),
            .I(N__32669));
    InMux I__5986 (
            .O(N__32673),
            .I(N__32666));
    CascadeMux I__5985 (
            .O(N__32672),
            .I(N__32663));
    LocalMux I__5984 (
            .O(N__32669),
            .I(N__32660));
    LocalMux I__5983 (
            .O(N__32666),
            .I(N__32657));
    InMux I__5982 (
            .O(N__32663),
            .I(N__32653));
    Span4Mux_v I__5981 (
            .O(N__32660),
            .I(N__32650));
    Span4Mux_h I__5980 (
            .O(N__32657),
            .I(N__32647));
    InMux I__5979 (
            .O(N__32656),
            .I(N__32644));
    LocalMux I__5978 (
            .O(N__32653),
            .I(measured_delay_hc_7));
    Odrv4 I__5977 (
            .O(N__32650),
            .I(measured_delay_hc_7));
    Odrv4 I__5976 (
            .O(N__32647),
            .I(measured_delay_hc_7));
    LocalMux I__5975 (
            .O(N__32644),
            .I(measured_delay_hc_7));
    InMux I__5974 (
            .O(N__32635),
            .I(N__32632));
    LocalMux I__5973 (
            .O(N__32632),
            .I(N__32629));
    Span4Mux_v I__5972 (
            .O(N__32629),
            .I(N__32626));
    Odrv4 I__5971 (
            .O(N__32626),
            .I(\current_shift_inst.un38_control_input_0_s0_19 ));
    InMux I__5970 (
            .O(N__32623),
            .I(\current_shift_inst.un38_control_input_cry_18_s0 ));
    InMux I__5969 (
            .O(N__32620),
            .I(N__32617));
    LocalMux I__5968 (
            .O(N__32617),
            .I(N__32614));
    Odrv12 I__5967 (
            .O(N__32614),
            .I(\current_shift_inst.un38_control_input_0_s0_20 ));
    InMux I__5966 (
            .O(N__32611),
            .I(\current_shift_inst.un38_control_input_cry_19_s0 ));
    InMux I__5965 (
            .O(N__32608),
            .I(N__32605));
    LocalMux I__5964 (
            .O(N__32605),
            .I(N__32602));
    Odrv12 I__5963 (
            .O(N__32602),
            .I(\current_shift_inst.un38_control_input_0_s0_21 ));
    InMux I__5962 (
            .O(N__32599),
            .I(\current_shift_inst.un38_control_input_cry_20_s0 ));
    CascadeMux I__5961 (
            .O(N__32596),
            .I(N__32593));
    InMux I__5960 (
            .O(N__32593),
            .I(N__32590));
    LocalMux I__5959 (
            .O(N__32590),
            .I(N__32587));
    Odrv12 I__5958 (
            .O(N__32587),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ));
    InMux I__5957 (
            .O(N__32584),
            .I(\current_shift_inst.un38_control_input_cry_21_s0 ));
    InMux I__5956 (
            .O(N__32581),
            .I(N__32578));
    LocalMux I__5955 (
            .O(N__32578),
            .I(N__32575));
    Odrv12 I__5954 (
            .O(N__32575),
            .I(\current_shift_inst.un38_control_input_0_s0_23 ));
    InMux I__5953 (
            .O(N__32572),
            .I(\current_shift_inst.un38_control_input_cry_22_s0 ));
    InMux I__5952 (
            .O(N__32569),
            .I(bfn_13_20_0_));
    InMux I__5951 (
            .O(N__32566),
            .I(\current_shift_inst.un38_control_input_cry_24_s0 ));
    InMux I__5950 (
            .O(N__32563),
            .I(\current_shift_inst.un38_control_input_cry_25_s0 ));
    InMux I__5949 (
            .O(N__32560),
            .I(\current_shift_inst.un38_control_input_cry_9_s0 ));
    InMux I__5948 (
            .O(N__32557),
            .I(\current_shift_inst.un38_control_input_cry_10_s0 ));
    InMux I__5947 (
            .O(N__32554),
            .I(N__32551));
    LocalMux I__5946 (
            .O(N__32551),
            .I(N__32548));
    Odrv12 I__5945 (
            .O(N__32548),
            .I(\current_shift_inst.un38_control_input_0_s0_12 ));
    InMux I__5944 (
            .O(N__32545),
            .I(\current_shift_inst.un38_control_input_cry_11_s0 ));
    InMux I__5943 (
            .O(N__32542),
            .I(N__32539));
    LocalMux I__5942 (
            .O(N__32539),
            .I(N__32536));
    Odrv12 I__5941 (
            .O(N__32536),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14 ));
    InMux I__5940 (
            .O(N__32533),
            .I(\current_shift_inst.un38_control_input_cry_12_s0 ));
    InMux I__5939 (
            .O(N__32530),
            .I(N__32527));
    LocalMux I__5938 (
            .O(N__32527),
            .I(N__32524));
    Odrv4 I__5937 (
            .O(N__32524),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15 ));
    InMux I__5936 (
            .O(N__32521),
            .I(N__32518));
    LocalMux I__5935 (
            .O(N__32518),
            .I(N__32515));
    Odrv12 I__5934 (
            .O(N__32515),
            .I(\current_shift_inst.un38_control_input_0_s0_14 ));
    InMux I__5933 (
            .O(N__32512),
            .I(\current_shift_inst.un38_control_input_cry_13_s0 ));
    InMux I__5932 (
            .O(N__32509),
            .I(N__32506));
    LocalMux I__5931 (
            .O(N__32506),
            .I(N__32503));
    Odrv12 I__5930 (
            .O(N__32503),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16 ));
    InMux I__5929 (
            .O(N__32500),
            .I(N__32497));
    LocalMux I__5928 (
            .O(N__32497),
            .I(N__32494));
    Odrv4 I__5927 (
            .O(N__32494),
            .I(\current_shift_inst.un38_control_input_0_s0_15 ));
    InMux I__5926 (
            .O(N__32491),
            .I(\current_shift_inst.un38_control_input_cry_14_s0 ));
    InMux I__5925 (
            .O(N__32488),
            .I(N__32485));
    LocalMux I__5924 (
            .O(N__32485),
            .I(N__32482));
    Span4Mux_v I__5923 (
            .O(N__32482),
            .I(N__32479));
    Odrv4 I__5922 (
            .O(N__32479),
            .I(\current_shift_inst.un38_control_input_0_s0_16 ));
    InMux I__5921 (
            .O(N__32476),
            .I(bfn_13_19_0_));
    InMux I__5920 (
            .O(N__32473),
            .I(N__32470));
    LocalMux I__5919 (
            .O(N__32470),
            .I(N__32467));
    Span4Mux_h I__5918 (
            .O(N__32467),
            .I(N__32464));
    Odrv4 I__5917 (
            .O(N__32464),
            .I(\current_shift_inst.un38_control_input_0_s0_17 ));
    InMux I__5916 (
            .O(N__32461),
            .I(\current_shift_inst.un38_control_input_cry_16_s0 ));
    InMux I__5915 (
            .O(N__32458),
            .I(N__32455));
    LocalMux I__5914 (
            .O(N__32455),
            .I(N__32452));
    Odrv12 I__5913 (
            .O(N__32452),
            .I(\current_shift_inst.un38_control_input_0_s0_18 ));
    InMux I__5912 (
            .O(N__32449),
            .I(\current_shift_inst.un38_control_input_cry_17_s0 ));
    InMux I__5911 (
            .O(N__32446),
            .I(N__32443));
    LocalMux I__5910 (
            .O(N__32443),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ));
    InMux I__5909 (
            .O(N__32440),
            .I(N__32437));
    LocalMux I__5908 (
            .O(N__32437),
            .I(N__32434));
    Odrv4 I__5907 (
            .O(N__32434),
            .I(\current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0 ));
    InMux I__5906 (
            .O(N__32431),
            .I(\current_shift_inst.un38_control_input_cry_5_s0 ));
    InMux I__5905 (
            .O(N__32428),
            .I(N__32425));
    LocalMux I__5904 (
            .O(N__32425),
            .I(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8 ));
    InMux I__5903 (
            .O(N__32422),
            .I(\current_shift_inst.un38_control_input_cry_6_s0 ));
    InMux I__5902 (
            .O(N__32419),
            .I(N__32416));
    LocalMux I__5901 (
            .O(N__32416),
            .I(N__32413));
    Odrv4 I__5900 (
            .O(N__32413),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9 ));
    InMux I__5899 (
            .O(N__32410),
            .I(N__32407));
    LocalMux I__5898 (
            .O(N__32407),
            .I(N__32404));
    Odrv4 I__5897 (
            .O(N__32404),
            .I(\current_shift_inst.un38_control_input_0_s0_8 ));
    InMux I__5896 (
            .O(N__32401),
            .I(bfn_13_18_0_));
    InMux I__5895 (
            .O(N__32398),
            .I(N__32395));
    LocalMux I__5894 (
            .O(N__32395),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10 ));
    InMux I__5893 (
            .O(N__32392),
            .I(N__32389));
    LocalMux I__5892 (
            .O(N__32389),
            .I(N__32386));
    Odrv4 I__5891 (
            .O(N__32386),
            .I(\current_shift_inst.un38_control_input_0_s0_9 ));
    InMux I__5890 (
            .O(N__32383),
            .I(\current_shift_inst.un38_control_input_cry_8_s0 ));
    InMux I__5889 (
            .O(N__32380),
            .I(N__32377));
    LocalMux I__5888 (
            .O(N__32377),
            .I(N__32374));
    Odrv4 I__5887 (
            .O(N__32374),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11 ));
    InMux I__5886 (
            .O(N__32371),
            .I(N__32368));
    LocalMux I__5885 (
            .O(N__32368),
            .I(N__32365));
    Odrv4 I__5884 (
            .O(N__32365),
            .I(\current_shift_inst.un38_control_input_0_s0_10 ));
    InMux I__5883 (
            .O(N__32362),
            .I(N__32359));
    LocalMux I__5882 (
            .O(N__32359),
            .I(\current_shift_inst.un38_control_input_cry_0_s0_sf ));
    InMux I__5881 (
            .O(N__32356),
            .I(N__32353));
    LocalMux I__5880 (
            .O(N__32353),
            .I(N__32350));
    Odrv12 I__5879 (
            .O(N__32350),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ));
    InMux I__5878 (
            .O(N__32347),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_24 ));
    InMux I__5877 (
            .O(N__32344),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_25 ));
    InMux I__5876 (
            .O(N__32341),
            .I(N__32338));
    LocalMux I__5875 (
            .O(N__32338),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25 ));
    InMux I__5874 (
            .O(N__32335),
            .I(N__32332));
    LocalMux I__5873 (
            .O(N__32332),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24 ));
    InMux I__5872 (
            .O(N__32329),
            .I(N__32326));
    LocalMux I__5871 (
            .O(N__32326),
            .I(N__32323));
    Odrv4 I__5870 (
            .O(N__32323),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21 ));
    InMux I__5869 (
            .O(N__32320),
            .I(bfn_13_12_0_));
    InMux I__5868 (
            .O(N__32317),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_16 ));
    InMux I__5867 (
            .O(N__32314),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_17 ));
    InMux I__5866 (
            .O(N__32311),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_18 ));
    InMux I__5865 (
            .O(N__32308),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_19 ));
    InMux I__5864 (
            .O(N__32305),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_20 ));
    InMux I__5863 (
            .O(N__32302),
            .I(N__32299));
    LocalMux I__5862 (
            .O(N__32299),
            .I(N__32296));
    Span4Mux_v I__5861 (
            .O(N__32296),
            .I(N__32293));
    Odrv4 I__5860 (
            .O(N__32293),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22 ));
    InMux I__5859 (
            .O(N__32290),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_21 ));
    InMux I__5858 (
            .O(N__32287),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_22 ));
    InMux I__5857 (
            .O(N__32284),
            .I(bfn_13_13_0_));
    InMux I__5856 (
            .O(N__32281),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ));
    InMux I__5855 (
            .O(N__32278),
            .I(bfn_13_11_0_));
    InMux I__5854 (
            .O(N__32275),
            .I(N__32272));
    LocalMux I__5853 (
            .O(N__32272),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ));
    InMux I__5852 (
            .O(N__32269),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ));
    InMux I__5851 (
            .O(N__32266),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ));
    InMux I__5850 (
            .O(N__32263),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ));
    InMux I__5849 (
            .O(N__32260),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ));
    InMux I__5848 (
            .O(N__32257),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ));
    InMux I__5847 (
            .O(N__32254),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ));
    InMux I__5846 (
            .O(N__32251),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_14 ));
    InMux I__5845 (
            .O(N__32248),
            .I(N__32245));
    LocalMux I__5844 (
            .O(N__32245),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ));
    InMux I__5843 (
            .O(N__32242),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ));
    InMux I__5842 (
            .O(N__32239),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ));
    InMux I__5841 (
            .O(N__32236),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ));
    InMux I__5840 (
            .O(N__32233),
            .I(N__32230));
    LocalMux I__5839 (
            .O(N__32230),
            .I(N__32227));
    Span4Mux_h I__5838 (
            .O(N__32227),
            .I(N__32224));
    Odrv4 I__5837 (
            .O(N__32224),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ));
    InMux I__5836 (
            .O(N__32221),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ));
    InMux I__5835 (
            .O(N__32218),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ));
    InMux I__5834 (
            .O(N__32215),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ));
    CascadeMux I__5833 (
            .O(N__32212),
            .I(N__32208));
    CascadeMux I__5832 (
            .O(N__32211),
            .I(N__32205));
    InMux I__5831 (
            .O(N__32208),
            .I(N__32202));
    InMux I__5830 (
            .O(N__32205),
            .I(N__32198));
    LocalMux I__5829 (
            .O(N__32202),
            .I(N__32195));
    InMux I__5828 (
            .O(N__32201),
            .I(N__32192));
    LocalMux I__5827 (
            .O(N__32198),
            .I(N__32188));
    Span4Mux_h I__5826 (
            .O(N__32195),
            .I(N__32183));
    LocalMux I__5825 (
            .O(N__32192),
            .I(N__32183));
    InMux I__5824 (
            .O(N__32191),
            .I(N__32180));
    Span4Mux_h I__5823 (
            .O(N__32188),
            .I(N__32177));
    Span4Mux_v I__5822 (
            .O(N__32183),
            .I(N__32174));
    LocalMux I__5821 (
            .O(N__32180),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    Odrv4 I__5820 (
            .O(N__32177),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    Odrv4 I__5819 (
            .O(N__32174),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    InMux I__5818 (
            .O(N__32167),
            .I(N__32163));
    InMux I__5817 (
            .O(N__32166),
            .I(N__32160));
    LocalMux I__5816 (
            .O(N__32163),
            .I(measured_delay_hc_23));
    LocalMux I__5815 (
            .O(N__32160),
            .I(measured_delay_hc_23));
    InMux I__5814 (
            .O(N__32155),
            .I(N__32151));
    InMux I__5813 (
            .O(N__32154),
            .I(N__32148));
    LocalMux I__5812 (
            .O(N__32151),
            .I(N__32144));
    LocalMux I__5811 (
            .O(N__32148),
            .I(N__32141));
    InMux I__5810 (
            .O(N__32147),
            .I(N__32138));
    Span4Mux_s3_v I__5809 (
            .O(N__32144),
            .I(N__32135));
    Span4Mux_s3_v I__5808 (
            .O(N__32141),
            .I(N__32132));
    LocalMux I__5807 (
            .O(N__32138),
            .I(N__32129));
    Span4Mux_v I__5806 (
            .O(N__32135),
            .I(N__32126));
    Span4Mux_v I__5805 (
            .O(N__32132),
            .I(N__32123));
    Span12Mux_h I__5804 (
            .O(N__32129),
            .I(N__32117));
    Sp12to4 I__5803 (
            .O(N__32126),
            .I(N__32112));
    Sp12to4 I__5802 (
            .O(N__32123),
            .I(N__32112));
    InMux I__5801 (
            .O(N__32122),
            .I(N__32109));
    InMux I__5800 (
            .O(N__32121),
            .I(N__32104));
    InMux I__5799 (
            .O(N__32120),
            .I(N__32104));
    Span12Mux_v I__5798 (
            .O(N__32117),
            .I(N__32101));
    Span12Mux_h I__5797 (
            .O(N__32112),
            .I(N__32096));
    LocalMux I__5796 (
            .O(N__32109),
            .I(N__32096));
    LocalMux I__5795 (
            .O(N__32104),
            .I(state_3));
    Odrv12 I__5794 (
            .O(N__32101),
            .I(state_3));
    Odrv12 I__5793 (
            .O(N__32096),
            .I(state_3));
    IoInMux I__5792 (
            .O(N__32089),
            .I(N__32086));
    LocalMux I__5791 (
            .O(N__32086),
            .I(N__32083));
    Span4Mux_s2_v I__5790 (
            .O(N__32083),
            .I(N__32079));
    CascadeMux I__5789 (
            .O(N__32082),
            .I(N__32076));
    Span4Mux_h I__5788 (
            .O(N__32079),
            .I(N__32072));
    InMux I__5787 (
            .O(N__32076),
            .I(N__32069));
    InMux I__5786 (
            .O(N__32075),
            .I(N__32066));
    Odrv4 I__5785 (
            .O(N__32072),
            .I(s1_phy_c));
    LocalMux I__5784 (
            .O(N__32069),
            .I(s1_phy_c));
    LocalMux I__5783 (
            .O(N__32066),
            .I(s1_phy_c));
    CascadeMux I__5782 (
            .O(N__32059),
            .I(N__32056));
    InMux I__5781 (
            .O(N__32056),
            .I(N__32053));
    LocalMux I__5780 (
            .O(N__32053),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_11 ));
    CascadeMux I__5779 (
            .O(N__32050),
            .I(\current_shift_inst.PI_CTRL.un1_enablelt3_0_cascade_ ));
    InMux I__5778 (
            .O(N__32047),
            .I(N__32044));
    LocalMux I__5777 (
            .O(N__32044),
            .I(N__32041));
    Odrv4 I__5776 (
            .O(N__32041),
            .I(\current_shift_inst.PI_CTRL.N_71 ));
    CascadeMux I__5775 (
            .O(N__32038),
            .I(N__32031));
    InMux I__5774 (
            .O(N__32037),
            .I(N__32028));
    InMux I__5773 (
            .O(N__32036),
            .I(N__32025));
    InMux I__5772 (
            .O(N__32035),
            .I(N__32020));
    InMux I__5771 (
            .O(N__32034),
            .I(N__32020));
    InMux I__5770 (
            .O(N__32031),
            .I(N__32017));
    LocalMux I__5769 (
            .O(N__32028),
            .I(N__32014));
    LocalMux I__5768 (
            .O(N__32025),
            .I(N__32009));
    LocalMux I__5767 (
            .O(N__32020),
            .I(N__32009));
    LocalMux I__5766 (
            .O(N__32017),
            .I(measured_delay_hc_11));
    Odrv12 I__5765 (
            .O(N__32014),
            .I(measured_delay_hc_11));
    Odrv4 I__5764 (
            .O(N__32009),
            .I(measured_delay_hc_11));
    CascadeMux I__5763 (
            .O(N__32002),
            .I(N__31997));
    InMux I__5762 (
            .O(N__32001),
            .I(N__31993));
    InMux I__5761 (
            .O(N__32000),
            .I(N__31987));
    InMux I__5760 (
            .O(N__31997),
            .I(N__31987));
    CascadeMux I__5759 (
            .O(N__31996),
            .I(N__31984));
    LocalMux I__5758 (
            .O(N__31993),
            .I(N__31981));
    InMux I__5757 (
            .O(N__31992),
            .I(N__31978));
    LocalMux I__5756 (
            .O(N__31987),
            .I(N__31975));
    InMux I__5755 (
            .O(N__31984),
            .I(N__31972));
    Span12Mux_v I__5754 (
            .O(N__31981),
            .I(N__31969));
    LocalMux I__5753 (
            .O(N__31978),
            .I(N__31964));
    Span4Mux_h I__5752 (
            .O(N__31975),
            .I(N__31964));
    LocalMux I__5751 (
            .O(N__31972),
            .I(measured_delay_hc_9));
    Odrv12 I__5750 (
            .O(N__31969),
            .I(measured_delay_hc_9));
    Odrv4 I__5749 (
            .O(N__31964),
            .I(measured_delay_hc_9));
    InMux I__5748 (
            .O(N__31957),
            .I(N__31954));
    LocalMux I__5747 (
            .O(N__31954),
            .I(N__31948));
    CascadeMux I__5746 (
            .O(N__31953),
            .I(N__31945));
    InMux I__5745 (
            .O(N__31952),
            .I(N__31942));
    CascadeMux I__5744 (
            .O(N__31951),
            .I(N__31938));
    Span4Mux_h I__5743 (
            .O(N__31948),
            .I(N__31935));
    InMux I__5742 (
            .O(N__31945),
            .I(N__31932));
    LocalMux I__5741 (
            .O(N__31942),
            .I(N__31929));
    InMux I__5740 (
            .O(N__31941),
            .I(N__31926));
    InMux I__5739 (
            .O(N__31938),
            .I(N__31923));
    Span4Mux_v I__5738 (
            .O(N__31935),
            .I(N__31920));
    LocalMux I__5737 (
            .O(N__31932),
            .I(N__31915));
    Span4Mux_h I__5736 (
            .O(N__31929),
            .I(N__31915));
    LocalMux I__5735 (
            .O(N__31926),
            .I(N__31912));
    LocalMux I__5734 (
            .O(N__31923),
            .I(measured_delay_hc_14));
    Odrv4 I__5733 (
            .O(N__31920),
            .I(measured_delay_hc_14));
    Odrv4 I__5732 (
            .O(N__31915),
            .I(measured_delay_hc_14));
    Odrv12 I__5731 (
            .O(N__31912),
            .I(measured_delay_hc_14));
    InMux I__5730 (
            .O(N__31903),
            .I(N__31898));
    CascadeMux I__5729 (
            .O(N__31902),
            .I(N__31894));
    CascadeMux I__5728 (
            .O(N__31901),
            .I(N__31891));
    LocalMux I__5727 (
            .O(N__31898),
            .I(N__31888));
    InMux I__5726 (
            .O(N__31897),
            .I(N__31885));
    InMux I__5725 (
            .O(N__31894),
            .I(N__31880));
    InMux I__5724 (
            .O(N__31891),
            .I(N__31880));
    Span4Mux_h I__5723 (
            .O(N__31888),
            .I(N__31876));
    LocalMux I__5722 (
            .O(N__31885),
            .I(N__31873));
    LocalMux I__5721 (
            .O(N__31880),
            .I(N__31870));
    InMux I__5720 (
            .O(N__31879),
            .I(N__31867));
    Span4Mux_v I__5719 (
            .O(N__31876),
            .I(N__31864));
    Span4Mux_h I__5718 (
            .O(N__31873),
            .I(N__31859));
    Span4Mux_h I__5717 (
            .O(N__31870),
            .I(N__31859));
    LocalMux I__5716 (
            .O(N__31867),
            .I(measured_delay_hc_6));
    Odrv4 I__5715 (
            .O(N__31864),
            .I(measured_delay_hc_6));
    Odrv4 I__5714 (
            .O(N__31859),
            .I(measured_delay_hc_6));
    InMux I__5713 (
            .O(N__31852),
            .I(N__31845));
    InMux I__5712 (
            .O(N__31851),
            .I(N__31842));
    InMux I__5711 (
            .O(N__31850),
            .I(N__31839));
    CascadeMux I__5710 (
            .O(N__31849),
            .I(N__31836));
    CascadeMux I__5709 (
            .O(N__31848),
            .I(N__31833));
    LocalMux I__5708 (
            .O(N__31845),
            .I(N__31830));
    LocalMux I__5707 (
            .O(N__31842),
            .I(N__31825));
    LocalMux I__5706 (
            .O(N__31839),
            .I(N__31825));
    InMux I__5705 (
            .O(N__31836),
            .I(N__31822));
    InMux I__5704 (
            .O(N__31833),
            .I(N__31819));
    Span12Mux_h I__5703 (
            .O(N__31830),
            .I(N__31812));
    Sp12to4 I__5702 (
            .O(N__31825),
            .I(N__31812));
    LocalMux I__5701 (
            .O(N__31822),
            .I(N__31812));
    LocalMux I__5700 (
            .O(N__31819),
            .I(measured_delay_hc_13));
    Odrv12 I__5699 (
            .O(N__31812),
            .I(measured_delay_hc_13));
    InMux I__5698 (
            .O(N__31807),
            .I(N__31803));
    InMux I__5697 (
            .O(N__31806),
            .I(N__31800));
    LocalMux I__5696 (
            .O(N__31803),
            .I(measured_delay_hc_24));
    LocalMux I__5695 (
            .O(N__31800),
            .I(measured_delay_hc_24));
    InMux I__5694 (
            .O(N__31795),
            .I(N__31791));
    InMux I__5693 (
            .O(N__31794),
            .I(N__31788));
    LocalMux I__5692 (
            .O(N__31791),
            .I(measured_delay_hc_25));
    LocalMux I__5691 (
            .O(N__31788),
            .I(measured_delay_hc_25));
    CascadeMux I__5690 (
            .O(N__31783),
            .I(N__31779));
    InMux I__5689 (
            .O(N__31782),
            .I(N__31776));
    InMux I__5688 (
            .O(N__31779),
            .I(N__31773));
    LocalMux I__5687 (
            .O(N__31776),
            .I(measured_delay_hc_26));
    LocalMux I__5686 (
            .O(N__31773),
            .I(measured_delay_hc_26));
    CascadeMux I__5685 (
            .O(N__31768),
            .I(N__31765));
    InMux I__5684 (
            .O(N__31765),
            .I(N__31762));
    LocalMux I__5683 (
            .O(N__31762),
            .I(N__31759));
    Odrv4 I__5682 (
            .O(N__31759),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ));
    InMux I__5681 (
            .O(N__31756),
            .I(N__31720));
    InMux I__5680 (
            .O(N__31755),
            .I(N__31720));
    InMux I__5679 (
            .O(N__31754),
            .I(N__31720));
    InMux I__5678 (
            .O(N__31753),
            .I(N__31720));
    InMux I__5677 (
            .O(N__31752),
            .I(N__31720));
    InMux I__5676 (
            .O(N__31751),
            .I(N__31704));
    InMux I__5675 (
            .O(N__31750),
            .I(N__31704));
    InMux I__5674 (
            .O(N__31749),
            .I(N__31704));
    InMux I__5673 (
            .O(N__31748),
            .I(N__31704));
    InMux I__5672 (
            .O(N__31747),
            .I(N__31704));
    InMux I__5671 (
            .O(N__31746),
            .I(N__31689));
    InMux I__5670 (
            .O(N__31745),
            .I(N__31689));
    InMux I__5669 (
            .O(N__31744),
            .I(N__31689));
    InMux I__5668 (
            .O(N__31743),
            .I(N__31689));
    InMux I__5667 (
            .O(N__31742),
            .I(N__31689));
    InMux I__5666 (
            .O(N__31741),
            .I(N__31689));
    InMux I__5665 (
            .O(N__31740),
            .I(N__31689));
    InMux I__5664 (
            .O(N__31739),
            .I(N__31678));
    InMux I__5663 (
            .O(N__31738),
            .I(N__31678));
    InMux I__5662 (
            .O(N__31737),
            .I(N__31678));
    InMux I__5661 (
            .O(N__31736),
            .I(N__31678));
    InMux I__5660 (
            .O(N__31735),
            .I(N__31678));
    InMux I__5659 (
            .O(N__31734),
            .I(N__31669));
    InMux I__5658 (
            .O(N__31733),
            .I(N__31669));
    InMux I__5657 (
            .O(N__31732),
            .I(N__31669));
    InMux I__5656 (
            .O(N__31731),
            .I(N__31669));
    LocalMux I__5655 (
            .O(N__31720),
            .I(N__31659));
    InMux I__5654 (
            .O(N__31719),
            .I(N__31648));
    InMux I__5653 (
            .O(N__31718),
            .I(N__31648));
    InMux I__5652 (
            .O(N__31717),
            .I(N__31648));
    InMux I__5651 (
            .O(N__31716),
            .I(N__31648));
    InMux I__5650 (
            .O(N__31715),
            .I(N__31648));
    LocalMux I__5649 (
            .O(N__31704),
            .I(N__31643));
    LocalMux I__5648 (
            .O(N__31689),
            .I(N__31643));
    LocalMux I__5647 (
            .O(N__31678),
            .I(N__31638));
    LocalMux I__5646 (
            .O(N__31669),
            .I(N__31638));
    InMux I__5645 (
            .O(N__31668),
            .I(N__31629));
    InMux I__5644 (
            .O(N__31667),
            .I(N__31629));
    InMux I__5643 (
            .O(N__31666),
            .I(N__31629));
    InMux I__5642 (
            .O(N__31665),
            .I(N__31629));
    InMux I__5641 (
            .O(N__31664),
            .I(N__31622));
    InMux I__5640 (
            .O(N__31663),
            .I(N__31622));
    InMux I__5639 (
            .O(N__31662),
            .I(N__31622));
    Odrv4 I__5638 (
            .O(N__31659),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt31_0 ));
    LocalMux I__5637 (
            .O(N__31648),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt31_0 ));
    Odrv4 I__5636 (
            .O(N__31643),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt31_0 ));
    Odrv4 I__5635 (
            .O(N__31638),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt31_0 ));
    LocalMux I__5634 (
            .O(N__31629),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt31_0 ));
    LocalMux I__5633 (
            .O(N__31622),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt31_0 ));
    CascadeMux I__5632 (
            .O(N__31609),
            .I(N__31606));
    InMux I__5631 (
            .O(N__31606),
            .I(N__31603));
    LocalMux I__5630 (
            .O(N__31603),
            .I(N__31600));
    Span4Mux_h I__5629 (
            .O(N__31600),
            .I(N__31597));
    Odrv4 I__5628 (
            .O(N__31597),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ));
    CEMux I__5627 (
            .O(N__31594),
            .I(N__31591));
    LocalMux I__5626 (
            .O(N__31591),
            .I(N__31588));
    Span4Mux_h I__5625 (
            .O(N__31588),
            .I(N__31585));
    Span4Mux_h I__5624 (
            .O(N__31585),
            .I(N__31579));
    CEMux I__5623 (
            .O(N__31584),
            .I(N__31576));
    CEMux I__5622 (
            .O(N__31583),
            .I(N__31573));
    CEMux I__5621 (
            .O(N__31582),
            .I(N__31570));
    Odrv4 I__5620 (
            .O(N__31579),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ));
    LocalMux I__5619 (
            .O(N__31576),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ));
    LocalMux I__5618 (
            .O(N__31573),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ));
    LocalMux I__5617 (
            .O(N__31570),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ));
    CascadeMux I__5616 (
            .O(N__31561),
            .I(N__31555));
    InMux I__5615 (
            .O(N__31560),
            .I(N__31552));
    InMux I__5614 (
            .O(N__31559),
            .I(N__31546));
    InMux I__5613 (
            .O(N__31558),
            .I(N__31546));
    InMux I__5612 (
            .O(N__31555),
            .I(N__31543));
    LocalMux I__5611 (
            .O(N__31552),
            .I(N__31540));
    InMux I__5610 (
            .O(N__31551),
            .I(N__31537));
    LocalMux I__5609 (
            .O(N__31546),
            .I(N__31534));
    LocalMux I__5608 (
            .O(N__31543),
            .I(measured_delay_hc_10));
    Odrv12 I__5607 (
            .O(N__31540),
            .I(measured_delay_hc_10));
    LocalMux I__5606 (
            .O(N__31537),
            .I(measured_delay_hc_10));
    Odrv4 I__5605 (
            .O(N__31534),
            .I(measured_delay_hc_10));
    CascadeMux I__5604 (
            .O(N__31525),
            .I(N__31517));
    CascadeMux I__5603 (
            .O(N__31524),
            .I(N__31514));
    CascadeMux I__5602 (
            .O(N__31523),
            .I(N__31503));
    CascadeMux I__5601 (
            .O(N__31522),
            .I(N__31494));
    CascadeMux I__5600 (
            .O(N__31521),
            .I(N__31489));
    CascadeMux I__5599 (
            .O(N__31520),
            .I(N__31486));
    InMux I__5598 (
            .O(N__31517),
            .I(N__31467));
    InMux I__5597 (
            .O(N__31514),
            .I(N__31467));
    InMux I__5596 (
            .O(N__31513),
            .I(N__31467));
    InMux I__5595 (
            .O(N__31512),
            .I(N__31467));
    InMux I__5594 (
            .O(N__31511),
            .I(N__31467));
    InMux I__5593 (
            .O(N__31510),
            .I(N__31456));
    InMux I__5592 (
            .O(N__31509),
            .I(N__31456));
    InMux I__5591 (
            .O(N__31508),
            .I(N__31456));
    InMux I__5590 (
            .O(N__31507),
            .I(N__31456));
    InMux I__5589 (
            .O(N__31506),
            .I(N__31456));
    InMux I__5588 (
            .O(N__31503),
            .I(N__31441));
    InMux I__5587 (
            .O(N__31502),
            .I(N__31441));
    InMux I__5586 (
            .O(N__31501),
            .I(N__31441));
    InMux I__5585 (
            .O(N__31500),
            .I(N__31441));
    InMux I__5584 (
            .O(N__31499),
            .I(N__31441));
    InMux I__5583 (
            .O(N__31498),
            .I(N__31441));
    InMux I__5582 (
            .O(N__31497),
            .I(N__31441));
    InMux I__5581 (
            .O(N__31494),
            .I(N__31437));
    InMux I__5580 (
            .O(N__31493),
            .I(N__31428));
    InMux I__5579 (
            .O(N__31492),
            .I(N__31428));
    InMux I__5578 (
            .O(N__31489),
            .I(N__31428));
    InMux I__5577 (
            .O(N__31486),
            .I(N__31428));
    InMux I__5576 (
            .O(N__31485),
            .I(N__31421));
    InMux I__5575 (
            .O(N__31484),
            .I(N__31421));
    InMux I__5574 (
            .O(N__31483),
            .I(N__31421));
    InMux I__5573 (
            .O(N__31482),
            .I(N__31410));
    InMux I__5572 (
            .O(N__31481),
            .I(N__31410));
    InMux I__5571 (
            .O(N__31480),
            .I(N__31410));
    InMux I__5570 (
            .O(N__31479),
            .I(N__31410));
    InMux I__5569 (
            .O(N__31478),
            .I(N__31410));
    LocalMux I__5568 (
            .O(N__31467),
            .I(N__31405));
    LocalMux I__5567 (
            .O(N__31456),
            .I(N__31405));
    LocalMux I__5566 (
            .O(N__31441),
            .I(N__31402));
    CascadeMux I__5565 (
            .O(N__31440),
            .I(N__31397));
    LocalMux I__5564 (
            .O(N__31437),
            .I(N__31384));
    LocalMux I__5563 (
            .O(N__31428),
            .I(N__31384));
    LocalMux I__5562 (
            .O(N__31421),
            .I(N__31379));
    LocalMux I__5561 (
            .O(N__31410),
            .I(N__31379));
    Span4Mux_v I__5560 (
            .O(N__31405),
            .I(N__31374));
    Span4Mux_v I__5559 (
            .O(N__31402),
            .I(N__31374));
    InMux I__5558 (
            .O(N__31401),
            .I(N__31371));
    InMux I__5557 (
            .O(N__31400),
            .I(N__31358));
    InMux I__5556 (
            .O(N__31397),
            .I(N__31358));
    InMux I__5555 (
            .O(N__31396),
            .I(N__31358));
    InMux I__5554 (
            .O(N__31395),
            .I(N__31358));
    InMux I__5553 (
            .O(N__31394),
            .I(N__31358));
    InMux I__5552 (
            .O(N__31393),
            .I(N__31358));
    InMux I__5551 (
            .O(N__31392),
            .I(N__31349));
    InMux I__5550 (
            .O(N__31391),
            .I(N__31349));
    InMux I__5549 (
            .O(N__31390),
            .I(N__31349));
    InMux I__5548 (
            .O(N__31389),
            .I(N__31349));
    Span4Mux_v I__5547 (
            .O(N__31384),
            .I(N__31346));
    Span4Mux_v I__5546 (
            .O(N__31379),
            .I(N__31343));
    Sp12to4 I__5545 (
            .O(N__31374),
            .I(N__31340));
    LocalMux I__5544 (
            .O(N__31371),
            .I(measured_delay_hc_31));
    LocalMux I__5543 (
            .O(N__31358),
            .I(measured_delay_hc_31));
    LocalMux I__5542 (
            .O(N__31349),
            .I(measured_delay_hc_31));
    Odrv4 I__5541 (
            .O(N__31346),
            .I(measured_delay_hc_31));
    Odrv4 I__5540 (
            .O(N__31343),
            .I(measured_delay_hc_31));
    Odrv12 I__5539 (
            .O(N__31340),
            .I(measured_delay_hc_31));
    InMux I__5538 (
            .O(N__31327),
            .I(N__31322));
    InMux I__5537 (
            .O(N__31326),
            .I(N__31319));
    InMux I__5536 (
            .O(N__31325),
            .I(N__31314));
    LocalMux I__5535 (
            .O(N__31322),
            .I(N__31311));
    LocalMux I__5534 (
            .O(N__31319),
            .I(N__31308));
    InMux I__5533 (
            .O(N__31318),
            .I(N__31305));
    InMux I__5532 (
            .O(N__31317),
            .I(N__31302));
    LocalMux I__5531 (
            .O(N__31314),
            .I(N__31299));
    Span4Mux_v I__5530 (
            .O(N__31311),
            .I(N__31294));
    Span4Mux_h I__5529 (
            .O(N__31308),
            .I(N__31294));
    LocalMux I__5528 (
            .O(N__31305),
            .I(N__31291));
    LocalMux I__5527 (
            .O(N__31302),
            .I(measured_delay_hc_3));
    Odrv4 I__5526 (
            .O(N__31299),
            .I(measured_delay_hc_3));
    Odrv4 I__5525 (
            .O(N__31294),
            .I(measured_delay_hc_3));
    Odrv12 I__5524 (
            .O(N__31291),
            .I(measured_delay_hc_3));
    CascadeMux I__5523 (
            .O(N__31282),
            .I(N__31275));
    InMux I__5522 (
            .O(N__31281),
            .I(N__31272));
    InMux I__5521 (
            .O(N__31280),
            .I(N__31269));
    InMux I__5520 (
            .O(N__31279),
            .I(N__31264));
    InMux I__5519 (
            .O(N__31278),
            .I(N__31264));
    InMux I__5518 (
            .O(N__31275),
            .I(N__31261));
    LocalMux I__5517 (
            .O(N__31272),
            .I(N__31258));
    LocalMux I__5516 (
            .O(N__31269),
            .I(N__31253));
    LocalMux I__5515 (
            .O(N__31264),
            .I(N__31253));
    LocalMux I__5514 (
            .O(N__31261),
            .I(measured_delay_hc_12));
    Odrv12 I__5513 (
            .O(N__31258),
            .I(measured_delay_hc_12));
    Odrv4 I__5512 (
            .O(N__31253),
            .I(measured_delay_hc_12));
    InMux I__5511 (
            .O(N__31246),
            .I(N__31241));
    CascadeMux I__5510 (
            .O(N__31245),
            .I(N__31236));
    InMux I__5509 (
            .O(N__31244),
            .I(N__31233));
    LocalMux I__5508 (
            .O(N__31241),
            .I(N__31230));
    InMux I__5507 (
            .O(N__31240),
            .I(N__31225));
    InMux I__5506 (
            .O(N__31239),
            .I(N__31225));
    InMux I__5505 (
            .O(N__31236),
            .I(N__31222));
    LocalMux I__5504 (
            .O(N__31233),
            .I(N__31219));
    Span4Mux_h I__5503 (
            .O(N__31230),
            .I(N__31216));
    LocalMux I__5502 (
            .O(N__31225),
            .I(N__31213));
    LocalMux I__5501 (
            .O(N__31222),
            .I(measured_delay_hc_18));
    Odrv4 I__5500 (
            .O(N__31219),
            .I(measured_delay_hc_18));
    Odrv4 I__5499 (
            .O(N__31216),
            .I(measured_delay_hc_18));
    Odrv12 I__5498 (
            .O(N__31213),
            .I(measured_delay_hc_18));
    InMux I__5497 (
            .O(N__31204),
            .I(N__31198));
    InMux I__5496 (
            .O(N__31203),
            .I(N__31192));
    InMux I__5495 (
            .O(N__31202),
            .I(N__31192));
    CascadeMux I__5494 (
            .O(N__31201),
            .I(N__31189));
    LocalMux I__5493 (
            .O(N__31198),
            .I(N__31186));
    InMux I__5492 (
            .O(N__31197),
            .I(N__31183));
    LocalMux I__5491 (
            .O(N__31192),
            .I(N__31180));
    InMux I__5490 (
            .O(N__31189),
            .I(N__31177));
    Span4Mux_v I__5489 (
            .O(N__31186),
            .I(N__31170));
    LocalMux I__5488 (
            .O(N__31183),
            .I(N__31170));
    Span4Mux_h I__5487 (
            .O(N__31180),
            .I(N__31170));
    LocalMux I__5486 (
            .O(N__31177),
            .I(measured_delay_hc_17));
    Odrv4 I__5485 (
            .O(N__31170),
            .I(measured_delay_hc_17));
    InMux I__5484 (
            .O(N__31165),
            .I(N__31160));
    InMux I__5483 (
            .O(N__31164),
            .I(N__31157));
    CascadeMux I__5482 (
            .O(N__31163),
            .I(N__31153));
    LocalMux I__5481 (
            .O(N__31160),
            .I(N__31147));
    LocalMux I__5480 (
            .O(N__31157),
            .I(N__31147));
    InMux I__5479 (
            .O(N__31156),
            .I(N__31144));
    InMux I__5478 (
            .O(N__31153),
            .I(N__31141));
    InMux I__5477 (
            .O(N__31152),
            .I(N__31138));
    Span4Mux_h I__5476 (
            .O(N__31147),
            .I(N__31135));
    LocalMux I__5475 (
            .O(N__31144),
            .I(N__31130));
    LocalMux I__5474 (
            .O(N__31141),
            .I(N__31130));
    LocalMux I__5473 (
            .O(N__31138),
            .I(measured_delay_hc_5));
    Odrv4 I__5472 (
            .O(N__31135),
            .I(measured_delay_hc_5));
    Odrv12 I__5471 (
            .O(N__31130),
            .I(measured_delay_hc_5));
    CascadeMux I__5470 (
            .O(N__31123),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt9_0_cascade_ ));
    InMux I__5469 (
            .O(N__31120),
            .I(N__31117));
    LocalMux I__5468 (
            .O(N__31117),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt15 ));
    InMux I__5467 (
            .O(N__31114),
            .I(N__31111));
    LocalMux I__5466 (
            .O(N__31111),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto13Z0Z_1 ));
    CascadeMux I__5465 (
            .O(N__31108),
            .I(N__31090));
    CascadeMux I__5464 (
            .O(N__31107),
            .I(N__31087));
    CascadeMux I__5463 (
            .O(N__31106),
            .I(N__31084));
    CascadeMux I__5462 (
            .O(N__31105),
            .I(N__31081));
    CascadeMux I__5461 (
            .O(N__31104),
            .I(N__31074));
    CascadeMux I__5460 (
            .O(N__31103),
            .I(N__31071));
    CascadeMux I__5459 (
            .O(N__31102),
            .I(N__31068));
    CascadeMux I__5458 (
            .O(N__31101),
            .I(N__31065));
    CascadeMux I__5457 (
            .O(N__31100),
            .I(N__31062));
    CascadeMux I__5456 (
            .O(N__31099),
            .I(N__31059));
    CascadeMux I__5455 (
            .O(N__31098),
            .I(N__31056));
    CascadeMux I__5454 (
            .O(N__31097),
            .I(N__31053));
    CascadeMux I__5453 (
            .O(N__31096),
            .I(N__31050));
    CascadeMux I__5452 (
            .O(N__31095),
            .I(N__31047));
    CascadeMux I__5451 (
            .O(N__31094),
            .I(N__31044));
    InMux I__5450 (
            .O(N__31093),
            .I(N__31027));
    InMux I__5449 (
            .O(N__31090),
            .I(N__31027));
    InMux I__5448 (
            .O(N__31087),
            .I(N__31027));
    InMux I__5447 (
            .O(N__31084),
            .I(N__31027));
    InMux I__5446 (
            .O(N__31081),
            .I(N__31027));
    InMux I__5445 (
            .O(N__31080),
            .I(N__31027));
    InMux I__5444 (
            .O(N__31079),
            .I(N__31027));
    InMux I__5443 (
            .O(N__31078),
            .I(N__31027));
    CascadeMux I__5442 (
            .O(N__31077),
            .I(N__31023));
    InMux I__5441 (
            .O(N__31074),
            .I(N__31013));
    InMux I__5440 (
            .O(N__31071),
            .I(N__31013));
    InMux I__5439 (
            .O(N__31068),
            .I(N__31013));
    InMux I__5438 (
            .O(N__31065),
            .I(N__31013));
    InMux I__5437 (
            .O(N__31062),
            .I(N__31004));
    InMux I__5436 (
            .O(N__31059),
            .I(N__31004));
    InMux I__5435 (
            .O(N__31056),
            .I(N__31004));
    InMux I__5434 (
            .O(N__31053),
            .I(N__31004));
    InMux I__5433 (
            .O(N__31050),
            .I(N__30999));
    InMux I__5432 (
            .O(N__31047),
            .I(N__30999));
    InMux I__5431 (
            .O(N__31044),
            .I(N__30996));
    LocalMux I__5430 (
            .O(N__31027),
            .I(N__30993));
    InMux I__5429 (
            .O(N__31026),
            .I(N__30990));
    InMux I__5428 (
            .O(N__31023),
            .I(N__30984));
    InMux I__5427 (
            .O(N__31022),
            .I(N__30984));
    LocalMux I__5426 (
            .O(N__31013),
            .I(N__30979));
    LocalMux I__5425 (
            .O(N__31004),
            .I(N__30979));
    LocalMux I__5424 (
            .O(N__30999),
            .I(N__30976));
    LocalMux I__5423 (
            .O(N__30996),
            .I(N__30973));
    Span4Mux_h I__5422 (
            .O(N__30993),
            .I(N__30967));
    LocalMux I__5421 (
            .O(N__30990),
            .I(N__30967));
    CascadeMux I__5420 (
            .O(N__30989),
            .I(N__30964));
    LocalMux I__5419 (
            .O(N__30984),
            .I(N__30959));
    Span4Mux_v I__5418 (
            .O(N__30979),
            .I(N__30959));
    Span4Mux_h I__5417 (
            .O(N__30976),
            .I(N__30954));
    Span4Mux_h I__5416 (
            .O(N__30973),
            .I(N__30954));
    InMux I__5415 (
            .O(N__30972),
            .I(N__30951));
    Span4Mux_v I__5414 (
            .O(N__30967),
            .I(N__30948));
    InMux I__5413 (
            .O(N__30964),
            .I(N__30945));
    Span4Mux_v I__5412 (
            .O(N__30959),
            .I(N__30942));
    Sp12to4 I__5411 (
            .O(N__30954),
            .I(N__30937));
    LocalMux I__5410 (
            .O(N__30951),
            .I(N__30937));
    Span4Mux_h I__5409 (
            .O(N__30948),
            .I(N__30934));
    LocalMux I__5408 (
            .O(N__30945),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__5407 (
            .O(N__30942),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv12 I__5406 (
            .O(N__30937),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__5405 (
            .O(N__30934),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    CascadeMux I__5404 (
            .O(N__30925),
            .I(N__30919));
    CascadeMux I__5403 (
            .O(N__30924),
            .I(N__30916));
    CascadeMux I__5402 (
            .O(N__30923),
            .I(N__30913));
    CascadeMux I__5401 (
            .O(N__30922),
            .I(N__30910));
    InMux I__5400 (
            .O(N__30919),
            .I(N__30883));
    InMux I__5399 (
            .O(N__30916),
            .I(N__30883));
    InMux I__5398 (
            .O(N__30913),
            .I(N__30883));
    InMux I__5397 (
            .O(N__30910),
            .I(N__30883));
    InMux I__5396 (
            .O(N__30909),
            .I(N__30880));
    InMux I__5395 (
            .O(N__30908),
            .I(N__30863));
    InMux I__5394 (
            .O(N__30907),
            .I(N__30863));
    InMux I__5393 (
            .O(N__30906),
            .I(N__30863));
    InMux I__5392 (
            .O(N__30905),
            .I(N__30863));
    InMux I__5391 (
            .O(N__30904),
            .I(N__30863));
    InMux I__5390 (
            .O(N__30903),
            .I(N__30863));
    InMux I__5389 (
            .O(N__30902),
            .I(N__30863));
    InMux I__5388 (
            .O(N__30901),
            .I(N__30863));
    InMux I__5387 (
            .O(N__30900),
            .I(N__30854));
    InMux I__5386 (
            .O(N__30899),
            .I(N__30854));
    InMux I__5385 (
            .O(N__30898),
            .I(N__30854));
    InMux I__5384 (
            .O(N__30897),
            .I(N__30854));
    InMux I__5383 (
            .O(N__30896),
            .I(N__30851));
    InMux I__5382 (
            .O(N__30895),
            .I(N__30848));
    InMux I__5381 (
            .O(N__30894),
            .I(N__30845));
    InMux I__5380 (
            .O(N__30893),
            .I(N__30838));
    InMux I__5379 (
            .O(N__30892),
            .I(N__30838));
    LocalMux I__5378 (
            .O(N__30883),
            .I(N__30829));
    LocalMux I__5377 (
            .O(N__30880),
            .I(N__30829));
    LocalMux I__5376 (
            .O(N__30863),
            .I(N__30829));
    LocalMux I__5375 (
            .O(N__30854),
            .I(N__30829));
    LocalMux I__5374 (
            .O(N__30851),
            .I(N__30826));
    LocalMux I__5373 (
            .O(N__30848),
            .I(N__30821));
    LocalMux I__5372 (
            .O(N__30845),
            .I(N__30821));
    InMux I__5371 (
            .O(N__30844),
            .I(N__30816));
    InMux I__5370 (
            .O(N__30843),
            .I(N__30816));
    LocalMux I__5369 (
            .O(N__30838),
            .I(N__30811));
    Span4Mux_v I__5368 (
            .O(N__30829),
            .I(N__30811));
    Span4Mux_v I__5367 (
            .O(N__30826),
            .I(N__30806));
    Span4Mux_v I__5366 (
            .O(N__30821),
            .I(N__30806));
    LocalMux I__5365 (
            .O(N__30816),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__5364 (
            .O(N__30811),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__5363 (
            .O(N__30806),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    InMux I__5362 (
            .O(N__30799),
            .I(N__30788));
    InMux I__5361 (
            .O(N__30798),
            .I(N__30771));
    InMux I__5360 (
            .O(N__30797),
            .I(N__30771));
    InMux I__5359 (
            .O(N__30796),
            .I(N__30771));
    InMux I__5358 (
            .O(N__30795),
            .I(N__30771));
    InMux I__5357 (
            .O(N__30794),
            .I(N__30771));
    InMux I__5356 (
            .O(N__30793),
            .I(N__30771));
    InMux I__5355 (
            .O(N__30792),
            .I(N__30771));
    InMux I__5354 (
            .O(N__30791),
            .I(N__30771));
    LocalMux I__5353 (
            .O(N__30788),
            .I(N__30752));
    LocalMux I__5352 (
            .O(N__30771),
            .I(N__30752));
    InMux I__5351 (
            .O(N__30770),
            .I(N__30749));
    InMux I__5350 (
            .O(N__30769),
            .I(N__30746));
    InMux I__5349 (
            .O(N__30768),
            .I(N__30741));
    InMux I__5348 (
            .O(N__30767),
            .I(N__30741));
    InMux I__5347 (
            .O(N__30766),
            .I(N__30724));
    InMux I__5346 (
            .O(N__30765),
            .I(N__30724));
    InMux I__5345 (
            .O(N__30764),
            .I(N__30724));
    InMux I__5344 (
            .O(N__30763),
            .I(N__30724));
    InMux I__5343 (
            .O(N__30762),
            .I(N__30724));
    InMux I__5342 (
            .O(N__30761),
            .I(N__30724));
    InMux I__5341 (
            .O(N__30760),
            .I(N__30724));
    InMux I__5340 (
            .O(N__30759),
            .I(N__30724));
    InMux I__5339 (
            .O(N__30758),
            .I(N__30721));
    CascadeMux I__5338 (
            .O(N__30757),
            .I(N__30718));
    Span4Mux_v I__5337 (
            .O(N__30752),
            .I(N__30712));
    LocalMux I__5336 (
            .O(N__30749),
            .I(N__30712));
    LocalMux I__5335 (
            .O(N__30746),
            .I(N__30709));
    LocalMux I__5334 (
            .O(N__30741),
            .I(N__30702));
    LocalMux I__5333 (
            .O(N__30724),
            .I(N__30702));
    LocalMux I__5332 (
            .O(N__30721),
            .I(N__30702));
    InMux I__5331 (
            .O(N__30718),
            .I(N__30697));
    InMux I__5330 (
            .O(N__30717),
            .I(N__30697));
    Span4Mux_v I__5329 (
            .O(N__30712),
            .I(N__30692));
    Span4Mux_v I__5328 (
            .O(N__30709),
            .I(N__30692));
    Span4Mux_v I__5327 (
            .O(N__30702),
            .I(N__30689));
    LocalMux I__5326 (
            .O(N__30697),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__5325 (
            .O(N__30692),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__5324 (
            .O(N__30689),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    InMux I__5323 (
            .O(N__30682),
            .I(N__30678));
    InMux I__5322 (
            .O(N__30681),
            .I(N__30675));
    LocalMux I__5321 (
            .O(N__30678),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto8Z0Z_0 ));
    LocalMux I__5320 (
            .O(N__30675),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto8Z0Z_0 ));
    InMux I__5319 (
            .O(N__30670),
            .I(N__30667));
    LocalMux I__5318 (
            .O(N__30667),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9 ));
    CascadeMux I__5317 (
            .O(N__30664),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6_cascade_ ));
    InMux I__5316 (
            .O(N__30661),
            .I(N__30658));
    LocalMux I__5315 (
            .O(N__30658),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_12 ));
    CascadeMux I__5314 (
            .O(N__30655),
            .I(N__30652));
    InMux I__5313 (
            .O(N__30652),
            .I(N__30649));
    LocalMux I__5312 (
            .O(N__30649),
            .I(N__30646));
    Span4Mux_h I__5311 (
            .O(N__30646),
            .I(N__30643));
    Odrv4 I__5310 (
            .O(N__30643),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ));
    CascadeMux I__5309 (
            .O(N__30640),
            .I(N__30637));
    InMux I__5308 (
            .O(N__30637),
            .I(N__30634));
    LocalMux I__5307 (
            .O(N__30634),
            .I(N__30631));
    Odrv4 I__5306 (
            .O(N__30631),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ));
    CascadeMux I__5305 (
            .O(N__30628),
            .I(N__30625));
    InMux I__5304 (
            .O(N__30625),
            .I(N__30622));
    LocalMux I__5303 (
            .O(N__30622),
            .I(N__30619));
    Span4Mux_h I__5302 (
            .O(N__30619),
            .I(N__30616));
    Odrv4 I__5301 (
            .O(N__30616),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ));
    CEMux I__5300 (
            .O(N__30613),
            .I(N__30608));
    CEMux I__5299 (
            .O(N__30612),
            .I(N__30605));
    CEMux I__5298 (
            .O(N__30611),
            .I(N__30602));
    LocalMux I__5297 (
            .O(N__30608),
            .I(N__30599));
    LocalMux I__5296 (
            .O(N__30605),
            .I(N__30596));
    LocalMux I__5295 (
            .O(N__30602),
            .I(N__30592));
    Span4Mux_h I__5294 (
            .O(N__30599),
            .I(N__30589));
    Span4Mux_h I__5293 (
            .O(N__30596),
            .I(N__30586));
    CEMux I__5292 (
            .O(N__30595),
            .I(N__30583));
    Span4Mux_v I__5291 (
            .O(N__30592),
            .I(N__30580));
    Span4Mux_h I__5290 (
            .O(N__30589),
            .I(N__30577));
    Span4Mux_h I__5289 (
            .O(N__30586),
            .I(N__30574));
    LocalMux I__5288 (
            .O(N__30583),
            .I(N__30571));
    Odrv4 I__5287 (
            .O(N__30580),
            .I(\phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa ));
    Odrv4 I__5286 (
            .O(N__30577),
            .I(\phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa ));
    Odrv4 I__5285 (
            .O(N__30574),
            .I(\phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa ));
    Odrv12 I__5284 (
            .O(N__30571),
            .I(\phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa ));
    CascadeMux I__5283 (
            .O(N__30562),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2_cascade_ ));
    CascadeMux I__5282 (
            .O(N__30559),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7_cascade_ ));
    CascadeMux I__5281 (
            .O(N__30556),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_11_cascade_ ));
    CascadeMux I__5280 (
            .O(N__30553),
            .I(N__30546));
    InMux I__5279 (
            .O(N__30552),
            .I(N__30540));
    InMux I__5278 (
            .O(N__30551),
            .I(N__30533));
    InMux I__5277 (
            .O(N__30550),
            .I(N__30533));
    InMux I__5276 (
            .O(N__30549),
            .I(N__30533));
    InMux I__5275 (
            .O(N__30546),
            .I(N__30530));
    InMux I__5274 (
            .O(N__30545),
            .I(N__30523));
    InMux I__5273 (
            .O(N__30544),
            .I(N__30523));
    InMux I__5272 (
            .O(N__30543),
            .I(N__30523));
    LocalMux I__5271 (
            .O(N__30540),
            .I(N__30520));
    LocalMux I__5270 (
            .O(N__30533),
            .I(N__30517));
    LocalMux I__5269 (
            .O(N__30530),
            .I(\phase_controller_inst1.stoper_hc.un2_startlt31 ));
    LocalMux I__5268 (
            .O(N__30523),
            .I(\phase_controller_inst1.stoper_hc.un2_startlt31 ));
    Odrv4 I__5267 (
            .O(N__30520),
            .I(\phase_controller_inst1.stoper_hc.un2_startlt31 ));
    Odrv12 I__5266 (
            .O(N__30517),
            .I(\phase_controller_inst1.stoper_hc.un2_startlt31 ));
    InMux I__5265 (
            .O(N__30508),
            .I(N__30505));
    LocalMux I__5264 (
            .O(N__30505),
            .I(N__30502));
    Span4Mux_h I__5263 (
            .O(N__30502),
            .I(N__30499));
    Span4Mux_v I__5262 (
            .O(N__30499),
            .I(N__30493));
    InMux I__5261 (
            .O(N__30498),
            .I(N__30490));
    InMux I__5260 (
            .O(N__30497),
            .I(N__30487));
    InMux I__5259 (
            .O(N__30496),
            .I(N__30484));
    Span4Mux_v I__5258 (
            .O(N__30493),
            .I(N__30481));
    LocalMux I__5257 (
            .O(N__30490),
            .I(N__30478));
    LocalMux I__5256 (
            .O(N__30487),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    LocalMux I__5255 (
            .O(N__30484),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    Odrv4 I__5254 (
            .O(N__30481),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    Odrv4 I__5253 (
            .O(N__30478),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    InMux I__5252 (
            .O(N__30469),
            .I(N__30466));
    LocalMux I__5251 (
            .O(N__30466),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto5Z0Z_3 ));
    CascadeMux I__5250 (
            .O(N__30463),
            .I(N__30460));
    InMux I__5249 (
            .O(N__30460),
            .I(N__30457));
    LocalMux I__5248 (
            .O(N__30457),
            .I(N__30454));
    Span4Mux_h I__5247 (
            .O(N__30454),
            .I(N__30451));
    Odrv4 I__5246 (
            .O(N__30451),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ));
    InMux I__5245 (
            .O(N__30448),
            .I(N__30430));
    InMux I__5244 (
            .O(N__30447),
            .I(N__30430));
    InMux I__5243 (
            .O(N__30446),
            .I(N__30405));
    InMux I__5242 (
            .O(N__30445),
            .I(N__30405));
    InMux I__5241 (
            .O(N__30444),
            .I(N__30405));
    InMux I__5240 (
            .O(N__30443),
            .I(N__30405));
    InMux I__5239 (
            .O(N__30442),
            .I(N__30405));
    InMux I__5238 (
            .O(N__30441),
            .I(N__30405));
    InMux I__5237 (
            .O(N__30440),
            .I(N__30405));
    InMux I__5236 (
            .O(N__30439),
            .I(N__30405));
    InMux I__5235 (
            .O(N__30438),
            .I(N__30402));
    InMux I__5234 (
            .O(N__30437),
            .I(N__30397));
    InMux I__5233 (
            .O(N__30436),
            .I(N__30397));
    InMux I__5232 (
            .O(N__30435),
            .I(N__30394));
    LocalMux I__5231 (
            .O(N__30430),
            .I(N__30391));
    InMux I__5230 (
            .O(N__30429),
            .I(N__30372));
    InMux I__5229 (
            .O(N__30428),
            .I(N__30372));
    InMux I__5228 (
            .O(N__30427),
            .I(N__30372));
    InMux I__5227 (
            .O(N__30426),
            .I(N__30372));
    InMux I__5226 (
            .O(N__30425),
            .I(N__30372));
    InMux I__5225 (
            .O(N__30424),
            .I(N__30372));
    InMux I__5224 (
            .O(N__30423),
            .I(N__30372));
    InMux I__5223 (
            .O(N__30422),
            .I(N__30372));
    LocalMux I__5222 (
            .O(N__30405),
            .I(N__30369));
    LocalMux I__5221 (
            .O(N__30402),
            .I(N__30366));
    LocalMux I__5220 (
            .O(N__30397),
            .I(N__30361));
    LocalMux I__5219 (
            .O(N__30394),
            .I(N__30361));
    Span4Mux_v I__5218 (
            .O(N__30391),
            .I(N__30358));
    InMux I__5217 (
            .O(N__30390),
            .I(N__30353));
    InMux I__5216 (
            .O(N__30389),
            .I(N__30353));
    LocalMux I__5215 (
            .O(N__30372),
            .I(N__30346));
    Span4Mux_h I__5214 (
            .O(N__30369),
            .I(N__30346));
    Span4Mux_h I__5213 (
            .O(N__30366),
            .I(N__30346));
    Sp12to4 I__5212 (
            .O(N__30361),
            .I(N__30343));
    Span4Mux_h I__5211 (
            .O(N__30358),
            .I(N__30340));
    LocalMux I__5210 (
            .O(N__30353),
            .I(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__5209 (
            .O(N__30346),
            .I(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv12 I__5208 (
            .O(N__30343),
            .I(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__5207 (
            .O(N__30340),
            .I(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0 ));
    CascadeMux I__5206 (
            .O(N__30331),
            .I(N__30328));
    InMux I__5205 (
            .O(N__30328),
            .I(N__30310));
    InMux I__5204 (
            .O(N__30327),
            .I(N__30310));
    CascadeMux I__5203 (
            .O(N__30326),
            .I(N__30304));
    CascadeMux I__5202 (
            .O(N__30325),
            .I(N__30301));
    CascadeMux I__5201 (
            .O(N__30324),
            .I(N__30298));
    CascadeMux I__5200 (
            .O(N__30323),
            .I(N__30295));
    InMux I__5199 (
            .O(N__30322),
            .I(N__30274));
    InMux I__5198 (
            .O(N__30321),
            .I(N__30274));
    InMux I__5197 (
            .O(N__30320),
            .I(N__30274));
    InMux I__5196 (
            .O(N__30319),
            .I(N__30274));
    InMux I__5195 (
            .O(N__30318),
            .I(N__30274));
    InMux I__5194 (
            .O(N__30317),
            .I(N__30274));
    InMux I__5193 (
            .O(N__30316),
            .I(N__30274));
    InMux I__5192 (
            .O(N__30315),
            .I(N__30274));
    LocalMux I__5191 (
            .O(N__30310),
            .I(N__30271));
    InMux I__5190 (
            .O(N__30309),
            .I(N__30268));
    CascadeMux I__5189 (
            .O(N__30308),
            .I(N__30265));
    CascadeMux I__5188 (
            .O(N__30307),
            .I(N__30262));
    InMux I__5187 (
            .O(N__30304),
            .I(N__30243));
    InMux I__5186 (
            .O(N__30301),
            .I(N__30243));
    InMux I__5185 (
            .O(N__30298),
            .I(N__30243));
    InMux I__5184 (
            .O(N__30295),
            .I(N__30243));
    InMux I__5183 (
            .O(N__30294),
            .I(N__30243));
    InMux I__5182 (
            .O(N__30293),
            .I(N__30243));
    InMux I__5181 (
            .O(N__30292),
            .I(N__30243));
    InMux I__5180 (
            .O(N__30291),
            .I(N__30243));
    LocalMux I__5179 (
            .O(N__30274),
            .I(N__30240));
    Span4Mux_v I__5178 (
            .O(N__30271),
            .I(N__30234));
    LocalMux I__5177 (
            .O(N__30268),
            .I(N__30234));
    InMux I__5176 (
            .O(N__30265),
            .I(N__30229));
    InMux I__5175 (
            .O(N__30262),
            .I(N__30229));
    InMux I__5174 (
            .O(N__30261),
            .I(N__30224));
    InMux I__5173 (
            .O(N__30260),
            .I(N__30224));
    LocalMux I__5172 (
            .O(N__30243),
            .I(N__30221));
    Span4Mux_v I__5171 (
            .O(N__30240),
            .I(N__30218));
    InMux I__5170 (
            .O(N__30239),
            .I(N__30215));
    Span4Mux_h I__5169 (
            .O(N__30234),
            .I(N__30212));
    LocalMux I__5168 (
            .O(N__30229),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    LocalMux I__5167 (
            .O(N__30224),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    Odrv4 I__5166 (
            .O(N__30221),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    Odrv4 I__5165 (
            .O(N__30218),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    LocalMux I__5164 (
            .O(N__30215),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    Odrv4 I__5163 (
            .O(N__30212),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    CascadeMux I__5162 (
            .O(N__30199),
            .I(N__30176));
    CascadeMux I__5161 (
            .O(N__30198),
            .I(N__30173));
    CascadeMux I__5160 (
            .O(N__30197),
            .I(N__30170));
    CascadeMux I__5159 (
            .O(N__30196),
            .I(N__30167));
    InMux I__5158 (
            .O(N__30195),
            .I(N__30149));
    InMux I__5157 (
            .O(N__30194),
            .I(N__30149));
    InMux I__5156 (
            .O(N__30193),
            .I(N__30149));
    InMux I__5155 (
            .O(N__30192),
            .I(N__30149));
    InMux I__5154 (
            .O(N__30191),
            .I(N__30149));
    InMux I__5153 (
            .O(N__30190),
            .I(N__30149));
    InMux I__5152 (
            .O(N__30189),
            .I(N__30149));
    InMux I__5151 (
            .O(N__30188),
            .I(N__30149));
    InMux I__5150 (
            .O(N__30187),
            .I(N__30143));
    InMux I__5149 (
            .O(N__30186),
            .I(N__30143));
    CascadeMux I__5148 (
            .O(N__30185),
            .I(N__30140));
    InMux I__5147 (
            .O(N__30184),
            .I(N__30134));
    InMux I__5146 (
            .O(N__30183),
            .I(N__30134));
    InMux I__5145 (
            .O(N__30182),
            .I(N__30117));
    InMux I__5144 (
            .O(N__30181),
            .I(N__30117));
    InMux I__5143 (
            .O(N__30180),
            .I(N__30117));
    InMux I__5142 (
            .O(N__30179),
            .I(N__30117));
    InMux I__5141 (
            .O(N__30176),
            .I(N__30117));
    InMux I__5140 (
            .O(N__30173),
            .I(N__30117));
    InMux I__5139 (
            .O(N__30170),
            .I(N__30117));
    InMux I__5138 (
            .O(N__30167),
            .I(N__30117));
    InMux I__5137 (
            .O(N__30166),
            .I(N__30114));
    LocalMux I__5136 (
            .O(N__30149),
            .I(N__30111));
    InMux I__5135 (
            .O(N__30148),
            .I(N__30108));
    LocalMux I__5134 (
            .O(N__30143),
            .I(N__30105));
    InMux I__5133 (
            .O(N__30140),
            .I(N__30100));
    InMux I__5132 (
            .O(N__30139),
            .I(N__30100));
    LocalMux I__5131 (
            .O(N__30134),
            .I(N__30097));
    LocalMux I__5130 (
            .O(N__30117),
            .I(N__30092));
    LocalMux I__5129 (
            .O(N__30114),
            .I(N__30092));
    Span4Mux_v I__5128 (
            .O(N__30111),
            .I(N__30085));
    LocalMux I__5127 (
            .O(N__30108),
            .I(N__30085));
    Span4Mux_v I__5126 (
            .O(N__30105),
            .I(N__30085));
    LocalMux I__5125 (
            .O(N__30100),
            .I(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv12 I__5124 (
            .O(N__30097),
            .I(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__5123 (
            .O(N__30092),
            .I(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__5122 (
            .O(N__30085),
            .I(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1 ));
    InMux I__5121 (
            .O(N__30076),
            .I(N__30072));
    InMux I__5120 (
            .O(N__30075),
            .I(N__30069));
    LocalMux I__5119 (
            .O(N__30072),
            .I(N__30066));
    LocalMux I__5118 (
            .O(N__30069),
            .I(N__30062));
    Span12Mux_h I__5117 (
            .O(N__30066),
            .I(N__30058));
    InMux I__5116 (
            .O(N__30065),
            .I(N__30055));
    Span4Mux_v I__5115 (
            .O(N__30062),
            .I(N__30052));
    InMux I__5114 (
            .O(N__30061),
            .I(N__30049));
    Odrv12 I__5113 (
            .O(N__30058),
            .I(\phase_controller_inst2.stoper_hc.time_passed11 ));
    LocalMux I__5112 (
            .O(N__30055),
            .I(\phase_controller_inst2.stoper_hc.time_passed11 ));
    Odrv4 I__5111 (
            .O(N__30052),
            .I(\phase_controller_inst2.stoper_hc.time_passed11 ));
    LocalMux I__5110 (
            .O(N__30049),
            .I(\phase_controller_inst2.stoper_hc.time_passed11 ));
    InMux I__5109 (
            .O(N__30040),
            .I(N__30037));
    LocalMux I__5108 (
            .O(N__30037),
            .I(N__30034));
    Span4Mux_v I__5107 (
            .O(N__30034),
            .I(N__30028));
    InMux I__5106 (
            .O(N__30033),
            .I(N__30021));
    InMux I__5105 (
            .O(N__30032),
            .I(N__30021));
    InMux I__5104 (
            .O(N__30031),
            .I(N__30021));
    Span4Mux_v I__5103 (
            .O(N__30028),
            .I(N__30016));
    LocalMux I__5102 (
            .O(N__30021),
            .I(N__30013));
    InMux I__5101 (
            .O(N__30020),
            .I(N__30008));
    InMux I__5100 (
            .O(N__30019),
            .I(N__30008));
    Odrv4 I__5099 (
            .O(N__30016),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__5098 (
            .O(N__30013),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__5097 (
            .O(N__30008),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    InMux I__5096 (
            .O(N__30001),
            .I(N__29998));
    LocalMux I__5095 (
            .O(N__29998),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIUO2PZ0 ));
    InMux I__5094 (
            .O(N__29995),
            .I(N__29984));
    InMux I__5093 (
            .O(N__29994),
            .I(N__29984));
    CascadeMux I__5092 (
            .O(N__29993),
            .I(N__29978));
    CascadeMux I__5091 (
            .O(N__29992),
            .I(N__29975));
    CascadeMux I__5090 (
            .O(N__29991),
            .I(N__29972));
    CascadeMux I__5089 (
            .O(N__29990),
            .I(N__29969));
    CascadeMux I__5088 (
            .O(N__29989),
            .I(N__29966));
    LocalMux I__5087 (
            .O(N__29984),
            .I(N__29960));
    InMux I__5086 (
            .O(N__29983),
            .I(N__29942));
    InMux I__5085 (
            .O(N__29982),
            .I(N__29942));
    InMux I__5084 (
            .O(N__29981),
            .I(N__29942));
    InMux I__5083 (
            .O(N__29978),
            .I(N__29942));
    InMux I__5082 (
            .O(N__29975),
            .I(N__29942));
    InMux I__5081 (
            .O(N__29972),
            .I(N__29942));
    InMux I__5080 (
            .O(N__29969),
            .I(N__29931));
    InMux I__5079 (
            .O(N__29966),
            .I(N__29931));
    InMux I__5078 (
            .O(N__29965),
            .I(N__29931));
    InMux I__5077 (
            .O(N__29964),
            .I(N__29931));
    InMux I__5076 (
            .O(N__29963),
            .I(N__29931));
    Span4Mux_v I__5075 (
            .O(N__29960),
            .I(N__29928));
    CascadeMux I__5074 (
            .O(N__29959),
            .I(N__29923));
    CascadeMux I__5073 (
            .O(N__29958),
            .I(N__29920));
    CascadeMux I__5072 (
            .O(N__29957),
            .I(N__29917));
    CascadeMux I__5071 (
            .O(N__29956),
            .I(N__29914));
    CascadeMux I__5070 (
            .O(N__29955),
            .I(N__29911));
    LocalMux I__5069 (
            .O(N__29942),
            .I(N__29900));
    LocalMux I__5068 (
            .O(N__29931),
            .I(N__29900));
    Span4Mux_h I__5067 (
            .O(N__29928),
            .I(N__29900));
    InMux I__5066 (
            .O(N__29927),
            .I(N__29895));
    InMux I__5065 (
            .O(N__29926),
            .I(N__29895));
    InMux I__5064 (
            .O(N__29923),
            .I(N__29892));
    InMux I__5063 (
            .O(N__29920),
            .I(N__29877));
    InMux I__5062 (
            .O(N__29917),
            .I(N__29877));
    InMux I__5061 (
            .O(N__29914),
            .I(N__29877));
    InMux I__5060 (
            .O(N__29911),
            .I(N__29877));
    InMux I__5059 (
            .O(N__29910),
            .I(N__29877));
    InMux I__5058 (
            .O(N__29909),
            .I(N__29877));
    InMux I__5057 (
            .O(N__29908),
            .I(N__29877));
    InMux I__5056 (
            .O(N__29907),
            .I(N__29874));
    Span4Mux_v I__5055 (
            .O(N__29900),
            .I(N__29869));
    LocalMux I__5054 (
            .O(N__29895),
            .I(N__29869));
    LocalMux I__5053 (
            .O(N__29892),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    LocalMux I__5052 (
            .O(N__29877),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    LocalMux I__5051 (
            .O(N__29874),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    Odrv4 I__5050 (
            .O(N__29869),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    InMux I__5049 (
            .O(N__29860),
            .I(N__29855));
    InMux I__5048 (
            .O(N__29859),
            .I(N__29852));
    InMux I__5047 (
            .O(N__29858),
            .I(N__29849));
    LocalMux I__5046 (
            .O(N__29855),
            .I(N__29845));
    LocalMux I__5045 (
            .O(N__29852),
            .I(N__29840));
    LocalMux I__5044 (
            .O(N__29849),
            .I(N__29840));
    CascadeMux I__5043 (
            .O(N__29848),
            .I(N__29837));
    Span4Mux_v I__5042 (
            .O(N__29845),
            .I(N__29830));
    Span4Mux_v I__5041 (
            .O(N__29840),
            .I(N__29830));
    InMux I__5040 (
            .O(N__29837),
            .I(N__29827));
    InMux I__5039 (
            .O(N__29836),
            .I(N__29822));
    InMux I__5038 (
            .O(N__29835),
            .I(N__29822));
    Odrv4 I__5037 (
            .O(N__29830),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__5036 (
            .O(N__29827),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__5035 (
            .O(N__29822),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    InMux I__5034 (
            .O(N__29815),
            .I(N__29794));
    InMux I__5033 (
            .O(N__29814),
            .I(N__29779));
    InMux I__5032 (
            .O(N__29813),
            .I(N__29779));
    InMux I__5031 (
            .O(N__29812),
            .I(N__29779));
    InMux I__5030 (
            .O(N__29811),
            .I(N__29779));
    InMux I__5029 (
            .O(N__29810),
            .I(N__29779));
    InMux I__5028 (
            .O(N__29809),
            .I(N__29779));
    InMux I__5027 (
            .O(N__29808),
            .I(N__29779));
    InMux I__5026 (
            .O(N__29807),
            .I(N__29766));
    InMux I__5025 (
            .O(N__29806),
            .I(N__29766));
    InMux I__5024 (
            .O(N__29805),
            .I(N__29766));
    InMux I__5023 (
            .O(N__29804),
            .I(N__29766));
    InMux I__5022 (
            .O(N__29803),
            .I(N__29766));
    InMux I__5021 (
            .O(N__29802),
            .I(N__29766));
    InMux I__5020 (
            .O(N__29801),
            .I(N__29755));
    InMux I__5019 (
            .O(N__29800),
            .I(N__29755));
    InMux I__5018 (
            .O(N__29799),
            .I(N__29755));
    InMux I__5017 (
            .O(N__29798),
            .I(N__29755));
    InMux I__5016 (
            .O(N__29797),
            .I(N__29755));
    LocalMux I__5015 (
            .O(N__29794),
            .I(N__29747));
    LocalMux I__5014 (
            .O(N__29779),
            .I(N__29747));
    LocalMux I__5013 (
            .O(N__29766),
            .I(N__29742));
    LocalMux I__5012 (
            .O(N__29755),
            .I(N__29742));
    InMux I__5011 (
            .O(N__29754),
            .I(N__29735));
    InMux I__5010 (
            .O(N__29753),
            .I(N__29735));
    InMux I__5009 (
            .O(N__29752),
            .I(N__29735));
    Span4Mux_v I__5008 (
            .O(N__29747),
            .I(N__29726));
    Span4Mux_v I__5007 (
            .O(N__29742),
            .I(N__29726));
    LocalMux I__5006 (
            .O(N__29735),
            .I(N__29726));
    CascadeMux I__5005 (
            .O(N__29734),
            .I(N__29723));
    CascadeMux I__5004 (
            .O(N__29733),
            .I(N__29720));
    Span4Mux_h I__5003 (
            .O(N__29726),
            .I(N__29717));
    InMux I__5002 (
            .O(N__29723),
            .I(N__29714));
    InMux I__5001 (
            .O(N__29720),
            .I(N__29711));
    Span4Mux_v I__5000 (
            .O(N__29717),
            .I(N__29708));
    LocalMux I__4999 (
            .O(N__29714),
            .I(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0 ));
    LocalMux I__4998 (
            .O(N__29711),
            .I(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__4997 (
            .O(N__29708),
            .I(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0 ));
    InMux I__4996 (
            .O(N__29701),
            .I(N__29686));
    InMux I__4995 (
            .O(N__29700),
            .I(N__29671));
    InMux I__4994 (
            .O(N__29699),
            .I(N__29671));
    InMux I__4993 (
            .O(N__29698),
            .I(N__29671));
    InMux I__4992 (
            .O(N__29697),
            .I(N__29671));
    InMux I__4991 (
            .O(N__29696),
            .I(N__29671));
    InMux I__4990 (
            .O(N__29695),
            .I(N__29671));
    InMux I__4989 (
            .O(N__29694),
            .I(N__29671));
    InMux I__4988 (
            .O(N__29693),
            .I(N__29660));
    InMux I__4987 (
            .O(N__29692),
            .I(N__29660));
    InMux I__4986 (
            .O(N__29691),
            .I(N__29660));
    InMux I__4985 (
            .O(N__29690),
            .I(N__29660));
    InMux I__4984 (
            .O(N__29689),
            .I(N__29660));
    LocalMux I__4983 (
            .O(N__29686),
            .I(N__29646));
    LocalMux I__4982 (
            .O(N__29671),
            .I(N__29646));
    LocalMux I__4981 (
            .O(N__29660),
            .I(N__29643));
    InMux I__4980 (
            .O(N__29659),
            .I(N__29640));
    InMux I__4979 (
            .O(N__29658),
            .I(N__29635));
    InMux I__4978 (
            .O(N__29657),
            .I(N__29635));
    InMux I__4977 (
            .O(N__29656),
            .I(N__29622));
    InMux I__4976 (
            .O(N__29655),
            .I(N__29622));
    InMux I__4975 (
            .O(N__29654),
            .I(N__29622));
    InMux I__4974 (
            .O(N__29653),
            .I(N__29622));
    InMux I__4973 (
            .O(N__29652),
            .I(N__29622));
    InMux I__4972 (
            .O(N__29651),
            .I(N__29622));
    Span4Mux_v I__4971 (
            .O(N__29646),
            .I(N__29613));
    Span4Mux_v I__4970 (
            .O(N__29643),
            .I(N__29613));
    LocalMux I__4969 (
            .O(N__29640),
            .I(N__29613));
    LocalMux I__4968 (
            .O(N__29635),
            .I(N__29613));
    LocalMux I__4967 (
            .O(N__29622),
            .I(N__29608));
    Span4Mux_h I__4966 (
            .O(N__29613),
            .I(N__29605));
    InMux I__4965 (
            .O(N__29612),
            .I(N__29600));
    InMux I__4964 (
            .O(N__29611),
            .I(N__29600));
    Span4Mux_h I__4963 (
            .O(N__29608),
            .I(N__29597));
    Span4Mux_v I__4962 (
            .O(N__29605),
            .I(N__29594));
    LocalMux I__4961 (
            .O(N__29600),
            .I(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__4960 (
            .O(N__29597),
            .I(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__4959 (
            .O(N__29594),
            .I(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1 ));
    CascadeMux I__4958 (
            .O(N__29587),
            .I(N__29584));
    InMux I__4957 (
            .O(N__29584),
            .I(N__29581));
    LocalMux I__4956 (
            .O(N__29581),
            .I(N__29578));
    Span4Mux_v I__4955 (
            .O(N__29578),
            .I(N__29575));
    Odrv4 I__4954 (
            .O(N__29575),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ));
    CascadeMux I__4953 (
            .O(N__29572),
            .I(N__29569));
    InMux I__4952 (
            .O(N__29569),
            .I(N__29566));
    LocalMux I__4951 (
            .O(N__29566),
            .I(N__29563));
    Span4Mux_h I__4950 (
            .O(N__29563),
            .I(N__29560));
    Odrv4 I__4949 (
            .O(N__29560),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ));
    InMux I__4948 (
            .O(N__29557),
            .I(N__29554));
    LocalMux I__4947 (
            .O(N__29554),
            .I(\current_shift_inst.un4_control_input1_1 ));
    CascadeMux I__4946 (
            .O(N__29551),
            .I(\current_shift_inst.un4_control_input1_1_cascade_ ));
    CascadeMux I__4945 (
            .O(N__29548),
            .I(N__29545));
    InMux I__4944 (
            .O(N__29545),
            .I(N__29542));
    LocalMux I__4943 (
            .O(N__29542),
            .I(N__29539));
    Odrv4 I__4942 (
            .O(N__29539),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ));
    CascadeMux I__4941 (
            .O(N__29536),
            .I(N__29533));
    InMux I__4940 (
            .O(N__29533),
            .I(N__29530));
    LocalMux I__4939 (
            .O(N__29530),
            .I(N__29527));
    Odrv4 I__4938 (
            .O(N__29527),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ));
    CascadeMux I__4937 (
            .O(N__29524),
            .I(N__29521));
    InMux I__4936 (
            .O(N__29521),
            .I(N__29518));
    LocalMux I__4935 (
            .O(N__29518),
            .I(N__29515));
    Odrv4 I__4934 (
            .O(N__29515),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ));
    CascadeMux I__4933 (
            .O(N__29512),
            .I(N__29509));
    InMux I__4932 (
            .O(N__29509),
            .I(N__29506));
    LocalMux I__4931 (
            .O(N__29506),
            .I(N__29503));
    Odrv4 I__4930 (
            .O(N__29503),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ));
    CascadeMux I__4929 (
            .O(N__29500),
            .I(\delay_measurement_inst.N_265_cascade_ ));
    InMux I__4928 (
            .O(N__29497),
            .I(N__29491));
    InMux I__4927 (
            .O(N__29496),
            .I(N__29491));
    LocalMux I__4926 (
            .O(N__29491),
            .I(N__29484));
    InMux I__4925 (
            .O(N__29490),
            .I(N__29475));
    InMux I__4924 (
            .O(N__29489),
            .I(N__29475));
    InMux I__4923 (
            .O(N__29488),
            .I(N__29475));
    InMux I__4922 (
            .O(N__29487),
            .I(N__29475));
    Odrv4 I__4921 (
            .O(N__29484),
            .I(\delay_measurement_inst.N_270 ));
    LocalMux I__4920 (
            .O(N__29475),
            .I(\delay_measurement_inst.N_270 ));
    InMux I__4919 (
            .O(N__29470),
            .I(N__29467));
    LocalMux I__4918 (
            .O(N__29467),
            .I(N__29464));
    Odrv4 I__4917 (
            .O(N__29464),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19 ));
    InMux I__4916 (
            .O(N__29461),
            .I(N__29458));
    LocalMux I__4915 (
            .O(N__29458),
            .I(N__29453));
    InMux I__4914 (
            .O(N__29457),
            .I(N__29450));
    InMux I__4913 (
            .O(N__29456),
            .I(N__29447));
    Span4Mux_v I__4912 (
            .O(N__29453),
            .I(N__29444));
    LocalMux I__4911 (
            .O(N__29450),
            .I(N__29440));
    LocalMux I__4910 (
            .O(N__29447),
            .I(N__29437));
    Span4Mux_h I__4909 (
            .O(N__29444),
            .I(N__29434));
    InMux I__4908 (
            .O(N__29443),
            .I(N__29431));
    Span4Mux_v I__4907 (
            .O(N__29440),
            .I(N__29426));
    Span4Mux_v I__4906 (
            .O(N__29437),
            .I(N__29426));
    Odrv4 I__4905 (
            .O(N__29434),
            .I(measured_delay_tr_17));
    LocalMux I__4904 (
            .O(N__29431),
            .I(measured_delay_tr_17));
    Odrv4 I__4903 (
            .O(N__29426),
            .I(measured_delay_tr_17));
    InMux I__4902 (
            .O(N__29419),
            .I(N__29414));
    InMux I__4901 (
            .O(N__29418),
            .I(N__29411));
    InMux I__4900 (
            .O(N__29417),
            .I(N__29408));
    LocalMux I__4899 (
            .O(N__29414),
            .I(N__29404));
    LocalMux I__4898 (
            .O(N__29411),
            .I(N__29399));
    LocalMux I__4897 (
            .O(N__29408),
            .I(N__29399));
    InMux I__4896 (
            .O(N__29407),
            .I(N__29396));
    Span4Mux_h I__4895 (
            .O(N__29404),
            .I(N__29391));
    Span4Mux_h I__4894 (
            .O(N__29399),
            .I(N__29391));
    LocalMux I__4893 (
            .O(N__29396),
            .I(measured_delay_tr_18));
    Odrv4 I__4892 (
            .O(N__29391),
            .I(measured_delay_tr_18));
    InMux I__4891 (
            .O(N__29386),
            .I(N__29376));
    InMux I__4890 (
            .O(N__29385),
            .I(N__29376));
    InMux I__4889 (
            .O(N__29384),
            .I(N__29376));
    InMux I__4888 (
            .O(N__29383),
            .I(N__29370));
    LocalMux I__4887 (
            .O(N__29376),
            .I(N__29367));
    InMux I__4886 (
            .O(N__29375),
            .I(N__29362));
    InMux I__4885 (
            .O(N__29374),
            .I(N__29362));
    InMux I__4884 (
            .O(N__29373),
            .I(N__29359));
    LocalMux I__4883 (
            .O(N__29370),
            .I(N__29354));
    Span4Mux_v I__4882 (
            .O(N__29367),
            .I(N__29347));
    LocalMux I__4881 (
            .O(N__29362),
            .I(N__29347));
    LocalMux I__4880 (
            .O(N__29359),
            .I(N__29347));
    InMux I__4879 (
            .O(N__29358),
            .I(N__29342));
    InMux I__4878 (
            .O(N__29357),
            .I(N__29342));
    Odrv4 I__4877 (
            .O(N__29354),
            .I(\delay_measurement_inst.N_325 ));
    Odrv4 I__4876 (
            .O(N__29347),
            .I(\delay_measurement_inst.N_325 ));
    LocalMux I__4875 (
            .O(N__29342),
            .I(\delay_measurement_inst.N_325 ));
    CascadeMux I__4874 (
            .O(N__29335),
            .I(N__29330));
    InMux I__4873 (
            .O(N__29334),
            .I(N__29326));
    InMux I__4872 (
            .O(N__29333),
            .I(N__29323));
    InMux I__4871 (
            .O(N__29330),
            .I(N__29320));
    CascadeMux I__4870 (
            .O(N__29329),
            .I(N__29317));
    LocalMux I__4869 (
            .O(N__29326),
            .I(N__29314));
    LocalMux I__4868 (
            .O(N__29323),
            .I(N__29309));
    LocalMux I__4867 (
            .O(N__29320),
            .I(N__29309));
    InMux I__4866 (
            .O(N__29317),
            .I(N__29306));
    Span4Mux_h I__4865 (
            .O(N__29314),
            .I(N__29301));
    Span4Mux_h I__4864 (
            .O(N__29309),
            .I(N__29301));
    LocalMux I__4863 (
            .O(N__29306),
            .I(measured_delay_tr_19));
    Odrv4 I__4862 (
            .O(N__29301),
            .I(measured_delay_tr_19));
    CEMux I__4861 (
            .O(N__29296),
            .I(N__29293));
    LocalMux I__4860 (
            .O(N__29293),
            .I(N__29290));
    Sp12to4 I__4859 (
            .O(N__29290),
            .I(N__29284));
    CEMux I__4858 (
            .O(N__29289),
            .I(N__29281));
    CEMux I__4857 (
            .O(N__29288),
            .I(N__29278));
    CEMux I__4856 (
            .O(N__29287),
            .I(N__29275));
    Odrv12 I__4855 (
            .O(N__29284),
            .I(\delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ));
    LocalMux I__4854 (
            .O(N__29281),
            .I(\delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ));
    LocalMux I__4853 (
            .O(N__29278),
            .I(\delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ));
    LocalMux I__4852 (
            .O(N__29275),
            .I(\delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ));
    InMux I__4851 (
            .O(N__29266),
            .I(N__29263));
    LocalMux I__4850 (
            .O(N__29263),
            .I(\current_shift_inst.elapsed_time_ns_s1_fast_31 ));
    CascadeMux I__4849 (
            .O(N__29260),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10_cascade_ ));
    InMux I__4848 (
            .O(N__29257),
            .I(N__29254));
    LocalMux I__4847 (
            .O(N__29254),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_5 ));
    CascadeMux I__4846 (
            .O(N__29251),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_0_cascade_ ));
    InMux I__4845 (
            .O(N__29248),
            .I(N__29244));
    InMux I__4844 (
            .O(N__29247),
            .I(N__29241));
    LocalMux I__4843 (
            .O(N__29244),
            .I(N__29236));
    LocalMux I__4842 (
            .O(N__29241),
            .I(N__29236));
    Odrv4 I__4841 (
            .O(N__29236),
            .I(\delay_measurement_inst.un3_elapsed_time_tr_0_i ));
    CascadeMux I__4840 (
            .O(N__29233),
            .I(\delay_measurement_inst.un3_elapsed_time_tr_0_i_cascade_ ));
    InMux I__4839 (
            .O(N__29230),
            .I(N__29227));
    LocalMux I__4838 (
            .O(N__29227),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_5 ));
    InMux I__4837 (
            .O(N__29224),
            .I(N__29218));
    InMux I__4836 (
            .O(N__29223),
            .I(N__29218));
    LocalMux I__4835 (
            .O(N__29218),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6Z0Z_7 ));
    InMux I__4834 (
            .O(N__29215),
            .I(N__29204));
    InMux I__4833 (
            .O(N__29214),
            .I(N__29204));
    InMux I__4832 (
            .O(N__29213),
            .I(N__29195));
    InMux I__4831 (
            .O(N__29212),
            .I(N__29195));
    InMux I__4830 (
            .O(N__29211),
            .I(N__29195));
    InMux I__4829 (
            .O(N__29210),
            .I(N__29195));
    InMux I__4828 (
            .O(N__29209),
            .I(N__29192));
    LocalMux I__4827 (
            .O(N__29204),
            .I(\delay_measurement_inst.N_299 ));
    LocalMux I__4826 (
            .O(N__29195),
            .I(\delay_measurement_inst.N_299 ));
    LocalMux I__4825 (
            .O(N__29192),
            .I(\delay_measurement_inst.N_299 ));
    CascadeMux I__4824 (
            .O(N__29185),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3_cascade_ ));
    InMux I__4823 (
            .O(N__29182),
            .I(N__29179));
    LocalMux I__4822 (
            .O(N__29179),
            .I(\delay_measurement_inst.delay_tr_timer.N_287_4 ));
    InMux I__4821 (
            .O(N__29176),
            .I(N__29173));
    LocalMux I__4820 (
            .O(N__29173),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6 ));
    InMux I__4819 (
            .O(N__29170),
            .I(N__29167));
    LocalMux I__4818 (
            .O(N__29167),
            .I(N__29163));
    InMux I__4817 (
            .O(N__29166),
            .I(N__29159));
    Span4Mux_v I__4816 (
            .O(N__29163),
            .I(N__29156));
    InMux I__4815 (
            .O(N__29162),
            .I(N__29153));
    LocalMux I__4814 (
            .O(N__29159),
            .I(\delay_measurement_inst.N_265 ));
    Odrv4 I__4813 (
            .O(N__29156),
            .I(\delay_measurement_inst.N_265 ));
    LocalMux I__4812 (
            .O(N__29153),
            .I(\delay_measurement_inst.N_265 ));
    InMux I__4811 (
            .O(N__29146),
            .I(N__29143));
    LocalMux I__4810 (
            .O(N__29143),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ));
    InMux I__4809 (
            .O(N__29140),
            .I(N__29137));
    LocalMux I__4808 (
            .O(N__29137),
            .I(N__29134));
    Span4Mux_h I__4807 (
            .O(N__29134),
            .I(N__29131));
    Odrv4 I__4806 (
            .O(N__29131),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ));
    InMux I__4805 (
            .O(N__29128),
            .I(N__29125));
    LocalMux I__4804 (
            .O(N__29125),
            .I(N__29122));
    Odrv4 I__4803 (
            .O(N__29122),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3 ));
    CascadeMux I__4802 (
            .O(N__29119),
            .I(\delay_measurement_inst.delay_tr_timer.N_287_4_cascade_ ));
    InMux I__4801 (
            .O(N__29116),
            .I(N__29113));
    LocalMux I__4800 (
            .O(N__29113),
            .I(N__29110));
    Odrv4 I__4799 (
            .O(N__29110),
            .I(\delay_measurement_inst.delay_tr_timer.N_290 ));
    CascadeMux I__4798 (
            .O(N__29107),
            .I(N__29104));
    InMux I__4797 (
            .O(N__29104),
            .I(N__29101));
    LocalMux I__4796 (
            .O(N__29101),
            .I(\delay_measurement_inst.N_59 ));
    InMux I__4795 (
            .O(N__29098),
            .I(N__29092));
    InMux I__4794 (
            .O(N__29097),
            .I(N__29092));
    LocalMux I__4793 (
            .O(N__29092),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10 ));
    CascadeMux I__4792 (
            .O(N__29089),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_ ));
    InMux I__4791 (
            .O(N__29086),
            .I(N__29083));
    LocalMux I__4790 (
            .O(N__29083),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ));
    InMux I__4789 (
            .O(N__29080),
            .I(N__29077));
    LocalMux I__4788 (
            .O(N__29077),
            .I(N__29074));
    Odrv12 I__4787 (
            .O(N__29074),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_7 ));
    InMux I__4786 (
            .O(N__29071),
            .I(N__29068));
    LocalMux I__4785 (
            .O(N__29068),
            .I(N__29065));
    Odrv12 I__4784 (
            .O(N__29065),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_15 ));
    InMux I__4783 (
            .O(N__29062),
            .I(N__29059));
    LocalMux I__4782 (
            .O(N__29059),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ));
    CascadeMux I__4781 (
            .O(N__29056),
            .I(N__29048));
    CascadeMux I__4780 (
            .O(N__29055),
            .I(N__29045));
    CascadeMux I__4779 (
            .O(N__29054),
            .I(N__29042));
    CascadeMux I__4778 (
            .O(N__29053),
            .I(N__29039));
    InMux I__4777 (
            .O(N__29052),
            .I(N__29030));
    InMux I__4776 (
            .O(N__29051),
            .I(N__29030));
    InMux I__4775 (
            .O(N__29048),
            .I(N__29030));
    InMux I__4774 (
            .O(N__29045),
            .I(N__29030));
    InMux I__4773 (
            .O(N__29042),
            .I(N__29023));
    InMux I__4772 (
            .O(N__29039),
            .I(N__29023));
    LocalMux I__4771 (
            .O(N__29030),
            .I(N__29020));
    InMux I__4770 (
            .O(N__29029),
            .I(N__29017));
    InMux I__4769 (
            .O(N__29028),
            .I(N__29014));
    LocalMux I__4768 (
            .O(N__29023),
            .I(N__29005));
    Span4Mux_h I__4767 (
            .O(N__29020),
            .I(N__29005));
    LocalMux I__4766 (
            .O(N__29017),
            .I(N__29005));
    LocalMux I__4765 (
            .O(N__29014),
            .I(N__29005));
    Odrv4 I__4764 (
            .O(N__29005),
            .I(\delay_measurement_inst.N_267 ));
    InMux I__4763 (
            .O(N__29002),
            .I(N__28999));
    LocalMux I__4762 (
            .O(N__28999),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3 ));
    CascadeMux I__4761 (
            .O(N__28996),
            .I(N__28993));
    InMux I__4760 (
            .O(N__28993),
            .I(N__28990));
    LocalMux I__4759 (
            .O(N__28990),
            .I(N__28987));
    Odrv4 I__4758 (
            .O(N__28987),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ));
    CascadeMux I__4757 (
            .O(N__28984),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_ ));
    CascadeMux I__4756 (
            .O(N__28981),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_ ));
    CascadeMux I__4755 (
            .O(N__28978),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ));
    InMux I__4754 (
            .O(N__28975),
            .I(N__28972));
    LocalMux I__4753 (
            .O(N__28972),
            .I(\current_shift_inst.PI_CTRL.N_72 ));
    InMux I__4752 (
            .O(N__28969),
            .I(N__28966));
    LocalMux I__4751 (
            .O(N__28966),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ));
    CascadeMux I__4750 (
            .O(N__28963),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_18_cascade_ ));
    InMux I__4749 (
            .O(N__28960),
            .I(N__28957));
    LocalMux I__4748 (
            .O(N__28957),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ));
    CascadeMux I__4747 (
            .O(N__28954),
            .I(N__28951));
    InMux I__4746 (
            .O(N__28951),
            .I(N__28948));
    LocalMux I__4745 (
            .O(N__28948),
            .I(N__28945));
    Span4Mux_h I__4744 (
            .O(N__28945),
            .I(N__28942));
    Odrv4 I__4743 (
            .O(N__28942),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ));
    CascadeMux I__4742 (
            .O(N__28939),
            .I(N__28936));
    InMux I__4741 (
            .O(N__28936),
            .I(N__28933));
    LocalMux I__4740 (
            .O(N__28933),
            .I(N__28930));
    Span4Mux_h I__4739 (
            .O(N__28930),
            .I(N__28927));
    Odrv4 I__4738 (
            .O(N__28927),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ));
    CascadeMux I__4737 (
            .O(N__28924),
            .I(N__28921));
    InMux I__4736 (
            .O(N__28921),
            .I(N__28918));
    LocalMux I__4735 (
            .O(N__28918),
            .I(N__28915));
    Span4Mux_h I__4734 (
            .O(N__28915),
            .I(N__28912));
    Odrv4 I__4733 (
            .O(N__28912),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ));
    CascadeMux I__4732 (
            .O(N__28909),
            .I(N__28906));
    InMux I__4731 (
            .O(N__28906),
            .I(N__28903));
    LocalMux I__4730 (
            .O(N__28903),
            .I(N__28900));
    Odrv12 I__4729 (
            .O(N__28900),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ));
    CascadeMux I__4728 (
            .O(N__28897),
            .I(N__28894));
    InMux I__4727 (
            .O(N__28894),
            .I(N__28891));
    LocalMux I__4726 (
            .O(N__28891),
            .I(N__28888));
    Span4Mux_h I__4725 (
            .O(N__28888),
            .I(N__28885));
    Odrv4 I__4724 (
            .O(N__28885),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ));
    CascadeMux I__4723 (
            .O(N__28882),
            .I(N__28879));
    InMux I__4722 (
            .O(N__28879),
            .I(N__28876));
    LocalMux I__4721 (
            .O(N__28876),
            .I(N__28873));
    Span4Mux_h I__4720 (
            .O(N__28873),
            .I(N__28870));
    Odrv4 I__4719 (
            .O(N__28870),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ));
    CascadeMux I__4718 (
            .O(N__28867),
            .I(N__28864));
    InMux I__4717 (
            .O(N__28864),
            .I(N__28861));
    LocalMux I__4716 (
            .O(N__28861),
            .I(N__28858));
    Odrv4 I__4715 (
            .O(N__28858),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ));
    CascadeMux I__4714 (
            .O(N__28855),
            .I(N__28852));
    InMux I__4713 (
            .O(N__28852),
            .I(N__28849));
    LocalMux I__4712 (
            .O(N__28849),
            .I(N__28846));
    Odrv4 I__4711 (
            .O(N__28846),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ));
    CascadeMux I__4710 (
            .O(N__28843),
            .I(N__28840));
    InMux I__4709 (
            .O(N__28840),
            .I(N__28837));
    LocalMux I__4708 (
            .O(N__28837),
            .I(N__28834));
    Odrv4 I__4707 (
            .O(N__28834),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ));
    InMux I__4706 (
            .O(N__28831),
            .I(N__28825));
    InMux I__4705 (
            .O(N__28830),
            .I(N__28818));
    InMux I__4704 (
            .O(N__28829),
            .I(N__28818));
    InMux I__4703 (
            .O(N__28828),
            .I(N__28818));
    LocalMux I__4702 (
            .O(N__28825),
            .I(N__28815));
    LocalMux I__4701 (
            .O(N__28818),
            .I(N__28812));
    Odrv4 I__4700 (
            .O(N__28815),
            .I(\phase_controller_inst1.stoper_hc.time_passed11 ));
    Odrv4 I__4699 (
            .O(N__28812),
            .I(\phase_controller_inst1.stoper_hc.time_passed11 ));
    InMux I__4698 (
            .O(N__28807),
            .I(N__28803));
    InMux I__4697 (
            .O(N__28806),
            .I(N__28800));
    LocalMux I__4696 (
            .O(N__28803),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    LocalMux I__4695 (
            .O(N__28800),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__4694 (
            .O(N__28795),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_17 ));
    CascadeMux I__4693 (
            .O(N__28792),
            .I(N__28789));
    InMux I__4692 (
            .O(N__28789),
            .I(N__28786));
    LocalMux I__4691 (
            .O(N__28786),
            .I(N__28783));
    Odrv4 I__4690 (
            .O(N__28783),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_19 ));
    CascadeMux I__4689 (
            .O(N__28780),
            .I(N__28777));
    InMux I__4688 (
            .O(N__28777),
            .I(N__28774));
    LocalMux I__4687 (
            .O(N__28774),
            .I(N__28771));
    Odrv4 I__4686 (
            .O(N__28771),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ));
    CascadeMux I__4685 (
            .O(N__28768),
            .I(N__28765));
    InMux I__4684 (
            .O(N__28765),
            .I(N__28762));
    LocalMux I__4683 (
            .O(N__28762),
            .I(N__28759));
    Span4Mux_h I__4682 (
            .O(N__28759),
            .I(N__28756));
    Odrv4 I__4681 (
            .O(N__28756),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ));
    CascadeMux I__4680 (
            .O(N__28753),
            .I(N__28750));
    InMux I__4679 (
            .O(N__28750),
            .I(N__28747));
    LocalMux I__4678 (
            .O(N__28747),
            .I(N__28744));
    Span4Mux_h I__4677 (
            .O(N__28744),
            .I(N__28741));
    Odrv4 I__4676 (
            .O(N__28741),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ));
    CascadeMux I__4675 (
            .O(N__28738),
            .I(N__28735));
    InMux I__4674 (
            .O(N__28735),
            .I(N__28732));
    LocalMux I__4673 (
            .O(N__28732),
            .I(N__28729));
    Span4Mux_v I__4672 (
            .O(N__28729),
            .I(N__28726));
    Odrv4 I__4671 (
            .O(N__28726),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ));
    CascadeMux I__4670 (
            .O(N__28723),
            .I(N__28720));
    InMux I__4669 (
            .O(N__28720),
            .I(N__28717));
    LocalMux I__4668 (
            .O(N__28717),
            .I(N__28714));
    Odrv4 I__4667 (
            .O(N__28714),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ));
    CascadeMux I__4666 (
            .O(N__28711),
            .I(N__28708));
    InMux I__4665 (
            .O(N__28708),
            .I(N__28705));
    LocalMux I__4664 (
            .O(N__28705),
            .I(N__28702));
    Span4Mux_h I__4663 (
            .O(N__28702),
            .I(N__28699));
    Odrv4 I__4662 (
            .O(N__28699),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ));
    CascadeMux I__4661 (
            .O(N__28696),
            .I(N__28693));
    InMux I__4660 (
            .O(N__28693),
            .I(N__28690));
    LocalMux I__4659 (
            .O(N__28690),
            .I(N__28687));
    Odrv12 I__4658 (
            .O(N__28687),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ1Z_6 ));
    CascadeMux I__4657 (
            .O(N__28684),
            .I(N__28681));
    InMux I__4656 (
            .O(N__28681),
            .I(N__28678));
    LocalMux I__4655 (
            .O(N__28678),
            .I(N__28675));
    Span4Mux_h I__4654 (
            .O(N__28675),
            .I(N__28672));
    Odrv4 I__4653 (
            .O(N__28672),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ));
    InMux I__4652 (
            .O(N__28669),
            .I(N__28666));
    LocalMux I__4651 (
            .O(N__28666),
            .I(N__28663));
    Span4Mux_h I__4650 (
            .O(N__28663),
            .I(N__28659));
    InMux I__4649 (
            .O(N__28662),
            .I(N__28656));
    Odrv4 I__4648 (
            .O(N__28659),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ));
    LocalMux I__4647 (
            .O(N__28656),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ));
    CascadeMux I__4646 (
            .O(N__28651),
            .I(N__28648));
    InMux I__4645 (
            .O(N__28648),
            .I(N__28645));
    LocalMux I__4644 (
            .O(N__28645),
            .I(N__28642));
    Span4Mux_h I__4643 (
            .O(N__28642),
            .I(N__28639));
    Odrv4 I__4642 (
            .O(N__28639),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_11 ));
    InMux I__4641 (
            .O(N__28636),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_9 ));
    InMux I__4640 (
            .O(N__28633),
            .I(N__28629));
    InMux I__4639 (
            .O(N__28632),
            .I(N__28626));
    LocalMux I__4638 (
            .O(N__28629),
            .I(N__28623));
    LocalMux I__4637 (
            .O(N__28626),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    Odrv4 I__4636 (
            .O(N__28623),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__4635 (
            .O(N__28618),
            .I(N__28615));
    LocalMux I__4634 (
            .O(N__28615),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_12 ));
    InMux I__4633 (
            .O(N__28612),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_10 ));
    InMux I__4632 (
            .O(N__28609),
            .I(N__28605));
    InMux I__4631 (
            .O(N__28608),
            .I(N__28602));
    LocalMux I__4630 (
            .O(N__28605),
            .I(N__28599));
    LocalMux I__4629 (
            .O(N__28602),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ));
    Odrv4 I__4628 (
            .O(N__28599),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ));
    CascadeMux I__4627 (
            .O(N__28594),
            .I(N__28591));
    InMux I__4626 (
            .O(N__28591),
            .I(N__28588));
    LocalMux I__4625 (
            .O(N__28588),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_13 ));
    InMux I__4624 (
            .O(N__28585),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_11 ));
    InMux I__4623 (
            .O(N__28582),
            .I(N__28578));
    InMux I__4622 (
            .O(N__28581),
            .I(N__28575));
    LocalMux I__4621 (
            .O(N__28578),
            .I(N__28572));
    LocalMux I__4620 (
            .O(N__28575),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    Odrv4 I__4619 (
            .O(N__28572),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    InMux I__4618 (
            .O(N__28567),
            .I(N__28564));
    LocalMux I__4617 (
            .O(N__28564),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_14 ));
    InMux I__4616 (
            .O(N__28561),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_12 ));
    InMux I__4615 (
            .O(N__28558),
            .I(N__28554));
    InMux I__4614 (
            .O(N__28557),
            .I(N__28551));
    LocalMux I__4613 (
            .O(N__28554),
            .I(N__28548));
    LocalMux I__4612 (
            .O(N__28551),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    Odrv4 I__4611 (
            .O(N__28548),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    CascadeMux I__4610 (
            .O(N__28543),
            .I(N__28540));
    InMux I__4609 (
            .O(N__28540),
            .I(N__28537));
    LocalMux I__4608 (
            .O(N__28537),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_15 ));
    InMux I__4607 (
            .O(N__28534),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_13 ));
    InMux I__4606 (
            .O(N__28531),
            .I(N__28527));
    InMux I__4605 (
            .O(N__28530),
            .I(N__28524));
    LocalMux I__4604 (
            .O(N__28527),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    LocalMux I__4603 (
            .O(N__28524),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    InMux I__4602 (
            .O(N__28519),
            .I(N__28516));
    LocalMux I__4601 (
            .O(N__28516),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_16 ));
    InMux I__4600 (
            .O(N__28513),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_14 ));
    InMux I__4599 (
            .O(N__28510),
            .I(N__28506));
    InMux I__4598 (
            .O(N__28509),
            .I(N__28503));
    LocalMux I__4597 (
            .O(N__28506),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ));
    LocalMux I__4596 (
            .O(N__28503),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ));
    CascadeMux I__4595 (
            .O(N__28498),
            .I(N__28495));
    InMux I__4594 (
            .O(N__28495),
            .I(N__28492));
    LocalMux I__4593 (
            .O(N__28492),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_17 ));
    InMux I__4592 (
            .O(N__28489),
            .I(bfn_11_20_0_));
    InMux I__4591 (
            .O(N__28486),
            .I(N__28482));
    InMux I__4590 (
            .O(N__28485),
            .I(N__28479));
    LocalMux I__4589 (
            .O(N__28482),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    LocalMux I__4588 (
            .O(N__28479),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__4587 (
            .O(N__28474),
            .I(N__28471));
    LocalMux I__4586 (
            .O(N__28471),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_18 ));
    InMux I__4585 (
            .O(N__28468),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_16 ));
    CascadeMux I__4584 (
            .O(N__28465),
            .I(N__28462));
    InMux I__4583 (
            .O(N__28462),
            .I(N__28458));
    InMux I__4582 (
            .O(N__28461),
            .I(N__28455));
    LocalMux I__4581 (
            .O(N__28458),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    LocalMux I__4580 (
            .O(N__28455),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    InMux I__4579 (
            .O(N__28450),
            .I(N__28447));
    LocalMux I__4578 (
            .O(N__28447),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_3 ));
    InMux I__4577 (
            .O(N__28444),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_1 ));
    InMux I__4576 (
            .O(N__28441),
            .I(N__28437));
    InMux I__4575 (
            .O(N__28440),
            .I(N__28434));
    LocalMux I__4574 (
            .O(N__28437),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    LocalMux I__4573 (
            .O(N__28434),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    CascadeMux I__4572 (
            .O(N__28429),
            .I(N__28426));
    InMux I__4571 (
            .O(N__28426),
            .I(N__28423));
    LocalMux I__4570 (
            .O(N__28423),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_4 ));
    InMux I__4569 (
            .O(N__28420),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_2 ));
    InMux I__4568 (
            .O(N__28417),
            .I(N__28413));
    InMux I__4567 (
            .O(N__28416),
            .I(N__28410));
    LocalMux I__4566 (
            .O(N__28413),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    LocalMux I__4565 (
            .O(N__28410),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    InMux I__4564 (
            .O(N__28405),
            .I(N__28402));
    LocalMux I__4563 (
            .O(N__28402),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_5 ));
    InMux I__4562 (
            .O(N__28399),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_3 ));
    InMux I__4561 (
            .O(N__28396),
            .I(N__28392));
    InMux I__4560 (
            .O(N__28395),
            .I(N__28389));
    LocalMux I__4559 (
            .O(N__28392),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    LocalMux I__4558 (
            .O(N__28389),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    CascadeMux I__4557 (
            .O(N__28384),
            .I(N__28381));
    InMux I__4556 (
            .O(N__28381),
            .I(N__28378));
    LocalMux I__4555 (
            .O(N__28378),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_6 ));
    InMux I__4554 (
            .O(N__28375),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_4 ));
    InMux I__4553 (
            .O(N__28372),
            .I(N__28368));
    InMux I__4552 (
            .O(N__28371),
            .I(N__28365));
    LocalMux I__4551 (
            .O(N__28368),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    LocalMux I__4550 (
            .O(N__28365),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    InMux I__4549 (
            .O(N__28360),
            .I(N__28357));
    LocalMux I__4548 (
            .O(N__28357),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_7 ));
    InMux I__4547 (
            .O(N__28354),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_5 ));
    InMux I__4546 (
            .O(N__28351),
            .I(N__28347));
    InMux I__4545 (
            .O(N__28350),
            .I(N__28344));
    LocalMux I__4544 (
            .O(N__28347),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    LocalMux I__4543 (
            .O(N__28344),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    CascadeMux I__4542 (
            .O(N__28339),
            .I(N__28336));
    InMux I__4541 (
            .O(N__28336),
            .I(N__28333));
    LocalMux I__4540 (
            .O(N__28333),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_8 ));
    InMux I__4539 (
            .O(N__28330),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_6 ));
    InMux I__4538 (
            .O(N__28327),
            .I(N__28324));
    LocalMux I__4537 (
            .O(N__28324),
            .I(N__28320));
    InMux I__4536 (
            .O(N__28323),
            .I(N__28317));
    Odrv4 I__4535 (
            .O(N__28320),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    LocalMux I__4534 (
            .O(N__28317),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    InMux I__4533 (
            .O(N__28312),
            .I(N__28309));
    LocalMux I__4532 (
            .O(N__28309),
            .I(N__28306));
    Odrv4 I__4531 (
            .O(N__28306),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_9 ));
    InMux I__4530 (
            .O(N__28303),
            .I(bfn_11_19_0_));
    InMux I__4529 (
            .O(N__28300),
            .I(N__28297));
    LocalMux I__4528 (
            .O(N__28297),
            .I(N__28293));
    InMux I__4527 (
            .O(N__28296),
            .I(N__28290));
    Odrv4 I__4526 (
            .O(N__28293),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ));
    LocalMux I__4525 (
            .O(N__28290),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ));
    InMux I__4524 (
            .O(N__28285),
            .I(N__28282));
    LocalMux I__4523 (
            .O(N__28282),
            .I(N__28279));
    Odrv4 I__4522 (
            .O(N__28279),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_10 ));
    InMux I__4521 (
            .O(N__28276),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_8 ));
    InMux I__4520 (
            .O(N__28273),
            .I(N__28270));
    LocalMux I__4519 (
            .O(N__28270),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1 ));
    CascadeMux I__4518 (
            .O(N__28267),
            .I(N__28264));
    InMux I__4517 (
            .O(N__28264),
            .I(N__28261));
    LocalMux I__4516 (
            .O(N__28261),
            .I(N__28256));
    InMux I__4515 (
            .O(N__28260),
            .I(N__28253));
    InMux I__4514 (
            .O(N__28259),
            .I(N__28250));
    Span4Mux_h I__4513 (
            .O(N__28256),
            .I(N__28247));
    LocalMux I__4512 (
            .O(N__28253),
            .I(N__28244));
    LocalMux I__4511 (
            .O(N__28250),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__4510 (
            .O(N__28247),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__4509 (
            .O(N__28244),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    InMux I__4508 (
            .O(N__28237),
            .I(N__28233));
    InMux I__4507 (
            .O(N__28236),
            .I(N__28230));
    LocalMux I__4506 (
            .O(N__28233),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    LocalMux I__4505 (
            .O(N__28230),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    CascadeMux I__4504 (
            .O(N__28225),
            .I(N__28222));
    InMux I__4503 (
            .O(N__28222),
            .I(N__28219));
    LocalMux I__4502 (
            .O(N__28219),
            .I(N__28216));
    Odrv4 I__4501 (
            .O(N__28216),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_2 ));
    InMux I__4500 (
            .O(N__28213),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0 ));
    InMux I__4499 (
            .O(N__28210),
            .I(N__28207));
    LocalMux I__4498 (
            .O(N__28207),
            .I(N__28204));
    Span4Mux_h I__4497 (
            .O(N__28204),
            .I(N__28199));
    InMux I__4496 (
            .O(N__28203),
            .I(N__28196));
    InMux I__4495 (
            .O(N__28202),
            .I(N__28193));
    Odrv4 I__4494 (
            .O(N__28199),
            .I(measured_delay_tr_12));
    LocalMux I__4493 (
            .O(N__28196),
            .I(measured_delay_tr_12));
    LocalMux I__4492 (
            .O(N__28193),
            .I(measured_delay_tr_12));
    InMux I__4491 (
            .O(N__28186),
            .I(N__28183));
    LocalMux I__4490 (
            .O(N__28183),
            .I(N__28180));
    Span4Mux_h I__4489 (
            .O(N__28180),
            .I(N__28175));
    InMux I__4488 (
            .O(N__28179),
            .I(N__28172));
    InMux I__4487 (
            .O(N__28178),
            .I(N__28169));
    Odrv4 I__4486 (
            .O(N__28175),
            .I(measured_delay_tr_11));
    LocalMux I__4485 (
            .O(N__28172),
            .I(measured_delay_tr_11));
    LocalMux I__4484 (
            .O(N__28169),
            .I(measured_delay_tr_11));
    InMux I__4483 (
            .O(N__28162),
            .I(N__28159));
    LocalMux I__4482 (
            .O(N__28159),
            .I(N__28155));
    CascadeMux I__4481 (
            .O(N__28158),
            .I(N__28151));
    Span4Mux_v I__4480 (
            .O(N__28155),
            .I(N__28148));
    InMux I__4479 (
            .O(N__28154),
            .I(N__28145));
    InMux I__4478 (
            .O(N__28151),
            .I(N__28142));
    Odrv4 I__4477 (
            .O(N__28148),
            .I(measured_delay_tr_13));
    LocalMux I__4476 (
            .O(N__28145),
            .I(measured_delay_tr_13));
    LocalMux I__4475 (
            .O(N__28142),
            .I(measured_delay_tr_13));
    InMux I__4474 (
            .O(N__28135),
            .I(N__28132));
    LocalMux I__4473 (
            .O(N__28132),
            .I(N__28128));
    InMux I__4472 (
            .O(N__28131),
            .I(N__28124));
    Span4Mux_v I__4471 (
            .O(N__28128),
            .I(N__28121));
    InMux I__4470 (
            .O(N__28127),
            .I(N__28118));
    LocalMux I__4469 (
            .O(N__28124),
            .I(N__28115));
    Odrv4 I__4468 (
            .O(N__28121),
            .I(measured_delay_tr_10));
    LocalMux I__4467 (
            .O(N__28118),
            .I(measured_delay_tr_10));
    Odrv4 I__4466 (
            .O(N__28115),
            .I(measured_delay_tr_10));
    InMux I__4465 (
            .O(N__28108),
            .I(N__28105));
    LocalMux I__4464 (
            .O(N__28105),
            .I(N__28102));
    Span4Mux_h I__4463 (
            .O(N__28102),
            .I(N__28096));
    InMux I__4462 (
            .O(N__28101),
            .I(N__28093));
    InMux I__4461 (
            .O(N__28100),
            .I(N__28088));
    InMux I__4460 (
            .O(N__28099),
            .I(N__28088));
    Odrv4 I__4459 (
            .O(N__28096),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6 ));
    LocalMux I__4458 (
            .O(N__28093),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6 ));
    LocalMux I__4457 (
            .O(N__28088),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6 ));
    InMux I__4456 (
            .O(N__28081),
            .I(N__28077));
    InMux I__4455 (
            .O(N__28080),
            .I(N__28074));
    LocalMux I__4454 (
            .O(N__28077),
            .I(N__28071));
    LocalMux I__4453 (
            .O(N__28074),
            .I(N__28068));
    Span4Mux_h I__4452 (
            .O(N__28071),
            .I(N__28061));
    Span4Mux_v I__4451 (
            .O(N__28068),
            .I(N__28061));
    InMux I__4450 (
            .O(N__28067),
            .I(N__28058));
    InMux I__4449 (
            .O(N__28066),
            .I(N__28055));
    Span4Mux_v I__4448 (
            .O(N__28061),
            .I(N__28052));
    LocalMux I__4447 (
            .O(N__28058),
            .I(measured_delay_tr_16));
    LocalMux I__4446 (
            .O(N__28055),
            .I(measured_delay_tr_16));
    Odrv4 I__4445 (
            .O(N__28052),
            .I(measured_delay_tr_16));
    CascadeMux I__4444 (
            .O(N__28045),
            .I(N__28042));
    InMux I__4443 (
            .O(N__28042),
            .I(N__28039));
    LocalMux I__4442 (
            .O(N__28039),
            .I(N__28036));
    Odrv12 I__4441 (
            .O(N__28036),
            .I(\phase_controller_inst2.stoper_hc.time_passed_1_sqmuxa ));
    InMux I__4440 (
            .O(N__28033),
            .I(N__28030));
    LocalMux I__4439 (
            .O(N__28030),
            .I(N__28026));
    InMux I__4438 (
            .O(N__28029),
            .I(N__28023));
    Span4Mux_h I__4437 (
            .O(N__28026),
            .I(N__28020));
    LocalMux I__4436 (
            .O(N__28023),
            .I(N__28016));
    Span4Mux_v I__4435 (
            .O(N__28020),
            .I(N__28013));
    InMux I__4434 (
            .O(N__28019),
            .I(N__28010));
    Span4Mux_v I__4433 (
            .O(N__28016),
            .I(N__28007));
    Odrv4 I__4432 (
            .O(N__28013),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    LocalMux I__4431 (
            .O(N__28010),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    Odrv4 I__4430 (
            .O(N__28007),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    InMux I__4429 (
            .O(N__28000),
            .I(N__27996));
    InMux I__4428 (
            .O(N__27999),
            .I(N__27993));
    LocalMux I__4427 (
            .O(N__27996),
            .I(N__27990));
    LocalMux I__4426 (
            .O(N__27993),
            .I(N__27985));
    Span4Mux_v I__4425 (
            .O(N__27990),
            .I(N__27982));
    InMux I__4424 (
            .O(N__27989),
            .I(N__27979));
    InMux I__4423 (
            .O(N__27988),
            .I(N__27976));
    Span4Mux_h I__4422 (
            .O(N__27985),
            .I(N__27971));
    Span4Mux_v I__4421 (
            .O(N__27982),
            .I(N__27971));
    LocalMux I__4420 (
            .O(N__27979),
            .I(N__27968));
    LocalMux I__4419 (
            .O(N__27976),
            .I(\phase_controller_inst2.hc_time_passed ));
    Odrv4 I__4418 (
            .O(N__27971),
            .I(\phase_controller_inst2.hc_time_passed ));
    Odrv12 I__4417 (
            .O(N__27968),
            .I(\phase_controller_inst2.hc_time_passed ));
    InMux I__4416 (
            .O(N__27961),
            .I(N__27958));
    LocalMux I__4415 (
            .O(N__27958),
            .I(N__27955));
    Span4Mux_h I__4414 (
            .O(N__27955),
            .I(N__27952));
    Odrv4 I__4413 (
            .O(N__27952),
            .I(\phase_controller_inst2.start_timer_hc_RNO_0_0 ));
    InMux I__4412 (
            .O(N__27949),
            .I(N__27945));
    InMux I__4411 (
            .O(N__27948),
            .I(N__27942));
    LocalMux I__4410 (
            .O(N__27945),
            .I(N__27938));
    LocalMux I__4409 (
            .O(N__27942),
            .I(N__27935));
    InMux I__4408 (
            .O(N__27941),
            .I(N__27932));
    Span12Mux_v I__4407 (
            .O(N__27938),
            .I(N__27929));
    Span4Mux_v I__4406 (
            .O(N__27935),
            .I(N__27926));
    LocalMux I__4405 (
            .O(N__27932),
            .I(measured_delay_tr_4));
    Odrv12 I__4404 (
            .O(N__27929),
            .I(measured_delay_tr_4));
    Odrv4 I__4403 (
            .O(N__27926),
            .I(measured_delay_tr_4));
    CascadeMux I__4402 (
            .O(N__27919),
            .I(N__27916));
    InMux I__4401 (
            .O(N__27916),
            .I(N__27912));
    InMux I__4400 (
            .O(N__27915),
            .I(N__27909));
    LocalMux I__4399 (
            .O(N__27912),
            .I(N__27905));
    LocalMux I__4398 (
            .O(N__27909),
            .I(N__27902));
    InMux I__4397 (
            .O(N__27908),
            .I(N__27899));
    Span4Mux_v I__4396 (
            .O(N__27905),
            .I(N__27896));
    Span4Mux_v I__4395 (
            .O(N__27902),
            .I(N__27893));
    LocalMux I__4394 (
            .O(N__27899),
            .I(measured_delay_tr_9));
    Odrv4 I__4393 (
            .O(N__27896),
            .I(measured_delay_tr_9));
    Odrv4 I__4392 (
            .O(N__27893),
            .I(measured_delay_tr_9));
    CascadeMux I__4391 (
            .O(N__27886),
            .I(N__27883));
    InMux I__4390 (
            .O(N__27883),
            .I(N__27878));
    InMux I__4389 (
            .O(N__27882),
            .I(N__27875));
    CascadeMux I__4388 (
            .O(N__27881),
            .I(N__27872));
    LocalMux I__4387 (
            .O(N__27878),
            .I(N__27867));
    LocalMux I__4386 (
            .O(N__27875),
            .I(N__27867));
    InMux I__4385 (
            .O(N__27872),
            .I(N__27864));
    Span4Mux_h I__4384 (
            .O(N__27867),
            .I(N__27861));
    LocalMux I__4383 (
            .O(N__27864),
            .I(measured_delay_tr_3));
    Odrv4 I__4382 (
            .O(N__27861),
            .I(measured_delay_tr_3));
    CascadeMux I__4381 (
            .O(N__27856),
            .I(N__27853));
    InMux I__4380 (
            .O(N__27853),
            .I(N__27850));
    LocalMux I__4379 (
            .O(N__27850),
            .I(N__27845));
    InMux I__4378 (
            .O(N__27849),
            .I(N__27842));
    InMux I__4377 (
            .O(N__27848),
            .I(N__27839));
    Span4Mux_h I__4376 (
            .O(N__27845),
            .I(N__27834));
    LocalMux I__4375 (
            .O(N__27842),
            .I(N__27834));
    LocalMux I__4374 (
            .O(N__27839),
            .I(measured_delay_tr_2));
    Odrv4 I__4373 (
            .O(N__27834),
            .I(measured_delay_tr_2));
    InMux I__4372 (
            .O(N__27829),
            .I(N__27825));
    InMux I__4371 (
            .O(N__27828),
            .I(N__27822));
    LocalMux I__4370 (
            .O(N__27825),
            .I(N__27818));
    LocalMux I__4369 (
            .O(N__27822),
            .I(N__27815));
    InMux I__4368 (
            .O(N__27821),
            .I(N__27812));
    Span4Mux_v I__4367 (
            .O(N__27818),
            .I(N__27809));
    Span4Mux_h I__4366 (
            .O(N__27815),
            .I(N__27804));
    LocalMux I__4365 (
            .O(N__27812),
            .I(N__27804));
    Odrv4 I__4364 (
            .O(N__27809),
            .I(measured_delay_tr_6));
    Odrv4 I__4363 (
            .O(N__27804),
            .I(measured_delay_tr_6));
    CascadeMux I__4362 (
            .O(N__27799),
            .I(N__27796));
    InMux I__4361 (
            .O(N__27796),
            .I(N__27793));
    LocalMux I__4360 (
            .O(N__27793),
            .I(N__27789));
    CascadeMux I__4359 (
            .O(N__27792),
            .I(N__27786));
    Span4Mux_h I__4358 (
            .O(N__27789),
            .I(N__27783));
    InMux I__4357 (
            .O(N__27786),
            .I(N__27780));
    Odrv4 I__4356 (
            .O(N__27783),
            .I(measured_delay_tr_1));
    LocalMux I__4355 (
            .O(N__27780),
            .I(measured_delay_tr_1));
    InMux I__4354 (
            .O(N__27775),
            .I(N__27772));
    LocalMux I__4353 (
            .O(N__27772),
            .I(N__27767));
    InMux I__4352 (
            .O(N__27771),
            .I(N__27760));
    InMux I__4351 (
            .O(N__27770),
            .I(N__27760));
    Span4Mux_v I__4350 (
            .O(N__27767),
            .I(N__27757));
    InMux I__4349 (
            .O(N__27766),
            .I(N__27752));
    InMux I__4348 (
            .O(N__27765),
            .I(N__27752));
    LocalMux I__4347 (
            .O(N__27760),
            .I(N__27749));
    Odrv4 I__4346 (
            .O(N__27757),
            .I(measured_delay_tr_14));
    LocalMux I__4345 (
            .O(N__27752),
            .I(measured_delay_tr_14));
    Odrv4 I__4344 (
            .O(N__27749),
            .I(measured_delay_tr_14));
    CascadeMux I__4343 (
            .O(N__27742),
            .I(N__27739));
    InMux I__4342 (
            .O(N__27739),
            .I(N__27736));
    LocalMux I__4341 (
            .O(N__27736),
            .I(N__27733));
    Odrv4 I__4340 (
            .O(N__27733),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_24 ));
    CascadeMux I__4339 (
            .O(N__27730),
            .I(N__27727));
    InMux I__4338 (
            .O(N__27727),
            .I(N__27724));
    LocalMux I__4337 (
            .O(N__27724),
            .I(N__27721));
    Span4Mux_v I__4336 (
            .O(N__27721),
            .I(N__27718));
    Odrv4 I__4335 (
            .O(N__27718),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_21 ));
    InMux I__4334 (
            .O(N__27715),
            .I(N__27712));
    LocalMux I__4333 (
            .O(N__27712),
            .I(N__27707));
    InMux I__4332 (
            .O(N__27711),
            .I(N__27703));
    CascadeMux I__4331 (
            .O(N__27710),
            .I(N__27700));
    Span4Mux_h I__4330 (
            .O(N__27707),
            .I(N__27697));
    InMux I__4329 (
            .O(N__27706),
            .I(N__27694));
    LocalMux I__4328 (
            .O(N__27703),
            .I(N__27691));
    InMux I__4327 (
            .O(N__27700),
            .I(N__27688));
    Span4Mux_v I__4326 (
            .O(N__27697),
            .I(N__27685));
    LocalMux I__4325 (
            .O(N__27694),
            .I(N__27680));
    Span4Mux_v I__4324 (
            .O(N__27691),
            .I(N__27680));
    LocalMux I__4323 (
            .O(N__27688),
            .I(measured_delay_tr_8));
    Odrv4 I__4322 (
            .O(N__27685),
            .I(measured_delay_tr_8));
    Odrv4 I__4321 (
            .O(N__27680),
            .I(measured_delay_tr_8));
    CascadeMux I__4320 (
            .O(N__27673),
            .I(N__27670));
    InMux I__4319 (
            .O(N__27670),
            .I(N__27667));
    LocalMux I__4318 (
            .O(N__27667),
            .I(N__27664));
    Span4Mux_h I__4317 (
            .O(N__27664),
            .I(N__27661));
    Odrv4 I__4316 (
            .O(N__27661),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ));
    CascadeMux I__4315 (
            .O(N__27658),
            .I(N__27655));
    InMux I__4314 (
            .O(N__27655),
            .I(N__27652));
    LocalMux I__4313 (
            .O(N__27652),
            .I(N__27649));
    Odrv4 I__4312 (
            .O(N__27649),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_25 ));
    InMux I__4311 (
            .O(N__27646),
            .I(N__27643));
    LocalMux I__4310 (
            .O(N__27643),
            .I(N__27639));
    InMux I__4309 (
            .O(N__27642),
            .I(N__27636));
    Span4Mux_v I__4308 (
            .O(N__27639),
            .I(N__27630));
    LocalMux I__4307 (
            .O(N__27636),
            .I(N__27630));
    InMux I__4306 (
            .O(N__27635),
            .I(N__27627));
    Span4Mux_v I__4305 (
            .O(N__27630),
            .I(N__27624));
    LocalMux I__4304 (
            .O(N__27627),
            .I(measured_delay_tr_5));
    Odrv4 I__4303 (
            .O(N__27624),
            .I(measured_delay_tr_5));
    CascadeMux I__4302 (
            .O(N__27619),
            .I(N__27616));
    InMux I__4301 (
            .O(N__27616),
            .I(N__27613));
    LocalMux I__4300 (
            .O(N__27613),
            .I(N__27610));
    Span4Mux_h I__4299 (
            .O(N__27610),
            .I(N__27607));
    Odrv4 I__4298 (
            .O(N__27607),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_19 ));
    InMux I__4297 (
            .O(N__27604),
            .I(N__27601));
    LocalMux I__4296 (
            .O(N__27601),
            .I(N__27598));
    Odrv12 I__4295 (
            .O(N__27598),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_17 ));
    CascadeMux I__4294 (
            .O(N__27595),
            .I(N__27592));
    InMux I__4293 (
            .O(N__27592),
            .I(N__27589));
    LocalMux I__4292 (
            .O(N__27589),
            .I(N__27586));
    Odrv12 I__4291 (
            .O(N__27586),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_20 ));
    CascadeMux I__4290 (
            .O(N__27583),
            .I(N__27580));
    InMux I__4289 (
            .O(N__27580),
            .I(N__27577));
    LocalMux I__4288 (
            .O(N__27577),
            .I(N__27574));
    Span4Mux_h I__4287 (
            .O(N__27574),
            .I(N__27571));
    Odrv4 I__4286 (
            .O(N__27571),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ));
    InMux I__4285 (
            .O(N__27568),
            .I(N__27563));
    CascadeMux I__4284 (
            .O(N__27567),
            .I(N__27559));
    InMux I__4283 (
            .O(N__27566),
            .I(N__27556));
    LocalMux I__4282 (
            .O(N__27563),
            .I(N__27553));
    InMux I__4281 (
            .O(N__27562),
            .I(N__27550));
    InMux I__4280 (
            .O(N__27559),
            .I(N__27547));
    LocalMux I__4279 (
            .O(N__27556),
            .I(N__27542));
    Span4Mux_v I__4278 (
            .O(N__27553),
            .I(N__27542));
    LocalMux I__4277 (
            .O(N__27550),
            .I(N__27539));
    LocalMux I__4276 (
            .O(N__27547),
            .I(N__27534));
    Span4Mux_v I__4275 (
            .O(N__27542),
            .I(N__27534));
    Span4Mux_v I__4274 (
            .O(N__27539),
            .I(N__27531));
    Odrv4 I__4273 (
            .O(N__27534),
            .I(measured_delay_tr_7));
    Odrv4 I__4272 (
            .O(N__27531),
            .I(measured_delay_tr_7));
    CascadeMux I__4271 (
            .O(N__27526),
            .I(N__27523));
    InMux I__4270 (
            .O(N__27523),
            .I(N__27520));
    LocalMux I__4269 (
            .O(N__27520),
            .I(N__27517));
    Odrv4 I__4268 (
            .O(N__27517),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_22 ));
    CascadeMux I__4267 (
            .O(N__27514),
            .I(N__27511));
    InMux I__4266 (
            .O(N__27511),
            .I(N__27508));
    LocalMux I__4265 (
            .O(N__27508),
            .I(N__27505));
    Odrv4 I__4264 (
            .O(N__27505),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_16 ));
    InMux I__4263 (
            .O(N__27502),
            .I(N__27498));
    InMux I__4262 (
            .O(N__27501),
            .I(N__27495));
    LocalMux I__4261 (
            .O(N__27498),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    LocalMux I__4260 (
            .O(N__27495),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    InMux I__4259 (
            .O(N__27490),
            .I(N__27487));
    LocalMux I__4258 (
            .O(N__27487),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16 ));
    InMux I__4257 (
            .O(N__27484),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ));
    InMux I__4256 (
            .O(N__27481),
            .I(N__27477));
    InMux I__4255 (
            .O(N__27480),
            .I(N__27474));
    LocalMux I__4254 (
            .O(N__27477),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    LocalMux I__4253 (
            .O(N__27474),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    InMux I__4252 (
            .O(N__27469),
            .I(N__27466));
    LocalMux I__4251 (
            .O(N__27466),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17 ));
    InMux I__4250 (
            .O(N__27463),
            .I(bfn_10_26_0_));
    InMux I__4249 (
            .O(N__27460),
            .I(N__27456));
    InMux I__4248 (
            .O(N__27459),
            .I(N__27453));
    LocalMux I__4247 (
            .O(N__27456),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    LocalMux I__4246 (
            .O(N__27453),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__4245 (
            .O(N__27448),
            .I(N__27445));
    LocalMux I__4244 (
            .O(N__27445),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18 ));
    InMux I__4243 (
            .O(N__27442),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ));
    InMux I__4242 (
            .O(N__27439),
            .I(N__27435));
    InMux I__4241 (
            .O(N__27438),
            .I(N__27432));
    LocalMux I__4240 (
            .O(N__27435),
            .I(N__27429));
    LocalMux I__4239 (
            .O(N__27432),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    Odrv4 I__4238 (
            .O(N__27429),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__4237 (
            .O(N__27424),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17 ));
    InMux I__4236 (
            .O(N__27421),
            .I(N__27418));
    LocalMux I__4235 (
            .O(N__27418),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19 ));
    InMux I__4234 (
            .O(N__27415),
            .I(N__27412));
    LocalMux I__4233 (
            .O(N__27412),
            .I(N__27409));
    Span12Mux_h I__4232 (
            .O(N__27409),
            .I(N__27406));
    Odrv12 I__4231 (
            .O(N__27406),
            .I(delay_hc_input_c));
    InMux I__4230 (
            .O(N__27403),
            .I(N__27400));
    LocalMux I__4229 (
            .O(N__27400),
            .I(delay_hc_d1));
    InMux I__4228 (
            .O(N__27397),
            .I(N__27394));
    LocalMux I__4227 (
            .O(N__27394),
            .I(N__27389));
    InMux I__4226 (
            .O(N__27393),
            .I(N__27386));
    InMux I__4225 (
            .O(N__27392),
            .I(N__27382));
    Span4Mux_h I__4224 (
            .O(N__27389),
            .I(N__27379));
    LocalMux I__4223 (
            .O(N__27386),
            .I(N__27376));
    InMux I__4222 (
            .O(N__27385),
            .I(N__27373));
    LocalMux I__4221 (
            .O(N__27382),
            .I(delay_hc_d2));
    Odrv4 I__4220 (
            .O(N__27379),
            .I(delay_hc_d2));
    Odrv4 I__4219 (
            .O(N__27376),
            .I(delay_hc_d2));
    LocalMux I__4218 (
            .O(N__27373),
            .I(delay_hc_d2));
    InMux I__4217 (
            .O(N__27364),
            .I(N__27360));
    InMux I__4216 (
            .O(N__27363),
            .I(N__27356));
    LocalMux I__4215 (
            .O(N__27360),
            .I(N__27353));
    InMux I__4214 (
            .O(N__27359),
            .I(N__27350));
    LocalMux I__4213 (
            .O(N__27356),
            .I(\delay_measurement_inst.prev_hc_sigZ0 ));
    Odrv4 I__4212 (
            .O(N__27353),
            .I(\delay_measurement_inst.prev_hc_sigZ0 ));
    LocalMux I__4211 (
            .O(N__27350),
            .I(\delay_measurement_inst.prev_hc_sigZ0 ));
    InMux I__4210 (
            .O(N__27343),
            .I(N__27339));
    InMux I__4209 (
            .O(N__27342),
            .I(N__27336));
    LocalMux I__4208 (
            .O(N__27339),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    LocalMux I__4207 (
            .O(N__27336),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    InMux I__4206 (
            .O(N__27331),
            .I(N__27328));
    LocalMux I__4205 (
            .O(N__27328),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8 ));
    InMux I__4204 (
            .O(N__27325),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ));
    InMux I__4203 (
            .O(N__27322),
            .I(N__27319));
    LocalMux I__4202 (
            .O(N__27319),
            .I(N__27315));
    InMux I__4201 (
            .O(N__27318),
            .I(N__27312));
    Odrv12 I__4200 (
            .O(N__27315),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    LocalMux I__4199 (
            .O(N__27312),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    InMux I__4198 (
            .O(N__27307),
            .I(N__27304));
    LocalMux I__4197 (
            .O(N__27304),
            .I(N__27301));
    Odrv4 I__4196 (
            .O(N__27301),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9 ));
    InMux I__4195 (
            .O(N__27298),
            .I(bfn_10_25_0_));
    InMux I__4194 (
            .O(N__27295),
            .I(N__27292));
    LocalMux I__4193 (
            .O(N__27292),
            .I(N__27288));
    InMux I__4192 (
            .O(N__27291),
            .I(N__27285));
    Odrv4 I__4191 (
            .O(N__27288),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    LocalMux I__4190 (
            .O(N__27285),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    InMux I__4189 (
            .O(N__27280),
            .I(N__27277));
    LocalMux I__4188 (
            .O(N__27277),
            .I(N__27274));
    Odrv4 I__4187 (
            .O(N__27274),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10 ));
    InMux I__4186 (
            .O(N__27271),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ));
    InMux I__4185 (
            .O(N__27268),
            .I(N__27264));
    InMux I__4184 (
            .O(N__27267),
            .I(N__27261));
    LocalMux I__4183 (
            .O(N__27264),
            .I(N__27258));
    LocalMux I__4182 (
            .O(N__27261),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    Odrv4 I__4181 (
            .O(N__27258),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    InMux I__4180 (
            .O(N__27253),
            .I(N__27250));
    LocalMux I__4179 (
            .O(N__27250),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11 ));
    InMux I__4178 (
            .O(N__27247),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ));
    InMux I__4177 (
            .O(N__27244),
            .I(N__27240));
    InMux I__4176 (
            .O(N__27243),
            .I(N__27237));
    LocalMux I__4175 (
            .O(N__27240),
            .I(N__27234));
    LocalMux I__4174 (
            .O(N__27237),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    Odrv4 I__4173 (
            .O(N__27234),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__4172 (
            .O(N__27229),
            .I(N__27226));
    LocalMux I__4171 (
            .O(N__27226),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12 ));
    InMux I__4170 (
            .O(N__27223),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ));
    InMux I__4169 (
            .O(N__27220),
            .I(N__27216));
    InMux I__4168 (
            .O(N__27219),
            .I(N__27213));
    LocalMux I__4167 (
            .O(N__27216),
            .I(N__27210));
    LocalMux I__4166 (
            .O(N__27213),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    Odrv4 I__4165 (
            .O(N__27210),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__4164 (
            .O(N__27205),
            .I(N__27202));
    LocalMux I__4163 (
            .O(N__27202),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13 ));
    InMux I__4162 (
            .O(N__27199),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ));
    InMux I__4161 (
            .O(N__27196),
            .I(N__27192));
    InMux I__4160 (
            .O(N__27195),
            .I(N__27189));
    LocalMux I__4159 (
            .O(N__27192),
            .I(N__27186));
    LocalMux I__4158 (
            .O(N__27189),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    Odrv4 I__4157 (
            .O(N__27186),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    InMux I__4156 (
            .O(N__27181),
            .I(N__27178));
    LocalMux I__4155 (
            .O(N__27178),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14 ));
    InMux I__4154 (
            .O(N__27175),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ));
    InMux I__4153 (
            .O(N__27172),
            .I(N__27168));
    InMux I__4152 (
            .O(N__27171),
            .I(N__27165));
    LocalMux I__4151 (
            .O(N__27168),
            .I(N__27162));
    LocalMux I__4150 (
            .O(N__27165),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    Odrv4 I__4149 (
            .O(N__27162),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__4148 (
            .O(N__27157),
            .I(N__27154));
    LocalMux I__4147 (
            .O(N__27154),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15 ));
    InMux I__4146 (
            .O(N__27151),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ));
    InMux I__4145 (
            .O(N__27148),
            .I(N__27145));
    LocalMux I__4144 (
            .O(N__27145),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0 ));
    CascadeMux I__4143 (
            .O(N__27142),
            .I(N__27138));
    CascadeMux I__4142 (
            .O(N__27141),
            .I(N__27135));
    InMux I__4141 (
            .O(N__27138),
            .I(N__27132));
    InMux I__4140 (
            .O(N__27135),
            .I(N__27129));
    LocalMux I__4139 (
            .O(N__27132),
            .I(N__27123));
    LocalMux I__4138 (
            .O(N__27129),
            .I(N__27123));
    InMux I__4137 (
            .O(N__27128),
            .I(N__27120));
    Odrv4 I__4136 (
            .O(N__27123),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__4135 (
            .O(N__27120),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    InMux I__4134 (
            .O(N__27115),
            .I(N__27111));
    InMux I__4133 (
            .O(N__27114),
            .I(N__27108));
    LocalMux I__4132 (
            .O(N__27111),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    LocalMux I__4131 (
            .O(N__27108),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    InMux I__4130 (
            .O(N__27103),
            .I(N__27100));
    LocalMux I__4129 (
            .O(N__27100),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2 ));
    InMux I__4128 (
            .O(N__27097),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ));
    InMux I__4127 (
            .O(N__27094),
            .I(N__27091));
    LocalMux I__4126 (
            .O(N__27091),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0 ));
    CascadeMux I__4125 (
            .O(N__27088),
            .I(N__27085));
    InMux I__4124 (
            .O(N__27085),
            .I(N__27081));
    InMux I__4123 (
            .O(N__27084),
            .I(N__27078));
    LocalMux I__4122 (
            .O(N__27081),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    LocalMux I__4121 (
            .O(N__27078),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    InMux I__4120 (
            .O(N__27073),
            .I(N__27070));
    LocalMux I__4119 (
            .O(N__27070),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3 ));
    InMux I__4118 (
            .O(N__27067),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ));
    InMux I__4117 (
            .O(N__27064),
            .I(N__27060));
    InMux I__4116 (
            .O(N__27063),
            .I(N__27057));
    LocalMux I__4115 (
            .O(N__27060),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    LocalMux I__4114 (
            .O(N__27057),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    InMux I__4113 (
            .O(N__27052),
            .I(N__27049));
    LocalMux I__4112 (
            .O(N__27049),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4 ));
    InMux I__4111 (
            .O(N__27046),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ));
    InMux I__4110 (
            .O(N__27043),
            .I(N__27039));
    InMux I__4109 (
            .O(N__27042),
            .I(N__27036));
    LocalMux I__4108 (
            .O(N__27039),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    LocalMux I__4107 (
            .O(N__27036),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    InMux I__4106 (
            .O(N__27031),
            .I(N__27028));
    LocalMux I__4105 (
            .O(N__27028),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5 ));
    InMux I__4104 (
            .O(N__27025),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ));
    InMux I__4103 (
            .O(N__27022),
            .I(N__27018));
    InMux I__4102 (
            .O(N__27021),
            .I(N__27015));
    LocalMux I__4101 (
            .O(N__27018),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    LocalMux I__4100 (
            .O(N__27015),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    InMux I__4099 (
            .O(N__27010),
            .I(N__27007));
    LocalMux I__4098 (
            .O(N__27007),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6 ));
    InMux I__4097 (
            .O(N__27004),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ));
    InMux I__4096 (
            .O(N__27001),
            .I(N__26997));
    InMux I__4095 (
            .O(N__27000),
            .I(N__26994));
    LocalMux I__4094 (
            .O(N__26997),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    LocalMux I__4093 (
            .O(N__26994),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    InMux I__4092 (
            .O(N__26989),
            .I(N__26986));
    LocalMux I__4091 (
            .O(N__26986),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7 ));
    InMux I__4090 (
            .O(N__26983),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ));
    CascadeMux I__4089 (
            .O(N__26980),
            .I(N__26977));
    InMux I__4088 (
            .O(N__26977),
            .I(N__26974));
    LocalMux I__4087 (
            .O(N__26974),
            .I(N__26971));
    Odrv12 I__4086 (
            .O(N__26971),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ));
    InMux I__4085 (
            .O(N__26968),
            .I(N__26965));
    LocalMux I__4084 (
            .O(N__26965),
            .I(N__26962));
    Span4Mux_h I__4083 (
            .O(N__26962),
            .I(N__26959));
    Odrv4 I__4082 (
            .O(N__26959),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0 ));
    CascadeMux I__4081 (
            .O(N__26956),
            .I(N__26953));
    InMux I__4080 (
            .O(N__26953),
            .I(N__26950));
    LocalMux I__4079 (
            .O(N__26950),
            .I(N__26947));
    Span4Mux_h I__4078 (
            .O(N__26947),
            .I(N__26944));
    Odrv4 I__4077 (
            .O(N__26944),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ1Z_6 ));
    CascadeMux I__4076 (
            .O(N__26941),
            .I(N__26938));
    InMux I__4075 (
            .O(N__26938),
            .I(N__26935));
    LocalMux I__4074 (
            .O(N__26935),
            .I(N__26932));
    Odrv4 I__4073 (
            .O(N__26932),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ));
    InMux I__4072 (
            .O(N__26929),
            .I(N__26926));
    LocalMux I__4071 (
            .O(N__26926),
            .I(N__26923));
    Span4Mux_h I__4070 (
            .O(N__26923),
            .I(N__26920));
    Odrv4 I__4069 (
            .O(N__26920),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_0 ));
    CascadeMux I__4068 (
            .O(N__26917),
            .I(N__26914));
    InMux I__4067 (
            .O(N__26914),
            .I(N__26911));
    LocalMux I__4066 (
            .O(N__26911),
            .I(N__26908));
    Odrv12 I__4065 (
            .O(N__26908),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ));
    CascadeMux I__4064 (
            .O(N__26905),
            .I(N__26902));
    InMux I__4063 (
            .O(N__26902),
            .I(N__26899));
    LocalMux I__4062 (
            .O(N__26899),
            .I(N__26896));
    Span4Mux_h I__4061 (
            .O(N__26896),
            .I(N__26893));
    Odrv4 I__4060 (
            .O(N__26893),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ));
    CascadeMux I__4059 (
            .O(N__26890),
            .I(N__26887));
    InMux I__4058 (
            .O(N__26887),
            .I(N__26884));
    LocalMux I__4057 (
            .O(N__26884),
            .I(N__26881));
    Span4Mux_v I__4056 (
            .O(N__26881),
            .I(N__26878));
    Odrv4 I__4055 (
            .O(N__26878),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ));
    InMux I__4054 (
            .O(N__26875),
            .I(N__26872));
    LocalMux I__4053 (
            .O(N__26872),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_19 ));
    InMux I__4052 (
            .O(N__26869),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ));
    InMux I__4051 (
            .O(N__26866),
            .I(N__26863));
    LocalMux I__4050 (
            .O(N__26863),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_axb_0 ));
    InMux I__4049 (
            .O(N__26860),
            .I(N__26857));
    LocalMux I__4048 (
            .O(N__26857),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ));
    InMux I__4047 (
            .O(N__26854),
            .I(N__26851));
    LocalMux I__4046 (
            .O(N__26851),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ));
    InMux I__4045 (
            .O(N__26848),
            .I(N__26845));
    LocalMux I__4044 (
            .O(N__26845),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ));
    InMux I__4043 (
            .O(N__26842),
            .I(N__26839));
    LocalMux I__4042 (
            .O(N__26839),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ));
    InMux I__4041 (
            .O(N__26836),
            .I(N__26833));
    LocalMux I__4040 (
            .O(N__26833),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ));
    InMux I__4039 (
            .O(N__26830),
            .I(N__26827));
    LocalMux I__4038 (
            .O(N__26827),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_16 ));
    InMux I__4037 (
            .O(N__26824),
            .I(N__26821));
    LocalMux I__4036 (
            .O(N__26821),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_17 ));
    InMux I__4035 (
            .O(N__26818),
            .I(N__26815));
    LocalMux I__4034 (
            .O(N__26815),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_18 ));
    InMux I__4033 (
            .O(N__26812),
            .I(N__26809));
    LocalMux I__4032 (
            .O(N__26809),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ));
    InMux I__4031 (
            .O(N__26806),
            .I(N__26803));
    LocalMux I__4030 (
            .O(N__26803),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ));
    InMux I__4029 (
            .O(N__26800),
            .I(N__26797));
    LocalMux I__4028 (
            .O(N__26797),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ));
    InMux I__4027 (
            .O(N__26794),
            .I(N__26791));
    LocalMux I__4026 (
            .O(N__26791),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ));
    InMux I__4025 (
            .O(N__26788),
            .I(N__26785));
    LocalMux I__4024 (
            .O(N__26785),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ));
    InMux I__4023 (
            .O(N__26782),
            .I(N__26779));
    LocalMux I__4022 (
            .O(N__26779),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ));
    InMux I__4021 (
            .O(N__26776),
            .I(N__26773));
    LocalMux I__4020 (
            .O(N__26773),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ));
    InMux I__4019 (
            .O(N__26770),
            .I(N__26767));
    LocalMux I__4018 (
            .O(N__26767),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ));
    CascadeMux I__4017 (
            .O(N__26764),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9_cascade_ ));
    CascadeMux I__4016 (
            .O(N__26761),
            .I(N__26756));
    CascadeMux I__4015 (
            .O(N__26760),
            .I(N__26751));
    InMux I__4014 (
            .O(N__26759),
            .I(N__26746));
    InMux I__4013 (
            .O(N__26756),
            .I(N__26733));
    InMux I__4012 (
            .O(N__26755),
            .I(N__26733));
    InMux I__4011 (
            .O(N__26754),
            .I(N__26733));
    InMux I__4010 (
            .O(N__26751),
            .I(N__26733));
    InMux I__4009 (
            .O(N__26750),
            .I(N__26733));
    InMux I__4008 (
            .O(N__26749),
            .I(N__26733));
    LocalMux I__4007 (
            .O(N__26746),
            .I(N__26725));
    LocalMux I__4006 (
            .O(N__26733),
            .I(N__26722));
    InMux I__4005 (
            .O(N__26732),
            .I(N__26719));
    InMux I__4004 (
            .O(N__26731),
            .I(N__26706));
    InMux I__4003 (
            .O(N__26730),
            .I(N__26706));
    InMux I__4002 (
            .O(N__26729),
            .I(N__26706));
    InMux I__4001 (
            .O(N__26728),
            .I(N__26706));
    Span4Mux_v I__4000 (
            .O(N__26725),
            .I(N__26699));
    Span4Mux_h I__3999 (
            .O(N__26722),
            .I(N__26699));
    LocalMux I__3998 (
            .O(N__26719),
            .I(N__26699));
    InMux I__3997 (
            .O(N__26718),
            .I(N__26690));
    InMux I__3996 (
            .O(N__26717),
            .I(N__26690));
    InMux I__3995 (
            .O(N__26716),
            .I(N__26690));
    InMux I__3994 (
            .O(N__26715),
            .I(N__26690));
    LocalMux I__3993 (
            .O(N__26706),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6 ));
    Odrv4 I__3992 (
            .O(N__26699),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6 ));
    LocalMux I__3991 (
            .O(N__26690),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6 ));
    CascadeMux I__3990 (
            .O(N__26683),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6_cascade_ ));
    InMux I__3989 (
            .O(N__26680),
            .I(N__26677));
    LocalMux I__3988 (
            .O(N__26677),
            .I(N__26667));
    InMux I__3987 (
            .O(N__26676),
            .I(N__26658));
    InMux I__3986 (
            .O(N__26675),
            .I(N__26658));
    InMux I__3985 (
            .O(N__26674),
            .I(N__26658));
    InMux I__3984 (
            .O(N__26673),
            .I(N__26658));
    InMux I__3983 (
            .O(N__26672),
            .I(N__26655));
    CascadeMux I__3982 (
            .O(N__26671),
            .I(N__26652));
    CascadeMux I__3981 (
            .O(N__26670),
            .I(N__26649));
    Span4Mux_h I__3980 (
            .O(N__26667),
            .I(N__26641));
    LocalMux I__3979 (
            .O(N__26658),
            .I(N__26641));
    LocalMux I__3978 (
            .O(N__26655),
            .I(N__26641));
    InMux I__3977 (
            .O(N__26652),
            .I(N__26631));
    InMux I__3976 (
            .O(N__26649),
            .I(N__26631));
    InMux I__3975 (
            .O(N__26648),
            .I(N__26631));
    Span4Mux_v I__3974 (
            .O(N__26641),
            .I(N__26628));
    InMux I__3973 (
            .O(N__26640),
            .I(N__26621));
    InMux I__3972 (
            .O(N__26639),
            .I(N__26621));
    InMux I__3971 (
            .O(N__26638),
            .I(N__26621));
    LocalMux I__3970 (
            .O(N__26631),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6 ));
    Odrv4 I__3969 (
            .O(N__26628),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6 ));
    LocalMux I__3968 (
            .O(N__26621),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6 ));
    InMux I__3967 (
            .O(N__26614),
            .I(N__26611));
    LocalMux I__3966 (
            .O(N__26611),
            .I(N__26608));
    Span4Mux_h I__3965 (
            .O(N__26608),
            .I(N__26605));
    Odrv4 I__3964 (
            .O(N__26605),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3Z0Z_3 ));
    InMux I__3963 (
            .O(N__26602),
            .I(N__26599));
    LocalMux I__3962 (
            .O(N__26599),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6 ));
    CascadeMux I__3961 (
            .O(N__26596),
            .I(N__26593));
    InMux I__3960 (
            .O(N__26593),
            .I(N__26590));
    LocalMux I__3959 (
            .O(N__26590),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4Z0Z_3 ));
    InMux I__3958 (
            .O(N__26587),
            .I(N__26584));
    LocalMux I__3957 (
            .O(N__26584),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9 ));
    InMux I__3956 (
            .O(N__26581),
            .I(N__26578));
    LocalMux I__3955 (
            .O(N__26578),
            .I(N__26574));
    InMux I__3954 (
            .O(N__26577),
            .I(N__26571));
    Odrv4 I__3953 (
            .O(N__26574),
            .I(\phase_controller_inst1.stoper_tr.N_248 ));
    LocalMux I__3952 (
            .O(N__26571),
            .I(\phase_controller_inst1.stoper_tr.N_248 ));
    CascadeMux I__3951 (
            .O(N__26566),
            .I(\phase_controller_inst1.stoper_tr.N_248_cascade_ ));
    InMux I__3950 (
            .O(N__26563),
            .I(N__26557));
    InMux I__3949 (
            .O(N__26562),
            .I(N__26557));
    LocalMux I__3948 (
            .O(N__26557),
            .I(N__26552));
    InMux I__3947 (
            .O(N__26556),
            .I(N__26547));
    InMux I__3946 (
            .O(N__26555),
            .I(N__26547));
    Odrv12 I__3945 (
            .O(N__26552),
            .I(\phase_controller_inst1.stoper_tr.N_55 ));
    LocalMux I__3944 (
            .O(N__26547),
            .I(\phase_controller_inst1.stoper_tr.N_55 ));
    InMux I__3943 (
            .O(N__26542),
            .I(N__26539));
    LocalMux I__3942 (
            .O(N__26539),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ));
    InMux I__3941 (
            .O(N__26536),
            .I(N__26533));
    LocalMux I__3940 (
            .O(N__26533),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ));
    CascadeMux I__3939 (
            .O(N__26530),
            .I(N__26527));
    InMux I__3938 (
            .O(N__26527),
            .I(N__26524));
    LocalMux I__3937 (
            .O(N__26524),
            .I(N__26521));
    Odrv4 I__3936 (
            .O(N__26521),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ));
    CascadeMux I__3935 (
            .O(N__26518),
            .I(N__26515));
    InMux I__3934 (
            .O(N__26515),
            .I(N__26512));
    LocalMux I__3933 (
            .O(N__26512),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ));
    CascadeMux I__3932 (
            .O(N__26509),
            .I(N__26506));
    InMux I__3931 (
            .O(N__26506),
            .I(N__26503));
    LocalMux I__3930 (
            .O(N__26503),
            .I(N__26500));
    Odrv4 I__3929 (
            .O(N__26500),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ));
    CascadeMux I__3928 (
            .O(N__26497),
            .I(N__26494));
    InMux I__3927 (
            .O(N__26494),
            .I(N__26491));
    LocalMux I__3926 (
            .O(N__26491),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ));
    CascadeMux I__3925 (
            .O(N__26488),
            .I(N__26485));
    InMux I__3924 (
            .O(N__26485),
            .I(N__26482));
    LocalMux I__3923 (
            .O(N__26482),
            .I(N__26479));
    Odrv4 I__3922 (
            .O(N__26479),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ));
    CascadeMux I__3921 (
            .O(N__26476),
            .I(N__26473));
    InMux I__3920 (
            .O(N__26473),
            .I(N__26470));
    LocalMux I__3919 (
            .O(N__26470),
            .I(N__26467));
    Odrv4 I__3918 (
            .O(N__26467),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ));
    InMux I__3917 (
            .O(N__26464),
            .I(N__26461));
    LocalMux I__3916 (
            .O(N__26461),
            .I(N__26454));
    InMux I__3915 (
            .O(N__26460),
            .I(N__26447));
    InMux I__3914 (
            .O(N__26459),
            .I(N__26447));
    InMux I__3913 (
            .O(N__26458),
            .I(N__26447));
    CascadeMux I__3912 (
            .O(N__26457),
            .I(N__26443));
    Span4Mux_h I__3911 (
            .O(N__26454),
            .I(N__26436));
    LocalMux I__3910 (
            .O(N__26447),
            .I(N__26433));
    InMux I__3909 (
            .O(N__26446),
            .I(N__26430));
    InMux I__3908 (
            .O(N__26443),
            .I(N__26419));
    InMux I__3907 (
            .O(N__26442),
            .I(N__26419));
    InMux I__3906 (
            .O(N__26441),
            .I(N__26419));
    InMux I__3905 (
            .O(N__26440),
            .I(N__26419));
    InMux I__3904 (
            .O(N__26439),
            .I(N__26419));
    Odrv4 I__3903 (
            .O(N__26436),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9 ));
    Odrv4 I__3902 (
            .O(N__26433),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9 ));
    LocalMux I__3901 (
            .O(N__26430),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9 ));
    LocalMux I__3900 (
            .O(N__26419),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9 ));
    CascadeMux I__3899 (
            .O(N__26410),
            .I(N__26407));
    InMux I__3898 (
            .O(N__26407),
            .I(N__26404));
    LocalMux I__3897 (
            .O(N__26404),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ));
    InMux I__3896 (
            .O(N__26401),
            .I(N__26397));
    InMux I__3895 (
            .O(N__26400),
            .I(N__26394));
    LocalMux I__3894 (
            .O(N__26397),
            .I(N__26389));
    LocalMux I__3893 (
            .O(N__26394),
            .I(N__26389));
    Odrv12 I__3892 (
            .O(N__26389),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    InMux I__3891 (
            .O(N__26386),
            .I(N__26381));
    InMux I__3890 (
            .O(N__26385),
            .I(N__26378));
    InMux I__3889 (
            .O(N__26384),
            .I(N__26375));
    LocalMux I__3888 (
            .O(N__26381),
            .I(N__26372));
    LocalMux I__3887 (
            .O(N__26378),
            .I(N__26367));
    LocalMux I__3886 (
            .O(N__26375),
            .I(N__26367));
    Span4Mux_h I__3885 (
            .O(N__26372),
            .I(N__26364));
    Span4Mux_v I__3884 (
            .O(N__26367),
            .I(N__26361));
    Span4Mux_v I__3883 (
            .O(N__26364),
            .I(N__26358));
    Odrv4 I__3882 (
            .O(N__26361),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    Odrv4 I__3881 (
            .O(N__26358),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    CascadeMux I__3880 (
            .O(N__26353),
            .I(N__26350));
    InMux I__3879 (
            .O(N__26350),
            .I(N__26347));
    LocalMux I__3878 (
            .O(N__26347),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ));
    CascadeMux I__3877 (
            .O(N__26344),
            .I(N__26341));
    InMux I__3876 (
            .O(N__26341),
            .I(N__26338));
    LocalMux I__3875 (
            .O(N__26338),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ));
    CascadeMux I__3874 (
            .O(N__26335),
            .I(N__26332));
    InMux I__3873 (
            .O(N__26332),
            .I(N__26329));
    LocalMux I__3872 (
            .O(N__26329),
            .I(N__26326));
    Odrv4 I__3871 (
            .O(N__26326),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ));
    CascadeMux I__3870 (
            .O(N__26323),
            .I(N__26320));
    InMux I__3869 (
            .O(N__26320),
            .I(N__26317));
    LocalMux I__3868 (
            .O(N__26317),
            .I(N__26314));
    Odrv4 I__3867 (
            .O(N__26314),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ));
    CascadeMux I__3866 (
            .O(N__26311),
            .I(N__26308));
    InMux I__3865 (
            .O(N__26308),
            .I(N__26305));
    LocalMux I__3864 (
            .O(N__26305),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ));
    CascadeMux I__3863 (
            .O(N__26302),
            .I(N__26299));
    InMux I__3862 (
            .O(N__26299),
            .I(N__26296));
    LocalMux I__3861 (
            .O(N__26296),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ));
    CascadeMux I__3860 (
            .O(N__26293),
            .I(N__26290));
    InMux I__3859 (
            .O(N__26290),
            .I(N__26287));
    LocalMux I__3858 (
            .O(N__26287),
            .I(N__26284));
    Odrv4 I__3857 (
            .O(N__26284),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ));
    CascadeMux I__3856 (
            .O(N__26281),
            .I(N__26278));
    InMux I__3855 (
            .O(N__26278),
            .I(N__26275));
    LocalMux I__3854 (
            .O(N__26275),
            .I(N__26272));
    Odrv4 I__3853 (
            .O(N__26272),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ));
    CascadeMux I__3852 (
            .O(N__26269),
            .I(N__26266));
    InMux I__3851 (
            .O(N__26266),
            .I(N__26263));
    LocalMux I__3850 (
            .O(N__26263),
            .I(N__26260));
    Odrv4 I__3849 (
            .O(N__26260),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ));
    CascadeMux I__3848 (
            .O(N__26257),
            .I(N__26254));
    InMux I__3847 (
            .O(N__26254),
            .I(N__26251));
    LocalMux I__3846 (
            .O(N__26251),
            .I(N__26248));
    Odrv4 I__3845 (
            .O(N__26248),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ));
    CascadeMux I__3844 (
            .O(N__26245),
            .I(N__26242));
    InMux I__3843 (
            .O(N__26242),
            .I(N__26239));
    LocalMux I__3842 (
            .O(N__26239),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ));
    CascadeMux I__3841 (
            .O(N__26236),
            .I(N__26233));
    InMux I__3840 (
            .O(N__26233),
            .I(N__26230));
    LocalMux I__3839 (
            .O(N__26230),
            .I(N__26227));
    Odrv4 I__3838 (
            .O(N__26227),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ));
    InMux I__3837 (
            .O(N__26224),
            .I(N__26221));
    LocalMux I__3836 (
            .O(N__26221),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_23 ));
    CascadeMux I__3835 (
            .O(N__26218),
            .I(N__26212));
    CascadeMux I__3834 (
            .O(N__26217),
            .I(N__26208));
    CascadeMux I__3833 (
            .O(N__26216),
            .I(N__26204));
    InMux I__3832 (
            .O(N__26215),
            .I(N__26191));
    InMux I__3831 (
            .O(N__26212),
            .I(N__26191));
    InMux I__3830 (
            .O(N__26211),
            .I(N__26191));
    InMux I__3829 (
            .O(N__26208),
            .I(N__26191));
    InMux I__3828 (
            .O(N__26207),
            .I(N__26191));
    InMux I__3827 (
            .O(N__26204),
            .I(N__26191));
    LocalMux I__3826 (
            .O(N__26191),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_26 ));
    CascadeMux I__3825 (
            .O(N__26188),
            .I(N__26185));
    InMux I__3824 (
            .O(N__26185),
            .I(N__26182));
    LocalMux I__3823 (
            .O(N__26182),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ));
    InMux I__3822 (
            .O(N__26179),
            .I(N__26174));
    InMux I__3821 (
            .O(N__26178),
            .I(N__26171));
    InMux I__3820 (
            .O(N__26177),
            .I(N__26168));
    LocalMux I__3819 (
            .O(N__26174),
            .I(\delay_measurement_inst.hc_stateZ0Z_0 ));
    LocalMux I__3818 (
            .O(N__26171),
            .I(\delay_measurement_inst.hc_stateZ0Z_0 ));
    LocalMux I__3817 (
            .O(N__26168),
            .I(\delay_measurement_inst.hc_stateZ0Z_0 ));
    CascadeMux I__3816 (
            .O(N__26161),
            .I(N__26158));
    InMux I__3815 (
            .O(N__26158),
            .I(N__26155));
    LocalMux I__3814 (
            .O(N__26155),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ));
    InMux I__3813 (
            .O(N__26152),
            .I(N__26149));
    LocalMux I__3812 (
            .O(N__26149),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ));
    CascadeMux I__3811 (
            .O(N__26146),
            .I(N__26143));
    InMux I__3810 (
            .O(N__26143),
            .I(N__26140));
    LocalMux I__3809 (
            .O(N__26140),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ));
    CascadeMux I__3808 (
            .O(N__26137),
            .I(N__26134));
    InMux I__3807 (
            .O(N__26134),
            .I(N__26131));
    LocalMux I__3806 (
            .O(N__26131),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ));
    InMux I__3805 (
            .O(N__26128),
            .I(N__26125));
    LocalMux I__3804 (
            .O(N__26125),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ));
    InMux I__3803 (
            .O(N__26122),
            .I(N__26119));
    LocalMux I__3802 (
            .O(N__26119),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_15 ));
    CascadeMux I__3801 (
            .O(N__26116),
            .I(N__26113));
    InMux I__3800 (
            .O(N__26113),
            .I(N__26110));
    LocalMux I__3799 (
            .O(N__26110),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_18 ));
    InMux I__3798 (
            .O(N__26107),
            .I(N__26104));
    LocalMux I__3797 (
            .O(N__26104),
            .I(N__26100));
    CascadeMux I__3796 (
            .O(N__26103),
            .I(N__26097));
    Span4Mux_v I__3795 (
            .O(N__26100),
            .I(N__26092));
    InMux I__3794 (
            .O(N__26097),
            .I(N__26087));
    InMux I__3793 (
            .O(N__26096),
            .I(N__26087));
    InMux I__3792 (
            .O(N__26095),
            .I(N__26084));
    Span4Mux_v I__3791 (
            .O(N__26092),
            .I(N__26079));
    LocalMux I__3790 (
            .O(N__26087),
            .I(N__26079));
    LocalMux I__3789 (
            .O(N__26084),
            .I(N__26074));
    Span4Mux_v I__3788 (
            .O(N__26079),
            .I(N__26074));
    Odrv4 I__3787 (
            .O(N__26074),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    IoInMux I__3786 (
            .O(N__26071),
            .I(N__26068));
    LocalMux I__3785 (
            .O(N__26068),
            .I(N__26065));
    Odrv12 I__3784 (
            .O(N__26065),
            .I(s3_phy_c));
    CascadeMux I__3783 (
            .O(N__26062),
            .I(N__26058));
    InMux I__3782 (
            .O(N__26061),
            .I(N__26055));
    InMux I__3781 (
            .O(N__26058),
            .I(N__26052));
    LocalMux I__3780 (
            .O(N__26055),
            .I(N__26048));
    LocalMux I__3779 (
            .O(N__26052),
            .I(N__26045));
    CascadeMux I__3778 (
            .O(N__26051),
            .I(N__26042));
    Span12Mux_v I__3777 (
            .O(N__26048),
            .I(N__26038));
    Span4Mux_v I__3776 (
            .O(N__26045),
            .I(N__26035));
    InMux I__3775 (
            .O(N__26042),
            .I(N__26032));
    InMux I__3774 (
            .O(N__26041),
            .I(N__26029));
    Odrv12 I__3773 (
            .O(N__26038),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv4 I__3772 (
            .O(N__26035),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    LocalMux I__3771 (
            .O(N__26032),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    LocalMux I__3770 (
            .O(N__26029),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    IoInMux I__3769 (
            .O(N__26020),
            .I(N__26017));
    LocalMux I__3768 (
            .O(N__26017),
            .I(N__26014));
    Span4Mux_s1_v I__3767 (
            .O(N__26014),
            .I(N__26011));
    Span4Mux_h I__3766 (
            .O(N__26011),
            .I(N__26008));
    Odrv4 I__3765 (
            .O(N__26008),
            .I(s2_phy_c));
    InMux I__3764 (
            .O(N__26005),
            .I(N__26002));
    LocalMux I__3763 (
            .O(N__26002),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_17 ));
    InMux I__3762 (
            .O(N__25999),
            .I(N__25996));
    LocalMux I__3761 (
            .O(N__25996),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_18 ));
    InMux I__3760 (
            .O(N__25993),
            .I(N__25990));
    LocalMux I__3759 (
            .O(N__25990),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_19 ));
    InMux I__3758 (
            .O(N__25987),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ));
    InMux I__3757 (
            .O(N__25984),
            .I(N__25978));
    InMux I__3756 (
            .O(N__25983),
            .I(N__25978));
    LocalMux I__3755 (
            .O(N__25978),
            .I(N__25971));
    InMux I__3754 (
            .O(N__25977),
            .I(N__25968));
    InMux I__3753 (
            .O(N__25976),
            .I(N__25961));
    InMux I__3752 (
            .O(N__25975),
            .I(N__25961));
    InMux I__3751 (
            .O(N__25974),
            .I(N__25961));
    Odrv12 I__3750 (
            .O(N__25971),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__3749 (
            .O(N__25968),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__3748 (
            .O(N__25961),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    InMux I__3747 (
            .O(N__25954),
            .I(N__25951));
    LocalMux I__3746 (
            .O(N__25951),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ));
    InMux I__3745 (
            .O(N__25948),
            .I(N__25945));
    LocalMux I__3744 (
            .O(N__25945),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ));
    InMux I__3743 (
            .O(N__25942),
            .I(N__25939));
    LocalMux I__3742 (
            .O(N__25939),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ));
    InMux I__3741 (
            .O(N__25936),
            .I(N__25933));
    LocalMux I__3740 (
            .O(N__25933),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ));
    InMux I__3739 (
            .O(N__25930),
            .I(N__25927));
    LocalMux I__3738 (
            .O(N__25927),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ));
    InMux I__3737 (
            .O(N__25924),
            .I(N__25921));
    LocalMux I__3736 (
            .O(N__25921),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ));
    InMux I__3735 (
            .O(N__25918),
            .I(N__25915));
    LocalMux I__3734 (
            .O(N__25915),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ));
    InMux I__3733 (
            .O(N__25912),
            .I(N__25909));
    LocalMux I__3732 (
            .O(N__25909),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_16 ));
    CascadeMux I__3731 (
            .O(N__25906),
            .I(N__25903));
    InMux I__3730 (
            .O(N__25903),
            .I(N__25900));
    LocalMux I__3729 (
            .O(N__25900),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ));
    InMux I__3728 (
            .O(N__25897),
            .I(N__25894));
    LocalMux I__3727 (
            .O(N__25894),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ));
    CascadeMux I__3726 (
            .O(N__25891),
            .I(N__25888));
    InMux I__3725 (
            .O(N__25888),
            .I(N__25885));
    LocalMux I__3724 (
            .O(N__25885),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ));
    InMux I__3723 (
            .O(N__25882),
            .I(N__25879));
    LocalMux I__3722 (
            .O(N__25879),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ));
    InMux I__3721 (
            .O(N__25876),
            .I(N__25873));
    LocalMux I__3720 (
            .O(N__25873),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ));
    CascadeMux I__3719 (
            .O(N__25870),
            .I(N__25867));
    InMux I__3718 (
            .O(N__25867),
            .I(N__25864));
    LocalMux I__3717 (
            .O(N__25864),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ));
    InMux I__3716 (
            .O(N__25861),
            .I(N__25858));
    LocalMux I__3715 (
            .O(N__25858),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ));
    CascadeMux I__3714 (
            .O(N__25855),
            .I(N__25852));
    InMux I__3713 (
            .O(N__25852),
            .I(N__25849));
    LocalMux I__3712 (
            .O(N__25849),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ));
    InMux I__3711 (
            .O(N__25846),
            .I(N__25843));
    LocalMux I__3710 (
            .O(N__25843),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ));
    InMux I__3709 (
            .O(N__25840),
            .I(N__25837));
    LocalMux I__3708 (
            .O(N__25837),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ));
    InMux I__3707 (
            .O(N__25834),
            .I(N__25831));
    LocalMux I__3706 (
            .O(N__25831),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ));
    InMux I__3705 (
            .O(N__25828),
            .I(N__25825));
    LocalMux I__3704 (
            .O(N__25825),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ));
    InMux I__3703 (
            .O(N__25822),
            .I(N__25819));
    LocalMux I__3702 (
            .O(N__25819),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0 ));
    InMux I__3701 (
            .O(N__25816),
            .I(N__25809));
    InMux I__3700 (
            .O(N__25815),
            .I(N__25809));
    InMux I__3699 (
            .O(N__25814),
            .I(N__25803));
    LocalMux I__3698 (
            .O(N__25809),
            .I(N__25800));
    InMux I__3697 (
            .O(N__25808),
            .I(N__25797));
    InMux I__3696 (
            .O(N__25807),
            .I(N__25792));
    InMux I__3695 (
            .O(N__25806),
            .I(N__25792));
    LocalMux I__3694 (
            .O(N__25803),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__3693 (
            .O(N__25800),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__3692 (
            .O(N__25797),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__3691 (
            .O(N__25792),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    InMux I__3690 (
            .O(N__25783),
            .I(N__25779));
    CascadeMux I__3689 (
            .O(N__25782),
            .I(N__25775));
    LocalMux I__3688 (
            .O(N__25779),
            .I(N__25771));
    InMux I__3687 (
            .O(N__25778),
            .I(N__25768));
    InMux I__3686 (
            .O(N__25775),
            .I(N__25763));
    InMux I__3685 (
            .O(N__25774),
            .I(N__25763));
    Span4Mux_h I__3684 (
            .O(N__25771),
            .I(N__25758));
    LocalMux I__3683 (
            .O(N__25768),
            .I(N__25758));
    LocalMux I__3682 (
            .O(N__25763),
            .I(N__25755));
    Odrv4 I__3681 (
            .O(N__25758),
            .I(\phase_controller_inst1.stoper_tr.time_passed11 ));
    Odrv4 I__3680 (
            .O(N__25755),
            .I(\phase_controller_inst1.stoper_tr.time_passed11 ));
    InMux I__3679 (
            .O(N__25750),
            .I(N__25747));
    LocalMux I__3678 (
            .O(N__25747),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0 ));
    InMux I__3677 (
            .O(N__25744),
            .I(N__25741));
    LocalMux I__3676 (
            .O(N__25741),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_0 ));
    InMux I__3675 (
            .O(N__25738),
            .I(N__25734));
    InMux I__3674 (
            .O(N__25737),
            .I(N__25731));
    LocalMux I__3673 (
            .O(N__25734),
            .I(N__25725));
    LocalMux I__3672 (
            .O(N__25731),
            .I(N__25725));
    InMux I__3671 (
            .O(N__25730),
            .I(N__25722));
    Span4Mux_h I__3670 (
            .O(N__25725),
            .I(N__25719));
    LocalMux I__3669 (
            .O(N__25722),
            .I(N__25714));
    Sp12to4 I__3668 (
            .O(N__25719),
            .I(N__25714));
    Odrv12 I__3667 (
            .O(N__25714),
            .I(il_max_comp2_D2));
    InMux I__3666 (
            .O(N__25711),
            .I(N__25708));
    LocalMux I__3665 (
            .O(N__25708),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7 ));
    InMux I__3664 (
            .O(N__25705),
            .I(N__25701));
    InMux I__3663 (
            .O(N__25704),
            .I(N__25698));
    LocalMux I__3662 (
            .O(N__25701),
            .I(N__25695));
    LocalMux I__3661 (
            .O(N__25698),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    Odrv4 I__3660 (
            .O(N__25695),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    CascadeMux I__3659 (
            .O(N__25690),
            .I(N__25687));
    InMux I__3658 (
            .O(N__25687),
            .I(N__25684));
    LocalMux I__3657 (
            .O(N__25684),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8 ));
    CascadeMux I__3656 (
            .O(N__25681),
            .I(N__25677));
    InMux I__3655 (
            .O(N__25680),
            .I(N__25674));
    InMux I__3654 (
            .O(N__25677),
            .I(N__25671));
    LocalMux I__3653 (
            .O(N__25674),
            .I(N__25668));
    LocalMux I__3652 (
            .O(N__25671),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    Odrv4 I__3651 (
            .O(N__25668),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__3650 (
            .O(N__25663),
            .I(N__25645));
    InMux I__3649 (
            .O(N__25662),
            .I(N__25645));
    InMux I__3648 (
            .O(N__25661),
            .I(N__25645));
    CascadeMux I__3647 (
            .O(N__25660),
            .I(N__25634));
    InMux I__3646 (
            .O(N__25659),
            .I(N__25626));
    InMux I__3645 (
            .O(N__25658),
            .I(N__25626));
    InMux I__3644 (
            .O(N__25657),
            .I(N__25613));
    InMux I__3643 (
            .O(N__25656),
            .I(N__25613));
    InMux I__3642 (
            .O(N__25655),
            .I(N__25613));
    InMux I__3641 (
            .O(N__25654),
            .I(N__25613));
    InMux I__3640 (
            .O(N__25653),
            .I(N__25613));
    InMux I__3639 (
            .O(N__25652),
            .I(N__25613));
    LocalMux I__3638 (
            .O(N__25645),
            .I(N__25610));
    InMux I__3637 (
            .O(N__25644),
            .I(N__25593));
    InMux I__3636 (
            .O(N__25643),
            .I(N__25593));
    InMux I__3635 (
            .O(N__25642),
            .I(N__25593));
    InMux I__3634 (
            .O(N__25641),
            .I(N__25593));
    InMux I__3633 (
            .O(N__25640),
            .I(N__25593));
    InMux I__3632 (
            .O(N__25639),
            .I(N__25593));
    InMux I__3631 (
            .O(N__25638),
            .I(N__25593));
    InMux I__3630 (
            .O(N__25637),
            .I(N__25593));
    InMux I__3629 (
            .O(N__25634),
            .I(N__25588));
    InMux I__3628 (
            .O(N__25633),
            .I(N__25588));
    InMux I__3627 (
            .O(N__25632),
            .I(N__25582));
    InMux I__3626 (
            .O(N__25631),
            .I(N__25582));
    LocalMux I__3625 (
            .O(N__25626),
            .I(N__25577));
    LocalMux I__3624 (
            .O(N__25613),
            .I(N__25577));
    Span4Mux_v I__3623 (
            .O(N__25610),
            .I(N__25574));
    LocalMux I__3622 (
            .O(N__25593),
            .I(N__25569));
    LocalMux I__3621 (
            .O(N__25588),
            .I(N__25569));
    InMux I__3620 (
            .O(N__25587),
            .I(N__25566));
    LocalMux I__3619 (
            .O(N__25582),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__3618 (
            .O(N__25577),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__3617 (
            .O(N__25574),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv12 I__3616 (
            .O(N__25569),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    LocalMux I__3615 (
            .O(N__25566),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    CascadeMux I__3614 (
            .O(N__25555),
            .I(N__25544));
    CascadeMux I__3613 (
            .O(N__25554),
            .I(N__25541));
    CascadeMux I__3612 (
            .O(N__25553),
            .I(N__25538));
    CascadeMux I__3611 (
            .O(N__25552),
            .I(N__25535));
    InMux I__3610 (
            .O(N__25551),
            .I(N__25524));
    InMux I__3609 (
            .O(N__25550),
            .I(N__25524));
    InMux I__3608 (
            .O(N__25549),
            .I(N__25517));
    InMux I__3607 (
            .O(N__25548),
            .I(N__25517));
    InMux I__3606 (
            .O(N__25547),
            .I(N__25517));
    InMux I__3605 (
            .O(N__25544),
            .I(N__25500));
    InMux I__3604 (
            .O(N__25541),
            .I(N__25500));
    InMux I__3603 (
            .O(N__25538),
            .I(N__25500));
    InMux I__3602 (
            .O(N__25535),
            .I(N__25500));
    InMux I__3601 (
            .O(N__25534),
            .I(N__25487));
    InMux I__3600 (
            .O(N__25533),
            .I(N__25487));
    InMux I__3599 (
            .O(N__25532),
            .I(N__25487));
    InMux I__3598 (
            .O(N__25531),
            .I(N__25487));
    InMux I__3597 (
            .O(N__25530),
            .I(N__25487));
    InMux I__3596 (
            .O(N__25529),
            .I(N__25487));
    LocalMux I__3595 (
            .O(N__25524),
            .I(N__25482));
    LocalMux I__3594 (
            .O(N__25517),
            .I(N__25482));
    InMux I__3593 (
            .O(N__25516),
            .I(N__25477));
    InMux I__3592 (
            .O(N__25515),
            .I(N__25477));
    InMux I__3591 (
            .O(N__25514),
            .I(N__25471));
    InMux I__3590 (
            .O(N__25513),
            .I(N__25471));
    InMux I__3589 (
            .O(N__25512),
            .I(N__25462));
    InMux I__3588 (
            .O(N__25511),
            .I(N__25462));
    InMux I__3587 (
            .O(N__25510),
            .I(N__25462));
    InMux I__3586 (
            .O(N__25509),
            .I(N__25462));
    LocalMux I__3585 (
            .O(N__25500),
            .I(N__25455));
    LocalMux I__3584 (
            .O(N__25487),
            .I(N__25455));
    Span4Mux_h I__3583 (
            .O(N__25482),
            .I(N__25455));
    LocalMux I__3582 (
            .O(N__25477),
            .I(N__25452));
    InMux I__3581 (
            .O(N__25476),
            .I(N__25449));
    LocalMux I__3580 (
            .O(N__25471),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    LocalMux I__3579 (
            .O(N__25462),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__3578 (
            .O(N__25455),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv12 I__3577 (
            .O(N__25452),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    LocalMux I__3576 (
            .O(N__25449),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    CascadeMux I__3575 (
            .O(N__25438),
            .I(N__25424));
    CascadeMux I__3574 (
            .O(N__25437),
            .I(N__25421));
    CascadeMux I__3573 (
            .O(N__25436),
            .I(N__25414));
    CascadeMux I__3572 (
            .O(N__25435),
            .I(N__25411));
    CascadeMux I__3571 (
            .O(N__25434),
            .I(N__25408));
    CascadeMux I__3570 (
            .O(N__25433),
            .I(N__25405));
    CascadeMux I__3569 (
            .O(N__25432),
            .I(N__25402));
    CascadeMux I__3568 (
            .O(N__25431),
            .I(N__25399));
    CascadeMux I__3567 (
            .O(N__25430),
            .I(N__25396));
    CascadeMux I__3566 (
            .O(N__25429),
            .I(N__25393));
    CascadeMux I__3565 (
            .O(N__25428),
            .I(N__25390));
    CascadeMux I__3564 (
            .O(N__25427),
            .I(N__25382));
    InMux I__3563 (
            .O(N__25424),
            .I(N__25375));
    InMux I__3562 (
            .O(N__25421),
            .I(N__25375));
    InMux I__3561 (
            .O(N__25420),
            .I(N__25375));
    InMux I__3560 (
            .O(N__25419),
            .I(N__25360));
    InMux I__3559 (
            .O(N__25418),
            .I(N__25360));
    InMux I__3558 (
            .O(N__25417),
            .I(N__25360));
    InMux I__3557 (
            .O(N__25414),
            .I(N__25360));
    InMux I__3556 (
            .O(N__25411),
            .I(N__25360));
    InMux I__3555 (
            .O(N__25408),
            .I(N__25360));
    InMux I__3554 (
            .O(N__25405),
            .I(N__25355));
    InMux I__3553 (
            .O(N__25402),
            .I(N__25355));
    InMux I__3552 (
            .O(N__25399),
            .I(N__25338));
    InMux I__3551 (
            .O(N__25396),
            .I(N__25338));
    InMux I__3550 (
            .O(N__25393),
            .I(N__25338));
    InMux I__3549 (
            .O(N__25390),
            .I(N__25338));
    InMux I__3548 (
            .O(N__25389),
            .I(N__25338));
    InMux I__3547 (
            .O(N__25388),
            .I(N__25338));
    InMux I__3546 (
            .O(N__25387),
            .I(N__25338));
    InMux I__3545 (
            .O(N__25386),
            .I(N__25338));
    InMux I__3544 (
            .O(N__25385),
            .I(N__25333));
    InMux I__3543 (
            .O(N__25382),
            .I(N__25333));
    LocalMux I__3542 (
            .O(N__25375),
            .I(N__25330));
    InMux I__3541 (
            .O(N__25374),
            .I(N__25325));
    InMux I__3540 (
            .O(N__25373),
            .I(N__25325));
    LocalMux I__3539 (
            .O(N__25360),
            .I(N__25321));
    LocalMux I__3538 (
            .O(N__25355),
            .I(N__25314));
    LocalMux I__3537 (
            .O(N__25338),
            .I(N__25314));
    LocalMux I__3536 (
            .O(N__25333),
            .I(N__25314));
    Span4Mux_v I__3535 (
            .O(N__25330),
            .I(N__25309));
    LocalMux I__3534 (
            .O(N__25325),
            .I(N__25309));
    InMux I__3533 (
            .O(N__25324),
            .I(N__25306));
    Span4Mux_v I__3532 (
            .O(N__25321),
            .I(N__25301));
    Span4Mux_v I__3531 (
            .O(N__25314),
            .I(N__25301));
    Span4Mux_h I__3530 (
            .O(N__25309),
            .I(N__25298));
    LocalMux I__3529 (
            .O(N__25306),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv4 I__3528 (
            .O(N__25301),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv4 I__3527 (
            .O(N__25298),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    InMux I__3526 (
            .O(N__25291),
            .I(N__25288));
    LocalMux I__3525 (
            .O(N__25288),
            .I(N__25285));
    Odrv4 I__3524 (
            .O(N__25285),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9 ));
    CascadeMux I__3523 (
            .O(N__25282),
            .I(N__25279));
    InMux I__3522 (
            .O(N__25279),
            .I(N__25276));
    LocalMux I__3521 (
            .O(N__25276),
            .I(N__25272));
    InMux I__3520 (
            .O(N__25275),
            .I(N__25269));
    Odrv4 I__3519 (
            .O(N__25272),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    LocalMux I__3518 (
            .O(N__25269),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    CascadeMux I__3517 (
            .O(N__25264),
            .I(N__25261));
    InMux I__3516 (
            .O(N__25261),
            .I(N__25258));
    LocalMux I__3515 (
            .O(N__25258),
            .I(N__25255));
    Span4Mux_h I__3514 (
            .O(N__25255),
            .I(N__25252));
    Odrv4 I__3513 (
            .O(N__25252),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ));
    CascadeMux I__3512 (
            .O(N__25249),
            .I(N__25246));
    InMux I__3511 (
            .O(N__25246),
            .I(N__25243));
    LocalMux I__3510 (
            .O(N__25243),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ));
    CascadeMux I__3509 (
            .O(N__25240),
            .I(N__25237));
    InMux I__3508 (
            .O(N__25237),
            .I(N__25234));
    LocalMux I__3507 (
            .O(N__25234),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ));
    CascadeMux I__3506 (
            .O(N__25231),
            .I(N__25228));
    InMux I__3505 (
            .O(N__25228),
            .I(N__25225));
    LocalMux I__3504 (
            .O(N__25225),
            .I(N__25222));
    Odrv12 I__3503 (
            .O(N__25222),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ));
    CascadeMux I__3502 (
            .O(N__25219),
            .I(N__25216));
    InMux I__3501 (
            .O(N__25216),
            .I(N__25213));
    LocalMux I__3500 (
            .O(N__25213),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ));
    CascadeMux I__3499 (
            .O(N__25210),
            .I(N__25207));
    InMux I__3498 (
            .O(N__25207),
            .I(N__25204));
    LocalMux I__3497 (
            .O(N__25204),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ));
    CascadeMux I__3496 (
            .O(N__25201),
            .I(N__25198));
    InMux I__3495 (
            .O(N__25198),
            .I(N__25195));
    LocalMux I__3494 (
            .O(N__25195),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ));
    CEMux I__3493 (
            .O(N__25192),
            .I(N__25186));
    CEMux I__3492 (
            .O(N__25191),
            .I(N__25183));
    CEMux I__3491 (
            .O(N__25190),
            .I(N__25180));
    CEMux I__3490 (
            .O(N__25189),
            .I(N__25177));
    LocalMux I__3489 (
            .O(N__25186),
            .I(N__25173));
    LocalMux I__3488 (
            .O(N__25183),
            .I(N__25170));
    LocalMux I__3487 (
            .O(N__25180),
            .I(N__25167));
    LocalMux I__3486 (
            .O(N__25177),
            .I(N__25164));
    CEMux I__3485 (
            .O(N__25176),
            .I(N__25161));
    Span4Mux_v I__3484 (
            .O(N__25173),
            .I(N__25158));
    Span4Mux_h I__3483 (
            .O(N__25170),
            .I(N__25155));
    Span4Mux_v I__3482 (
            .O(N__25167),
            .I(N__25152));
    Span4Mux_h I__3481 (
            .O(N__25164),
            .I(N__25147));
    LocalMux I__3480 (
            .O(N__25161),
            .I(N__25147));
    Odrv4 I__3479 (
            .O(N__25158),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv4 I__3478 (
            .O(N__25155),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv4 I__3477 (
            .O(N__25152),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv4 I__3476 (
            .O(N__25147),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ));
    CascadeMux I__3475 (
            .O(N__25138),
            .I(\phase_controller_inst2.start_timer_hc_0_sqmuxa_cascade_ ));
    InMux I__3474 (
            .O(N__25135),
            .I(N__25129));
    InMux I__3473 (
            .O(N__25134),
            .I(N__25126));
    InMux I__3472 (
            .O(N__25133),
            .I(N__25123));
    InMux I__3471 (
            .O(N__25132),
            .I(N__25120));
    LocalMux I__3470 (
            .O(N__25129),
            .I(N__25117));
    LocalMux I__3469 (
            .O(N__25126),
            .I(N__25114));
    LocalMux I__3468 (
            .O(N__25123),
            .I(N__25111));
    LocalMux I__3467 (
            .O(N__25120),
            .I(N__25104));
    Span4Mux_h I__3466 (
            .O(N__25117),
            .I(N__25104));
    Span4Mux_h I__3465 (
            .O(N__25114),
            .I(N__25099));
    Span4Mux_h I__3464 (
            .O(N__25111),
            .I(N__25099));
    InMux I__3463 (
            .O(N__25110),
            .I(N__25096));
    InMux I__3462 (
            .O(N__25109),
            .I(N__25093));
    Odrv4 I__3461 (
            .O(N__25104),
            .I(phase_controller_inst1_state_4));
    Odrv4 I__3460 (
            .O(N__25099),
            .I(phase_controller_inst1_state_4));
    LocalMux I__3459 (
            .O(N__25096),
            .I(phase_controller_inst1_state_4));
    LocalMux I__3458 (
            .O(N__25093),
            .I(phase_controller_inst1_state_4));
    CascadeMux I__3457 (
            .O(N__25084),
            .I(N__25081));
    InMux I__3456 (
            .O(N__25081),
            .I(N__25078));
    LocalMux I__3455 (
            .O(N__25078),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ));
    CascadeMux I__3454 (
            .O(N__25075),
            .I(N__25072));
    InMux I__3453 (
            .O(N__25072),
            .I(N__25069));
    LocalMux I__3452 (
            .O(N__25069),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ));
    CascadeMux I__3451 (
            .O(N__25066),
            .I(N__25063));
    InMux I__3450 (
            .O(N__25063),
            .I(N__25060));
    LocalMux I__3449 (
            .O(N__25060),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ));
    CascadeMux I__3448 (
            .O(N__25057),
            .I(N__25054));
    InMux I__3447 (
            .O(N__25054),
            .I(N__25051));
    LocalMux I__3446 (
            .O(N__25051),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ));
    CascadeMux I__3445 (
            .O(N__25048),
            .I(N__25045));
    InMux I__3444 (
            .O(N__25045),
            .I(N__25042));
    LocalMux I__3443 (
            .O(N__25042),
            .I(N__25039));
    Span4Mux_v I__3442 (
            .O(N__25039),
            .I(N__25036));
    Odrv4 I__3441 (
            .O(N__25036),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ));
    InMux I__3440 (
            .O(N__25033),
            .I(N__25030));
    LocalMux I__3439 (
            .O(N__25030),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ));
    CascadeMux I__3438 (
            .O(N__25027),
            .I(N__25024));
    InMux I__3437 (
            .O(N__25024),
            .I(N__25021));
    LocalMux I__3436 (
            .O(N__25021),
            .I(N__25018));
    Odrv4 I__3435 (
            .O(N__25018),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ));
    CascadeMux I__3434 (
            .O(N__25015),
            .I(N__25012));
    InMux I__3433 (
            .O(N__25012),
            .I(N__25009));
    LocalMux I__3432 (
            .O(N__25009),
            .I(N__25006));
    Span4Mux_v I__3431 (
            .O(N__25006),
            .I(N__25003));
    Odrv4 I__3430 (
            .O(N__25003),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ));
    CascadeMux I__3429 (
            .O(N__25000),
            .I(N__24997));
    InMux I__3428 (
            .O(N__24997),
            .I(N__24994));
    LocalMux I__3427 (
            .O(N__24994),
            .I(N__24991));
    Span4Mux_h I__3426 (
            .O(N__24991),
            .I(N__24988));
    Odrv4 I__3425 (
            .O(N__24988),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ));
    InMux I__3424 (
            .O(N__24985),
            .I(N__24981));
    InMux I__3423 (
            .O(N__24984),
            .I(N__24978));
    LocalMux I__3422 (
            .O(N__24981),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    LocalMux I__3421 (
            .O(N__24978),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__3420 (
            .O(N__24973),
            .I(N__24970));
    LocalMux I__3419 (
            .O(N__24970),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ));
    InMux I__3418 (
            .O(N__24967),
            .I(N__24963));
    InMux I__3417 (
            .O(N__24966),
            .I(N__24960));
    LocalMux I__3416 (
            .O(N__24963),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    LocalMux I__3415 (
            .O(N__24960),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__3414 (
            .O(N__24955),
            .I(N__24952));
    LocalMux I__3413 (
            .O(N__24952),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ));
    InMux I__3412 (
            .O(N__24949),
            .I(N__24945));
    InMux I__3411 (
            .O(N__24948),
            .I(N__24942));
    LocalMux I__3410 (
            .O(N__24945),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    LocalMux I__3409 (
            .O(N__24942),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__3408 (
            .O(N__24937),
            .I(N__24934));
    LocalMux I__3407 (
            .O(N__24934),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ));
    InMux I__3406 (
            .O(N__24931),
            .I(N__24928));
    LocalMux I__3405 (
            .O(N__24928),
            .I(N__24924));
    InMux I__3404 (
            .O(N__24927),
            .I(N__24921));
    Span4Mux_h I__3403 (
            .O(N__24924),
            .I(N__24918));
    LocalMux I__3402 (
            .O(N__24921),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv4 I__3401 (
            .O(N__24918),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    InMux I__3400 (
            .O(N__24913),
            .I(N__24910));
    LocalMux I__3399 (
            .O(N__24910),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_16 ));
    InMux I__3398 (
            .O(N__24907),
            .I(N__24903));
    InMux I__3397 (
            .O(N__24906),
            .I(N__24900));
    LocalMux I__3396 (
            .O(N__24903),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    LocalMux I__3395 (
            .O(N__24900),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__3394 (
            .O(N__24895),
            .I(N__24892));
    LocalMux I__3393 (
            .O(N__24892),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_17 ));
    InMux I__3392 (
            .O(N__24889),
            .I(N__24885));
    InMux I__3391 (
            .O(N__24888),
            .I(N__24882));
    LocalMux I__3390 (
            .O(N__24885),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    LocalMux I__3389 (
            .O(N__24882),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__3388 (
            .O(N__24877),
            .I(N__24874));
    LocalMux I__3387 (
            .O(N__24874),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_18 ));
    InMux I__3386 (
            .O(N__24871),
            .I(N__24867));
    InMux I__3385 (
            .O(N__24870),
            .I(N__24864));
    LocalMux I__3384 (
            .O(N__24867),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    LocalMux I__3383 (
            .O(N__24864),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__3382 (
            .O(N__24859),
            .I(N__24856));
    LocalMux I__3381 (
            .O(N__24856),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_19 ));
    InMux I__3380 (
            .O(N__24853),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ));
    InMux I__3379 (
            .O(N__24850),
            .I(N__24847));
    LocalMux I__3378 (
            .O(N__24847),
            .I(N__24843));
    InMux I__3377 (
            .O(N__24846),
            .I(N__24840));
    Odrv4 I__3376 (
            .O(N__24843),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    LocalMux I__3375 (
            .O(N__24840),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__3374 (
            .O(N__24835),
            .I(N__24832));
    LocalMux I__3373 (
            .O(N__24832),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ));
    CascadeMux I__3372 (
            .O(N__24829),
            .I(N__24826));
    InMux I__3371 (
            .O(N__24826),
            .I(N__24823));
    LocalMux I__3370 (
            .O(N__24823),
            .I(N__24820));
    Odrv4 I__3369 (
            .O(N__24820),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ));
    CascadeMux I__3368 (
            .O(N__24817),
            .I(N__24814));
    InMux I__3367 (
            .O(N__24814),
            .I(N__24811));
    LocalMux I__3366 (
            .O(N__24811),
            .I(N__24807));
    InMux I__3365 (
            .O(N__24810),
            .I(N__24804));
    Odrv4 I__3364 (
            .O(N__24807),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    LocalMux I__3363 (
            .O(N__24804),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__3362 (
            .O(N__24799),
            .I(N__24796));
    LocalMux I__3361 (
            .O(N__24796),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ));
    CascadeMux I__3360 (
            .O(N__24793),
            .I(N__24790));
    InMux I__3359 (
            .O(N__24790),
            .I(N__24787));
    LocalMux I__3358 (
            .O(N__24787),
            .I(N__24783));
    InMux I__3357 (
            .O(N__24786),
            .I(N__24780));
    Odrv4 I__3356 (
            .O(N__24783),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    LocalMux I__3355 (
            .O(N__24780),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__3354 (
            .O(N__24775),
            .I(N__24772));
    LocalMux I__3353 (
            .O(N__24772),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ));
    CascadeMux I__3352 (
            .O(N__24769),
            .I(N__24766));
    InMux I__3351 (
            .O(N__24766),
            .I(N__24763));
    LocalMux I__3350 (
            .O(N__24763),
            .I(N__24759));
    InMux I__3349 (
            .O(N__24762),
            .I(N__24756));
    Odrv4 I__3348 (
            .O(N__24759),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    LocalMux I__3347 (
            .O(N__24756),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__3346 (
            .O(N__24751),
            .I(N__24748));
    LocalMux I__3345 (
            .O(N__24748),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ));
    InMux I__3344 (
            .O(N__24745),
            .I(N__24741));
    InMux I__3343 (
            .O(N__24744),
            .I(N__24738));
    LocalMux I__3342 (
            .O(N__24741),
            .I(N__24735));
    LocalMux I__3341 (
            .O(N__24738),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    Odrv4 I__3340 (
            .O(N__24735),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__3339 (
            .O(N__24730),
            .I(N__24727));
    LocalMux I__3338 (
            .O(N__24727),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ));
    InMux I__3337 (
            .O(N__24724),
            .I(N__24720));
    InMux I__3336 (
            .O(N__24723),
            .I(N__24717));
    LocalMux I__3335 (
            .O(N__24720),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    LocalMux I__3334 (
            .O(N__24717),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__3333 (
            .O(N__24712),
            .I(N__24709));
    LocalMux I__3332 (
            .O(N__24709),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ));
    InMux I__3331 (
            .O(N__24706),
            .I(N__24702));
    InMux I__3330 (
            .O(N__24705),
            .I(N__24699));
    LocalMux I__3329 (
            .O(N__24702),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    LocalMux I__3328 (
            .O(N__24699),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__3327 (
            .O(N__24694),
            .I(N__24691));
    LocalMux I__3326 (
            .O(N__24691),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ));
    InMux I__3325 (
            .O(N__24688),
            .I(N__24684));
    InMux I__3324 (
            .O(N__24687),
            .I(N__24681));
    LocalMux I__3323 (
            .O(N__24684),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    LocalMux I__3322 (
            .O(N__24681),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__3321 (
            .O(N__24676),
            .I(N__24673));
    LocalMux I__3320 (
            .O(N__24673),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ));
    InMux I__3319 (
            .O(N__24670),
            .I(N__24666));
    InMux I__3318 (
            .O(N__24669),
            .I(N__24663));
    LocalMux I__3317 (
            .O(N__24666),
            .I(N__24658));
    LocalMux I__3316 (
            .O(N__24663),
            .I(N__24658));
    Span4Mux_v I__3315 (
            .O(N__24658),
            .I(N__24655));
    Odrv4 I__3314 (
            .O(N__24655),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    InMux I__3313 (
            .O(N__24652),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ));
    InMux I__3312 (
            .O(N__24649),
            .I(N__24646));
    LocalMux I__3311 (
            .O(N__24646),
            .I(N__24642));
    InMux I__3310 (
            .O(N__24645),
            .I(N__24639));
    Span4Mux_v I__3309 (
            .O(N__24642),
            .I(N__24634));
    LocalMux I__3308 (
            .O(N__24639),
            .I(N__24634));
    Odrv4 I__3307 (
            .O(N__24634),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    InMux I__3306 (
            .O(N__24631),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ));
    InMux I__3305 (
            .O(N__24628),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ));
    CascadeMux I__3304 (
            .O(N__24625),
            .I(N__24621));
    CascadeMux I__3303 (
            .O(N__24624),
            .I(N__24618));
    InMux I__3302 (
            .O(N__24621),
            .I(N__24609));
    InMux I__3301 (
            .O(N__24618),
            .I(N__24609));
    CascadeMux I__3300 (
            .O(N__24617),
            .I(N__24605));
    CascadeMux I__3299 (
            .O(N__24616),
            .I(N__24602));
    CascadeMux I__3298 (
            .O(N__24615),
            .I(N__24597));
    CascadeMux I__3297 (
            .O(N__24614),
            .I(N__24594));
    LocalMux I__3296 (
            .O(N__24609),
            .I(N__24590));
    InMux I__3295 (
            .O(N__24608),
            .I(N__24581));
    InMux I__3294 (
            .O(N__24605),
            .I(N__24581));
    InMux I__3293 (
            .O(N__24602),
            .I(N__24581));
    InMux I__3292 (
            .O(N__24601),
            .I(N__24581));
    InMux I__3291 (
            .O(N__24600),
            .I(N__24578));
    InMux I__3290 (
            .O(N__24597),
            .I(N__24575));
    InMux I__3289 (
            .O(N__24594),
            .I(N__24570));
    InMux I__3288 (
            .O(N__24593),
            .I(N__24570));
    Span4Mux_v I__3287 (
            .O(N__24590),
            .I(N__24563));
    LocalMux I__3286 (
            .O(N__24581),
            .I(N__24563));
    LocalMux I__3285 (
            .O(N__24578),
            .I(N__24563));
    LocalMux I__3284 (
            .O(N__24575),
            .I(N__24558));
    LocalMux I__3283 (
            .O(N__24570),
            .I(N__24558));
    Span4Mux_h I__3282 (
            .O(N__24563),
            .I(N__24555));
    Span4Mux_h I__3281 (
            .O(N__24558),
            .I(N__24552));
    Span4Mux_v I__3280 (
            .O(N__24555),
            .I(N__24549));
    Span4Mux_v I__3279 (
            .O(N__24552),
            .I(N__24546));
    Span4Mux_h I__3278 (
            .O(N__24549),
            .I(N__24543));
    Span4Mux_h I__3277 (
            .O(N__24546),
            .I(N__24540));
    Odrv4 I__3276 (
            .O(N__24543),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    Odrv4 I__3275 (
            .O(N__24540),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    CascadeMux I__3274 (
            .O(N__24535),
            .I(N__24531));
    InMux I__3273 (
            .O(N__24534),
            .I(N__24528));
    InMux I__3272 (
            .O(N__24531),
            .I(N__24525));
    LocalMux I__3271 (
            .O(N__24528),
            .I(N__24519));
    LocalMux I__3270 (
            .O(N__24525),
            .I(N__24519));
    InMux I__3269 (
            .O(N__24524),
            .I(N__24516));
    Odrv4 I__3268 (
            .O(N__24519),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__3267 (
            .O(N__24516),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    InMux I__3266 (
            .O(N__24511),
            .I(N__24508));
    LocalMux I__3265 (
            .O(N__24508),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ));
    InMux I__3264 (
            .O(N__24505),
            .I(N__24502));
    LocalMux I__3263 (
            .O(N__24502),
            .I(N__24498));
    InMux I__3262 (
            .O(N__24501),
            .I(N__24495));
    Odrv4 I__3261 (
            .O(N__24498),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    LocalMux I__3260 (
            .O(N__24495),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__3259 (
            .O(N__24490),
            .I(N__24487));
    LocalMux I__3258 (
            .O(N__24487),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ));
    CascadeMux I__3257 (
            .O(N__24484),
            .I(N__24481));
    InMux I__3256 (
            .O(N__24481),
            .I(N__24478));
    LocalMux I__3255 (
            .O(N__24478),
            .I(N__24474));
    InMux I__3254 (
            .O(N__24477),
            .I(N__24471));
    Odrv4 I__3253 (
            .O(N__24474),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    LocalMux I__3252 (
            .O(N__24471),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__3251 (
            .O(N__24466),
            .I(N__24463));
    LocalMux I__3250 (
            .O(N__24463),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ));
    InMux I__3249 (
            .O(N__24460),
            .I(N__24456));
    InMux I__3248 (
            .O(N__24459),
            .I(N__24453));
    LocalMux I__3247 (
            .O(N__24456),
            .I(N__24450));
    LocalMux I__3246 (
            .O(N__24453),
            .I(N__24447));
    Odrv4 I__3245 (
            .O(N__24450),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    Odrv4 I__3244 (
            .O(N__24447),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__3243 (
            .O(N__24442),
            .I(N__24439));
    LocalMux I__3242 (
            .O(N__24439),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ));
    InMux I__3241 (
            .O(N__24436),
            .I(N__24430));
    InMux I__3240 (
            .O(N__24435),
            .I(N__24430));
    LocalMux I__3239 (
            .O(N__24430),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    InMux I__3238 (
            .O(N__24427),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ));
    InMux I__3237 (
            .O(N__24424),
            .I(N__24420));
    InMux I__3236 (
            .O(N__24423),
            .I(N__24417));
    LocalMux I__3235 (
            .O(N__24420),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    LocalMux I__3234 (
            .O(N__24417),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    InMux I__3233 (
            .O(N__24412),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ));
    CascadeMux I__3232 (
            .O(N__24409),
            .I(N__24405));
    CascadeMux I__3231 (
            .O(N__24408),
            .I(N__24402));
    InMux I__3230 (
            .O(N__24405),
            .I(N__24397));
    InMux I__3229 (
            .O(N__24402),
            .I(N__24397));
    LocalMux I__3228 (
            .O(N__24397),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    InMux I__3227 (
            .O(N__24394),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ));
    InMux I__3226 (
            .O(N__24391),
            .I(N__24385));
    InMux I__3225 (
            .O(N__24390),
            .I(N__24385));
    LocalMux I__3224 (
            .O(N__24385),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ));
    InMux I__3223 (
            .O(N__24382),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ));
    InMux I__3222 (
            .O(N__24379),
            .I(N__24376));
    LocalMux I__3221 (
            .O(N__24376),
            .I(N__24372));
    InMux I__3220 (
            .O(N__24375),
            .I(N__24369));
    Odrv4 I__3219 (
            .O(N__24372),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ));
    LocalMux I__3218 (
            .O(N__24369),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ));
    InMux I__3217 (
            .O(N__24364),
            .I(bfn_9_11_0_));
    InMux I__3216 (
            .O(N__24361),
            .I(N__24357));
    InMux I__3215 (
            .O(N__24360),
            .I(N__24354));
    LocalMux I__3214 (
            .O(N__24357),
            .I(N__24351));
    LocalMux I__3213 (
            .O(N__24354),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ));
    Odrv4 I__3212 (
            .O(N__24351),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ));
    InMux I__3211 (
            .O(N__24346),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ));
    InMux I__3210 (
            .O(N__24343),
            .I(N__24339));
    InMux I__3209 (
            .O(N__24342),
            .I(N__24336));
    LocalMux I__3208 (
            .O(N__24339),
            .I(N__24333));
    LocalMux I__3207 (
            .O(N__24336),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ));
    Odrv4 I__3206 (
            .O(N__24333),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ));
    InMux I__3205 (
            .O(N__24328),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ));
    CascadeMux I__3204 (
            .O(N__24325),
            .I(N__24321));
    InMux I__3203 (
            .O(N__24324),
            .I(N__24318));
    InMux I__3202 (
            .O(N__24321),
            .I(N__24315));
    LocalMux I__3201 (
            .O(N__24318),
            .I(N__24312));
    LocalMux I__3200 (
            .O(N__24315),
            .I(N__24309));
    Odrv4 I__3199 (
            .O(N__24312),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    Odrv4 I__3198 (
            .O(N__24309),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    InMux I__3197 (
            .O(N__24304),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ));
    InMux I__3196 (
            .O(N__24301),
            .I(N__24298));
    LocalMux I__3195 (
            .O(N__24298),
            .I(N__24294));
    InMux I__3194 (
            .O(N__24297),
            .I(N__24291));
    Span4Mux_v I__3193 (
            .O(N__24294),
            .I(N__24288));
    LocalMux I__3192 (
            .O(N__24291),
            .I(N__24285));
    Odrv4 I__3191 (
            .O(N__24288),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    Odrv4 I__3190 (
            .O(N__24285),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    InMux I__3189 (
            .O(N__24280),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ));
    InMux I__3188 (
            .O(N__24277),
            .I(N__24271));
    InMux I__3187 (
            .O(N__24276),
            .I(N__24271));
    LocalMux I__3186 (
            .O(N__24271),
            .I(N__24268));
    Odrv4 I__3185 (
            .O(N__24268),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    InMux I__3184 (
            .O(N__24265),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ));
    InMux I__3183 (
            .O(N__24262),
            .I(N__24256));
    InMux I__3182 (
            .O(N__24261),
            .I(N__24256));
    LocalMux I__3181 (
            .O(N__24256),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    InMux I__3180 (
            .O(N__24253),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ));
    CascadeMux I__3179 (
            .O(N__24250),
            .I(N__24247));
    InMux I__3178 (
            .O(N__24247),
            .I(N__24244));
    LocalMux I__3177 (
            .O(N__24244),
            .I(N__24241));
    Odrv4 I__3176 (
            .O(N__24241),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ));
    CascadeMux I__3175 (
            .O(N__24238),
            .I(N__24235));
    InMux I__3174 (
            .O(N__24235),
            .I(N__24229));
    InMux I__3173 (
            .O(N__24234),
            .I(N__24229));
    LocalMux I__3172 (
            .O(N__24229),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    InMux I__3171 (
            .O(N__24226),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ));
    InMux I__3170 (
            .O(N__24223),
            .I(N__24219));
    InMux I__3169 (
            .O(N__24222),
            .I(N__24216));
    LocalMux I__3168 (
            .O(N__24219),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    LocalMux I__3167 (
            .O(N__24216),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    InMux I__3166 (
            .O(N__24211),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ));
    InMux I__3165 (
            .O(N__24208),
            .I(N__24204));
    CascadeMux I__3164 (
            .O(N__24207),
            .I(N__24201));
    LocalMux I__3163 (
            .O(N__24204),
            .I(N__24198));
    InMux I__3162 (
            .O(N__24201),
            .I(N__24195));
    Odrv4 I__3161 (
            .O(N__24198),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    LocalMux I__3160 (
            .O(N__24195),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    InMux I__3159 (
            .O(N__24190),
            .I(bfn_9_10_0_));
    InMux I__3158 (
            .O(N__24187),
            .I(N__24183));
    InMux I__3157 (
            .O(N__24186),
            .I(N__24180));
    LocalMux I__3156 (
            .O(N__24183),
            .I(N__24177));
    LocalMux I__3155 (
            .O(N__24180),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    Odrv4 I__3154 (
            .O(N__24177),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    InMux I__3153 (
            .O(N__24172),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ));
    CascadeMux I__3152 (
            .O(N__24169),
            .I(N__24166));
    InMux I__3151 (
            .O(N__24166),
            .I(N__24162));
    InMux I__3150 (
            .O(N__24165),
            .I(N__24159));
    LocalMux I__3149 (
            .O(N__24162),
            .I(N__24156));
    LocalMux I__3148 (
            .O(N__24159),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    Odrv4 I__3147 (
            .O(N__24156),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    InMux I__3146 (
            .O(N__24151),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ));
    InMux I__3145 (
            .O(N__24148),
            .I(N__24142));
    InMux I__3144 (
            .O(N__24147),
            .I(N__24142));
    LocalMux I__3143 (
            .O(N__24142),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    InMux I__3142 (
            .O(N__24139),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ));
    InMux I__3141 (
            .O(N__24136),
            .I(N__24132));
    InMux I__3140 (
            .O(N__24135),
            .I(N__24127));
    LocalMux I__3139 (
            .O(N__24132),
            .I(N__24124));
    InMux I__3138 (
            .O(N__24131),
            .I(N__24121));
    InMux I__3137 (
            .O(N__24130),
            .I(N__24118));
    LocalMux I__3136 (
            .O(N__24127),
            .I(N__24115));
    Span4Mux_v I__3135 (
            .O(N__24124),
            .I(N__24110));
    LocalMux I__3134 (
            .O(N__24121),
            .I(N__24110));
    LocalMux I__3133 (
            .O(N__24118),
            .I(N__24107));
    Span4Mux_v I__3132 (
            .O(N__24115),
            .I(N__24104));
    Span4Mux_h I__3131 (
            .O(N__24110),
            .I(N__24101));
    Span12Mux_s7_v I__3130 (
            .O(N__24107),
            .I(N__24098));
    Span4Mux_h I__3129 (
            .O(N__24104),
            .I(N__24095));
    Span4Mux_h I__3128 (
            .O(N__24101),
            .I(N__24092));
    Odrv12 I__3127 (
            .O(N__24098),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    Odrv4 I__3126 (
            .O(N__24095),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    Odrv4 I__3125 (
            .O(N__24092),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    InMux I__3124 (
            .O(N__24085),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ));
    InMux I__3123 (
            .O(N__24082),
            .I(N__24079));
    LocalMux I__3122 (
            .O(N__24079),
            .I(N__24074));
    InMux I__3121 (
            .O(N__24078),
            .I(N__24071));
    InMux I__3120 (
            .O(N__24077),
            .I(N__24068));
    Span4Mux_v I__3119 (
            .O(N__24074),
            .I(N__24061));
    LocalMux I__3118 (
            .O(N__24071),
            .I(N__24061));
    LocalMux I__3117 (
            .O(N__24068),
            .I(N__24061));
    Span4Mux_h I__3116 (
            .O(N__24061),
            .I(N__24058));
    Span4Mux_h I__3115 (
            .O(N__24058),
            .I(N__24055));
    Odrv4 I__3114 (
            .O(N__24055),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    InMux I__3113 (
            .O(N__24052),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ));
    InMux I__3112 (
            .O(N__24049),
            .I(N__24044));
    InMux I__3111 (
            .O(N__24048),
            .I(N__24041));
    InMux I__3110 (
            .O(N__24047),
            .I(N__24038));
    LocalMux I__3109 (
            .O(N__24044),
            .I(N__24031));
    LocalMux I__3108 (
            .O(N__24041),
            .I(N__24031));
    LocalMux I__3107 (
            .O(N__24038),
            .I(N__24031));
    Span4Mux_h I__3106 (
            .O(N__24031),
            .I(N__24028));
    Span4Mux_h I__3105 (
            .O(N__24028),
            .I(N__24025));
    Odrv4 I__3104 (
            .O(N__24025),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    InMux I__3103 (
            .O(N__24022),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ));
    InMux I__3102 (
            .O(N__24019),
            .I(N__24014));
    InMux I__3101 (
            .O(N__24018),
            .I(N__24011));
    InMux I__3100 (
            .O(N__24017),
            .I(N__24008));
    LocalMux I__3099 (
            .O(N__24014),
            .I(N__24001));
    LocalMux I__3098 (
            .O(N__24011),
            .I(N__24001));
    LocalMux I__3097 (
            .O(N__24008),
            .I(N__24001));
    Span4Mux_h I__3096 (
            .O(N__24001),
            .I(N__23998));
    Span4Mux_h I__3095 (
            .O(N__23998),
            .I(N__23995));
    Odrv4 I__3094 (
            .O(N__23995),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    InMux I__3093 (
            .O(N__23992),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ));
    InMux I__3092 (
            .O(N__23989),
            .I(N__23986));
    LocalMux I__3091 (
            .O(N__23986),
            .I(N__23981));
    InMux I__3090 (
            .O(N__23985),
            .I(N__23978));
    InMux I__3089 (
            .O(N__23984),
            .I(N__23975));
    Span4Mux_v I__3088 (
            .O(N__23981),
            .I(N__23968));
    LocalMux I__3087 (
            .O(N__23978),
            .I(N__23968));
    LocalMux I__3086 (
            .O(N__23975),
            .I(N__23968));
    Span4Mux_h I__3085 (
            .O(N__23968),
            .I(N__23965));
    Span4Mux_h I__3084 (
            .O(N__23965),
            .I(N__23962));
    Odrv4 I__3083 (
            .O(N__23962),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    InMux I__3082 (
            .O(N__23959),
            .I(bfn_9_9_0_));
    InMux I__3081 (
            .O(N__23956),
            .I(N__23952));
    InMux I__3080 (
            .O(N__23955),
            .I(N__23949));
    LocalMux I__3079 (
            .O(N__23952),
            .I(N__23943));
    LocalMux I__3078 (
            .O(N__23949),
            .I(N__23943));
    InMux I__3077 (
            .O(N__23948),
            .I(N__23940));
    Sp12to4 I__3076 (
            .O(N__23943),
            .I(N__23935));
    LocalMux I__3075 (
            .O(N__23940),
            .I(N__23935));
    Span12Mux_s9_h I__3074 (
            .O(N__23935),
            .I(N__23932));
    Odrv12 I__3073 (
            .O(N__23932),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    InMux I__3072 (
            .O(N__23929),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ));
    CascadeMux I__3071 (
            .O(N__23926),
            .I(N__23923));
    InMux I__3070 (
            .O(N__23923),
            .I(N__23920));
    LocalMux I__3069 (
            .O(N__23920),
            .I(N__23916));
    InMux I__3068 (
            .O(N__23919),
            .I(N__23913));
    Odrv4 I__3067 (
            .O(N__23916),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ));
    LocalMux I__3066 (
            .O(N__23913),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ));
    InMux I__3065 (
            .O(N__23908),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ));
    InMux I__3064 (
            .O(N__23905),
            .I(N__23899));
    InMux I__3063 (
            .O(N__23904),
            .I(N__23899));
    LocalMux I__3062 (
            .O(N__23899),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ));
    InMux I__3061 (
            .O(N__23896),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ));
    CascadeMux I__3060 (
            .O(N__23893),
            .I(N__23890));
    InMux I__3059 (
            .O(N__23890),
            .I(N__23887));
    LocalMux I__3058 (
            .O(N__23887),
            .I(\phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa ));
    InMux I__3057 (
            .O(N__23884),
            .I(N__23881));
    LocalMux I__3056 (
            .O(N__23881),
            .I(N__23877));
    InMux I__3055 (
            .O(N__23880),
            .I(N__23874));
    Span4Mux_v I__3054 (
            .O(N__23877),
            .I(N__23868));
    LocalMux I__3053 (
            .O(N__23874),
            .I(N__23868));
    InMux I__3052 (
            .O(N__23873),
            .I(N__23865));
    Span4Mux_h I__3051 (
            .O(N__23868),
            .I(N__23859));
    LocalMux I__3050 (
            .O(N__23865),
            .I(N__23859));
    InMux I__3049 (
            .O(N__23864),
            .I(N__23856));
    Sp12to4 I__3048 (
            .O(N__23859),
            .I(N__23853));
    LocalMux I__3047 (
            .O(N__23856),
            .I(\phase_controller_inst1.hc_time_passed ));
    Odrv12 I__3046 (
            .O(N__23853),
            .I(\phase_controller_inst1.hc_time_passed ));
    InMux I__3045 (
            .O(N__23848),
            .I(N__23845));
    LocalMux I__3044 (
            .O(N__23845),
            .I(N__23842));
    Glb2LocalMux I__3043 (
            .O(N__23842),
            .I(N__23839));
    GlobalMux I__3042 (
            .O(N__23839),
            .I(clk_12mhz));
    IoInMux I__3041 (
            .O(N__23836),
            .I(N__23833));
    LocalMux I__3040 (
            .O(N__23833),
            .I(N__23830));
    Span4Mux_s0_v I__3039 (
            .O(N__23830),
            .I(N__23827));
    Odrv4 I__3038 (
            .O(N__23827),
            .I(GB_BUFFER_clk_12mhz_THRU_CO));
    InMux I__3037 (
            .O(N__23824),
            .I(N__23821));
    LocalMux I__3036 (
            .O(N__23821),
            .I(N__23818));
    Odrv12 I__3035 (
            .O(N__23818),
            .I(il_min_comp1_c));
    InMux I__3034 (
            .O(N__23815),
            .I(N__23812));
    LocalMux I__3033 (
            .O(N__23812),
            .I(N__23809));
    Span4Mux_h I__3032 (
            .O(N__23809),
            .I(N__23806));
    Odrv4 I__3031 (
            .O(N__23806),
            .I(il_min_comp1_D1));
    InMux I__3030 (
            .O(N__23803),
            .I(N__23800));
    LocalMux I__3029 (
            .O(N__23800),
            .I(N__23797));
    Span4Mux_h I__3028 (
            .O(N__23797),
            .I(N__23794));
    Span4Mux_h I__3027 (
            .O(N__23794),
            .I(N__23791));
    Odrv4 I__3026 (
            .O(N__23791),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ));
    InMux I__3025 (
            .O(N__23788),
            .I(N__23785));
    LocalMux I__3024 (
            .O(N__23785),
            .I(N__23782));
    Span12Mux_s9_h I__3023 (
            .O(N__23782),
            .I(N__23779));
    Odrv12 I__3022 (
            .O(N__23779),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ));
    InMux I__3021 (
            .O(N__23776),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ));
    InMux I__3020 (
            .O(N__23773),
            .I(N__23770));
    LocalMux I__3019 (
            .O(N__23770),
            .I(N__23767));
    Span4Mux_h I__3018 (
            .O(N__23767),
            .I(N__23764));
    Span4Mux_h I__3017 (
            .O(N__23764),
            .I(N__23761));
    Odrv4 I__3016 (
            .O(N__23761),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ));
    InMux I__3015 (
            .O(N__23758),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ));
    InMux I__3014 (
            .O(N__23755),
            .I(N__23752));
    LocalMux I__3013 (
            .O(N__23752),
            .I(N__23748));
    InMux I__3012 (
            .O(N__23751),
            .I(N__23745));
    Span4Mux_s2_h I__3011 (
            .O(N__23748),
            .I(N__23739));
    LocalMux I__3010 (
            .O(N__23745),
            .I(N__23739));
    InMux I__3009 (
            .O(N__23744),
            .I(N__23736));
    Sp12to4 I__3008 (
            .O(N__23739),
            .I(N__23731));
    LocalMux I__3007 (
            .O(N__23736),
            .I(N__23731));
    Span12Mux_s7_v I__3006 (
            .O(N__23731),
            .I(N__23728));
    Odrv12 I__3005 (
            .O(N__23728),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    InMux I__3004 (
            .O(N__23725),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ));
    InMux I__3003 (
            .O(N__23722),
            .I(N__23718));
    InMux I__3002 (
            .O(N__23721),
            .I(N__23715));
    LocalMux I__3001 (
            .O(N__23718),
            .I(N__23712));
    LocalMux I__3000 (
            .O(N__23715),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    Odrv4 I__2999 (
            .O(N__23712),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__2998 (
            .O(N__23707),
            .I(N__23704));
    LocalMux I__2997 (
            .O(N__23704),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14 ));
    InMux I__2996 (
            .O(N__23701),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ));
    InMux I__2995 (
            .O(N__23698),
            .I(N__23694));
    InMux I__2994 (
            .O(N__23697),
            .I(N__23691));
    LocalMux I__2993 (
            .O(N__23694),
            .I(N__23688));
    LocalMux I__2992 (
            .O(N__23691),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    Odrv4 I__2991 (
            .O(N__23688),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    CascadeMux I__2990 (
            .O(N__23683),
            .I(N__23680));
    InMux I__2989 (
            .O(N__23680),
            .I(N__23677));
    LocalMux I__2988 (
            .O(N__23677),
            .I(N__23674));
    Odrv4 I__2987 (
            .O(N__23674),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15 ));
    InMux I__2986 (
            .O(N__23671),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ));
    InMux I__2985 (
            .O(N__23668),
            .I(N__23665));
    LocalMux I__2984 (
            .O(N__23665),
            .I(N__23661));
    InMux I__2983 (
            .O(N__23664),
            .I(N__23658));
    Odrv4 I__2982 (
            .O(N__23661),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    LocalMux I__2981 (
            .O(N__23658),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    CascadeMux I__2980 (
            .O(N__23653),
            .I(N__23650));
    InMux I__2979 (
            .O(N__23650),
            .I(N__23647));
    LocalMux I__2978 (
            .O(N__23647),
            .I(N__23644));
    Span4Mux_h I__2977 (
            .O(N__23644),
            .I(N__23641));
    Odrv4 I__2976 (
            .O(N__23641),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16 ));
    InMux I__2975 (
            .O(N__23638),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ));
    InMux I__2974 (
            .O(N__23635),
            .I(N__23631));
    InMux I__2973 (
            .O(N__23634),
            .I(N__23628));
    LocalMux I__2972 (
            .O(N__23631),
            .I(N__23625));
    LocalMux I__2971 (
            .O(N__23628),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    Odrv4 I__2970 (
            .O(N__23625),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__2969 (
            .O(N__23620),
            .I(N__23617));
    LocalMux I__2968 (
            .O(N__23617),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17 ));
    InMux I__2967 (
            .O(N__23614),
            .I(bfn_8_22_0_));
    InMux I__2966 (
            .O(N__23611),
            .I(N__23607));
    InMux I__2965 (
            .O(N__23610),
            .I(N__23604));
    LocalMux I__2964 (
            .O(N__23607),
            .I(N__23601));
    LocalMux I__2963 (
            .O(N__23604),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    Odrv4 I__2962 (
            .O(N__23601),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__2961 (
            .O(N__23596),
            .I(N__23593));
    LocalMux I__2960 (
            .O(N__23593),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18 ));
    InMux I__2959 (
            .O(N__23590),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ));
    InMux I__2958 (
            .O(N__23587),
            .I(N__23583));
    InMux I__2957 (
            .O(N__23586),
            .I(N__23580));
    LocalMux I__2956 (
            .O(N__23583),
            .I(N__23577));
    LocalMux I__2955 (
            .O(N__23580),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    Odrv4 I__2954 (
            .O(N__23577),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__2953 (
            .O(N__23572),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17 ));
    InMux I__2952 (
            .O(N__23569),
            .I(N__23566));
    LocalMux I__2951 (
            .O(N__23566),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19 ));
    InMux I__2950 (
            .O(N__23563),
            .I(N__23560));
    LocalMux I__2949 (
            .O(N__23560),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5 ));
    InMux I__2948 (
            .O(N__23557),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ));
    InMux I__2947 (
            .O(N__23554),
            .I(N__23550));
    InMux I__2946 (
            .O(N__23553),
            .I(N__23547));
    LocalMux I__2945 (
            .O(N__23550),
            .I(N__23542));
    LocalMux I__2944 (
            .O(N__23547),
            .I(N__23542));
    Span4Mux_v I__2943 (
            .O(N__23542),
            .I(N__23539));
    Odrv4 I__2942 (
            .O(N__23539),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__2941 (
            .O(N__23536),
            .I(N__23533));
    LocalMux I__2940 (
            .O(N__23533),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6 ));
    InMux I__2939 (
            .O(N__23530),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ));
    InMux I__2938 (
            .O(N__23527),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ));
    InMux I__2937 (
            .O(N__23524),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ));
    InMux I__2936 (
            .O(N__23521),
            .I(bfn_8_21_0_));
    InMux I__2935 (
            .O(N__23518),
            .I(N__23514));
    InMux I__2934 (
            .O(N__23517),
            .I(N__23511));
    LocalMux I__2933 (
            .O(N__23514),
            .I(N__23508));
    LocalMux I__2932 (
            .O(N__23511),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    Odrv4 I__2931 (
            .O(N__23508),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__2930 (
            .O(N__23503),
            .I(N__23500));
    LocalMux I__2929 (
            .O(N__23500),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10 ));
    InMux I__2928 (
            .O(N__23497),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ));
    InMux I__2927 (
            .O(N__23494),
            .I(N__23490));
    InMux I__2926 (
            .O(N__23493),
            .I(N__23487));
    LocalMux I__2925 (
            .O(N__23490),
            .I(N__23484));
    LocalMux I__2924 (
            .O(N__23487),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    Odrv4 I__2923 (
            .O(N__23484),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    CascadeMux I__2922 (
            .O(N__23479),
            .I(N__23476));
    InMux I__2921 (
            .O(N__23476),
            .I(N__23473));
    LocalMux I__2920 (
            .O(N__23473),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11 ));
    InMux I__2919 (
            .O(N__23470),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ));
    CascadeMux I__2918 (
            .O(N__23467),
            .I(N__23463));
    InMux I__2917 (
            .O(N__23466),
            .I(N__23460));
    InMux I__2916 (
            .O(N__23463),
            .I(N__23457));
    LocalMux I__2915 (
            .O(N__23460),
            .I(N__23454));
    LocalMux I__2914 (
            .O(N__23457),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    Odrv4 I__2913 (
            .O(N__23454),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__2912 (
            .O(N__23449),
            .I(N__23446));
    LocalMux I__2911 (
            .O(N__23446),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12 ));
    InMux I__2910 (
            .O(N__23443),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ));
    InMux I__2909 (
            .O(N__23440),
            .I(N__23436));
    InMux I__2908 (
            .O(N__23439),
            .I(N__23433));
    LocalMux I__2907 (
            .O(N__23436),
            .I(N__23430));
    LocalMux I__2906 (
            .O(N__23433),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    Odrv4 I__2905 (
            .O(N__23430),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    CascadeMux I__2904 (
            .O(N__23425),
            .I(N__23422));
    InMux I__2903 (
            .O(N__23422),
            .I(N__23419));
    LocalMux I__2902 (
            .O(N__23419),
            .I(N__23416));
    Span4Mux_h I__2901 (
            .O(N__23416),
            .I(N__23413));
    Odrv4 I__2900 (
            .O(N__23413),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13 ));
    InMux I__2899 (
            .O(N__23410),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ));
    InMux I__2898 (
            .O(N__23407),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ));
    CascadeMux I__2897 (
            .O(N__23404),
            .I(N__23401));
    InMux I__2896 (
            .O(N__23401),
            .I(N__23398));
    LocalMux I__2895 (
            .O(N__23398),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ));
    CascadeMux I__2894 (
            .O(N__23395),
            .I(N__23392));
    InMux I__2893 (
            .O(N__23392),
            .I(N__23389));
    LocalMux I__2892 (
            .O(N__23389),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ));
    CascadeMux I__2891 (
            .O(N__23386),
            .I(N__23383));
    InMux I__2890 (
            .O(N__23383),
            .I(N__23380));
    LocalMux I__2889 (
            .O(N__23380),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ));
    CascadeMux I__2888 (
            .O(N__23377),
            .I(N__23372));
    InMux I__2887 (
            .O(N__23376),
            .I(N__23369));
    InMux I__2886 (
            .O(N__23375),
            .I(N__23366));
    InMux I__2885 (
            .O(N__23372),
            .I(N__23363));
    LocalMux I__2884 (
            .O(N__23369),
            .I(N__23360));
    LocalMux I__2883 (
            .O(N__23366),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__2882 (
            .O(N__23363),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv4 I__2881 (
            .O(N__23360),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    InMux I__2880 (
            .O(N__23353),
            .I(N__23350));
    LocalMux I__2879 (
            .O(N__23350),
            .I(N__23346));
    InMux I__2878 (
            .O(N__23349),
            .I(N__23343));
    Span4Mux_h I__2877 (
            .O(N__23346),
            .I(N__23340));
    LocalMux I__2876 (
            .O(N__23343),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    Odrv4 I__2875 (
            .O(N__23340),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__2874 (
            .O(N__23335),
            .I(N__23332));
    LocalMux I__2873 (
            .O(N__23332),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2 ));
    InMux I__2872 (
            .O(N__23329),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ));
    InMux I__2871 (
            .O(N__23326),
            .I(N__23322));
    CascadeMux I__2870 (
            .O(N__23325),
            .I(N__23319));
    LocalMux I__2869 (
            .O(N__23322),
            .I(N__23316));
    InMux I__2868 (
            .O(N__23319),
            .I(N__23313));
    Span4Mux_h I__2867 (
            .O(N__23316),
            .I(N__23310));
    LocalMux I__2866 (
            .O(N__23313),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    Odrv4 I__2865 (
            .O(N__23310),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__2864 (
            .O(N__23305),
            .I(N__23302));
    LocalMux I__2863 (
            .O(N__23302),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3 ));
    InMux I__2862 (
            .O(N__23299),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ));
    InMux I__2861 (
            .O(N__23296),
            .I(N__23293));
    LocalMux I__2860 (
            .O(N__23293),
            .I(N__23289));
    InMux I__2859 (
            .O(N__23292),
            .I(N__23286));
    Span4Mux_h I__2858 (
            .O(N__23289),
            .I(N__23283));
    LocalMux I__2857 (
            .O(N__23286),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    Odrv4 I__2856 (
            .O(N__23283),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__2855 (
            .O(N__23278),
            .I(N__23275));
    LocalMux I__2854 (
            .O(N__23275),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4 ));
    InMux I__2853 (
            .O(N__23272),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ));
    InMux I__2852 (
            .O(N__23269),
            .I(N__23265));
    InMux I__2851 (
            .O(N__23268),
            .I(N__23262));
    LocalMux I__2850 (
            .O(N__23265),
            .I(N__23257));
    LocalMux I__2849 (
            .O(N__23262),
            .I(N__23257));
    Span4Mux_v I__2848 (
            .O(N__23257),
            .I(N__23254));
    Odrv4 I__2847 (
            .O(N__23254),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__2846 (
            .O(N__23251),
            .I(N__23248));
    LocalMux I__2845 (
            .O(N__23248),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ));
    InMux I__2844 (
            .O(N__23245),
            .I(N__23242));
    LocalMux I__2843 (
            .O(N__23242),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ));
    InMux I__2842 (
            .O(N__23239),
            .I(N__23236));
    LocalMux I__2841 (
            .O(N__23236),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ));
    InMux I__2840 (
            .O(N__23233),
            .I(N__23230));
    LocalMux I__2839 (
            .O(N__23230),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ));
    CascadeMux I__2838 (
            .O(N__23227),
            .I(N__23224));
    InMux I__2837 (
            .O(N__23224),
            .I(N__23221));
    LocalMux I__2836 (
            .O(N__23221),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ));
    InMux I__2835 (
            .O(N__23218),
            .I(N__23215));
    LocalMux I__2834 (
            .O(N__23215),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_16 ));
    InMux I__2833 (
            .O(N__23212),
            .I(N__23209));
    LocalMux I__2832 (
            .O(N__23209),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_17 ));
    InMux I__2831 (
            .O(N__23206),
            .I(N__23203));
    LocalMux I__2830 (
            .O(N__23203),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_18 ));
    InMux I__2829 (
            .O(N__23200),
            .I(N__23197));
    LocalMux I__2828 (
            .O(N__23197),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_19 ));
    InMux I__2827 (
            .O(N__23194),
            .I(N__23191));
    LocalMux I__2826 (
            .O(N__23191),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ));
    InMux I__2825 (
            .O(N__23188),
            .I(N__23185));
    LocalMux I__2824 (
            .O(N__23185),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ));
    InMux I__2823 (
            .O(N__23182),
            .I(N__23179));
    LocalMux I__2822 (
            .O(N__23179),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ));
    InMux I__2821 (
            .O(N__23176),
            .I(N__23173));
    LocalMux I__2820 (
            .O(N__23173),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ));
    CascadeMux I__2819 (
            .O(N__23170),
            .I(N__23167));
    InMux I__2818 (
            .O(N__23167),
            .I(N__23164));
    LocalMux I__2817 (
            .O(N__23164),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ));
    InMux I__2816 (
            .O(N__23161),
            .I(N__23158));
    LocalMux I__2815 (
            .O(N__23158),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ));
    InMux I__2814 (
            .O(N__23155),
            .I(N__23152));
    LocalMux I__2813 (
            .O(N__23152),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ));
    InMux I__2812 (
            .O(N__23149),
            .I(N__23146));
    LocalMux I__2811 (
            .O(N__23146),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ));
    CascadeMux I__2810 (
            .O(N__23143),
            .I(N__23140));
    InMux I__2809 (
            .O(N__23140),
            .I(N__23137));
    LocalMux I__2808 (
            .O(N__23137),
            .I(N__23134));
    Odrv12 I__2807 (
            .O(N__23134),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ));
    InMux I__2806 (
            .O(N__23131),
            .I(N__23128));
    LocalMux I__2805 (
            .O(N__23128),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ));
    InMux I__2804 (
            .O(N__23125),
            .I(N__23122));
    LocalMux I__2803 (
            .O(N__23122),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_15 ));
    CascadeMux I__2802 (
            .O(N__23119),
            .I(N__23116));
    InMux I__2801 (
            .O(N__23116),
            .I(N__23113));
    LocalMux I__2800 (
            .O(N__23113),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_17 ));
    InMux I__2799 (
            .O(N__23110),
            .I(N__23107));
    LocalMux I__2798 (
            .O(N__23107),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_18 ));
    CascadeMux I__2797 (
            .O(N__23104),
            .I(N__23101));
    InMux I__2796 (
            .O(N__23101),
            .I(N__23098));
    LocalMux I__2795 (
            .O(N__23098),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_19 ));
    InMux I__2794 (
            .O(N__23095),
            .I(N__23092));
    LocalMux I__2793 (
            .O(N__23092),
            .I(N__23089));
    Span4Mux_h I__2792 (
            .O(N__23089),
            .I(N__23086));
    Odrv4 I__2791 (
            .O(N__23086),
            .I(\phase_controller_inst1.start_timer_hc_0_sqmuxa ));
    InMux I__2790 (
            .O(N__23083),
            .I(N__23080));
    LocalMux I__2789 (
            .O(N__23080),
            .I(\phase_controller_inst1.start_timer_hc_RNOZ0Z_0 ));
    CascadeMux I__2788 (
            .O(N__23077),
            .I(N__23074));
    InMux I__2787 (
            .O(N__23074),
            .I(N__23071));
    LocalMux I__2786 (
            .O(N__23071),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_9 ));
    InMux I__2785 (
            .O(N__23068),
            .I(N__23065));
    LocalMux I__2784 (
            .O(N__23065),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_16 ));
    InMux I__2783 (
            .O(N__23062),
            .I(N__23059));
    LocalMux I__2782 (
            .O(N__23059),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ));
    InMux I__2781 (
            .O(N__23056),
            .I(N__23053));
    LocalMux I__2780 (
            .O(N__23053),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ));
    InMux I__2779 (
            .O(N__23050),
            .I(N__23047));
    LocalMux I__2778 (
            .O(N__23047),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2 ));
    CascadeMux I__2777 (
            .O(N__23044),
            .I(\phase_controller_inst2.stoper_tr.time_passed11_cascade_ ));
    InMux I__2776 (
            .O(N__23041),
            .I(N__23038));
    LocalMux I__2775 (
            .O(N__23038),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNIF9HJZ0 ));
    InMux I__2774 (
            .O(N__23035),
            .I(N__23030));
    InMux I__2773 (
            .O(N__23034),
            .I(N__23027));
    InMux I__2772 (
            .O(N__23033),
            .I(N__23024));
    LocalMux I__2771 (
            .O(N__23030),
            .I(\phase_controller_inst2.stoper_tr.time_passed11 ));
    LocalMux I__2770 (
            .O(N__23027),
            .I(\phase_controller_inst2.stoper_tr.time_passed11 ));
    LocalMux I__2769 (
            .O(N__23024),
            .I(\phase_controller_inst2.stoper_tr.time_passed11 ));
    CascadeMux I__2768 (
            .O(N__23017),
            .I(N__23014));
    InMux I__2767 (
            .O(N__23014),
            .I(N__23011));
    LocalMux I__2766 (
            .O(N__23011),
            .I(N__23008));
    Odrv4 I__2765 (
            .O(N__23008),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_axb_0 ));
    CascadeMux I__2764 (
            .O(N__23005),
            .I(N__23002));
    InMux I__2763 (
            .O(N__23002),
            .I(N__22999));
    LocalMux I__2762 (
            .O(N__22999),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_10 ));
    InMux I__2761 (
            .O(N__22996),
            .I(N__22993));
    LocalMux I__2760 (
            .O(N__22993),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_11 ));
    CascadeMux I__2759 (
            .O(N__22990),
            .I(N__22987));
    InMux I__2758 (
            .O(N__22987),
            .I(N__22984));
    LocalMux I__2757 (
            .O(N__22984),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_12 ));
    InMux I__2756 (
            .O(N__22981),
            .I(N__22978));
    LocalMux I__2755 (
            .O(N__22978),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_13 ));
    CascadeMux I__2754 (
            .O(N__22975),
            .I(N__22972));
    InMux I__2753 (
            .O(N__22972),
            .I(N__22969));
    LocalMux I__2752 (
            .O(N__22969),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_14 ));
    CascadeMux I__2751 (
            .O(N__22966),
            .I(N__22963));
    InMux I__2750 (
            .O(N__22963),
            .I(N__22960));
    LocalMux I__2749 (
            .O(N__22960),
            .I(N__22957));
    Span4Mux_h I__2748 (
            .O(N__22957),
            .I(N__22954));
    Odrv4 I__2747 (
            .O(N__22954),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_7 ));
    InMux I__2746 (
            .O(N__22951),
            .I(N__22948));
    LocalMux I__2745 (
            .O(N__22948),
            .I(N__22945));
    Odrv4 I__2744 (
            .O(N__22945),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_3 ));
    InMux I__2743 (
            .O(N__22942),
            .I(N__22939));
    LocalMux I__2742 (
            .O(N__22939),
            .I(N__22936));
    Odrv4 I__2741 (
            .O(N__22936),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_2 ));
    InMux I__2740 (
            .O(N__22933),
            .I(N__22930));
    LocalMux I__2739 (
            .O(N__22930),
            .I(N__22927));
    Odrv4 I__2738 (
            .O(N__22927),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_8 ));
    CascadeMux I__2737 (
            .O(N__22924),
            .I(N__22921));
    InMux I__2736 (
            .O(N__22921),
            .I(N__22918));
    LocalMux I__2735 (
            .O(N__22918),
            .I(N__22915));
    Span4Mux_h I__2734 (
            .O(N__22915),
            .I(N__22912));
    Odrv4 I__2733 (
            .O(N__22912),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_6 ));
    InMux I__2732 (
            .O(N__22909),
            .I(N__22906));
    LocalMux I__2731 (
            .O(N__22906),
            .I(N__22903));
    Odrv4 I__2730 (
            .O(N__22903),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_5 ));
    CascadeMux I__2729 (
            .O(N__22900),
            .I(N__22897));
    InMux I__2728 (
            .O(N__22897),
            .I(N__22894));
    LocalMux I__2727 (
            .O(N__22894),
            .I(\phase_controller_inst2.stoper_tr.time_passed_1_sqmuxa ));
    CascadeMux I__2726 (
            .O(N__22891),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_ ));
    InMux I__2725 (
            .O(N__22888),
            .I(N__22885));
    LocalMux I__2724 (
            .O(N__22885),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ));
    InMux I__2723 (
            .O(N__22882),
            .I(N__22879));
    LocalMux I__2722 (
            .O(N__22879),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ));
    CascadeMux I__2721 (
            .O(N__22876),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ));
    InMux I__2720 (
            .O(N__22873),
            .I(N__22870));
    LocalMux I__2719 (
            .O(N__22870),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ));
    InMux I__2718 (
            .O(N__22867),
            .I(N__22864));
    LocalMux I__2717 (
            .O(N__22864),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ));
    InMux I__2716 (
            .O(N__22861),
            .I(N__22858));
    LocalMux I__2715 (
            .O(N__22858),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ));
    InMux I__2714 (
            .O(N__22855),
            .I(N__22852));
    LocalMux I__2713 (
            .O(N__22852),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9 ));
    InMux I__2712 (
            .O(N__22849),
            .I(N__22846));
    LocalMux I__2711 (
            .O(N__22846),
            .I(N__22843));
    Odrv4 I__2710 (
            .O(N__22843),
            .I(il_max_comp1_c));
    InMux I__2709 (
            .O(N__22840),
            .I(N__22837));
    LocalMux I__2708 (
            .O(N__22837),
            .I(il_max_comp1_D1));
    CascadeMux I__2707 (
            .O(N__22834),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_ ));
    InMux I__2706 (
            .O(N__22831),
            .I(N__22828));
    LocalMux I__2705 (
            .O(N__22828),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ));
    CascadeMux I__2704 (
            .O(N__22825),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_ ));
    CascadeMux I__2703 (
            .O(N__22822),
            .I(N__22817));
    InMux I__2702 (
            .O(N__22821),
            .I(N__22807));
    InMux I__2701 (
            .O(N__22820),
            .I(N__22807));
    InMux I__2700 (
            .O(N__22817),
            .I(N__22800));
    InMux I__2699 (
            .O(N__22816),
            .I(N__22800));
    InMux I__2698 (
            .O(N__22815),
            .I(N__22800));
    InMux I__2697 (
            .O(N__22814),
            .I(N__22797));
    InMux I__2696 (
            .O(N__22813),
            .I(N__22792));
    InMux I__2695 (
            .O(N__22812),
            .I(N__22792));
    LocalMux I__2694 (
            .O(N__22807),
            .I(N__22789));
    LocalMux I__2693 (
            .O(N__22800),
            .I(N__22786));
    LocalMux I__2692 (
            .O(N__22797),
            .I(N__22781));
    LocalMux I__2691 (
            .O(N__22792),
            .I(N__22781));
    Span4Mux_h I__2690 (
            .O(N__22789),
            .I(N__22778));
    Span4Mux_h I__2689 (
            .O(N__22786),
            .I(N__22775));
    Span4Mux_h I__2688 (
            .O(N__22781),
            .I(N__22772));
    Span4Mux_v I__2687 (
            .O(N__22778),
            .I(N__22769));
    Span4Mux_h I__2686 (
            .O(N__22775),
            .I(N__22766));
    Span4Mux_h I__2685 (
            .O(N__22772),
            .I(N__22763));
    Odrv4 I__2684 (
            .O(N__22769),
            .I(\current_shift_inst.PI_CTRL.N_53 ));
    Odrv4 I__2683 (
            .O(N__22766),
            .I(\current_shift_inst.PI_CTRL.N_53 ));
    Odrv4 I__2682 (
            .O(N__22763),
            .I(\current_shift_inst.PI_CTRL.N_53 ));
    InMux I__2681 (
            .O(N__22756),
            .I(N__22753));
    LocalMux I__2680 (
            .O(N__22753),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ));
    CascadeMux I__2679 (
            .O(N__22750),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9_cascade_ ));
    InMux I__2678 (
            .O(N__22747),
            .I(N__22735));
    InMux I__2677 (
            .O(N__22746),
            .I(N__22735));
    InMux I__2676 (
            .O(N__22745),
            .I(N__22735));
    InMux I__2675 (
            .O(N__22744),
            .I(N__22730));
    InMux I__2674 (
            .O(N__22743),
            .I(N__22730));
    InMux I__2673 (
            .O(N__22742),
            .I(N__22727));
    LocalMux I__2672 (
            .O(N__22735),
            .I(N__22723));
    LocalMux I__2671 (
            .O(N__22730),
            .I(N__22718));
    LocalMux I__2670 (
            .O(N__22727),
            .I(N__22718));
    InMux I__2669 (
            .O(N__22726),
            .I(N__22715));
    Span4Mux_h I__2668 (
            .O(N__22723),
            .I(N__22712));
    Sp12to4 I__2667 (
            .O(N__22718),
            .I(N__22707));
    LocalMux I__2666 (
            .O(N__22715),
            .I(N__22707));
    Span4Mux_h I__2665 (
            .O(N__22712),
            .I(N__22704));
    Span12Mux_s8_v I__2664 (
            .O(N__22707),
            .I(N__22701));
    Odrv4 I__2663 (
            .O(N__22704),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    Odrv12 I__2662 (
            .O(N__22701),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    InMux I__2661 (
            .O(N__22696),
            .I(N__22693));
    LocalMux I__2660 (
            .O(N__22693),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ));
    InMux I__2659 (
            .O(N__22690),
            .I(N__22687));
    LocalMux I__2658 (
            .O(N__22687),
            .I(N__22682));
    InMux I__2657 (
            .O(N__22686),
            .I(N__22679));
    CascadeMux I__2656 (
            .O(N__22685),
            .I(N__22676));
    Span12Mux_v I__2655 (
            .O(N__22682),
            .I(N__22670));
    LocalMux I__2654 (
            .O(N__22679),
            .I(N__22670));
    InMux I__2653 (
            .O(N__22676),
            .I(N__22667));
    InMux I__2652 (
            .O(N__22675),
            .I(N__22664));
    Odrv12 I__2651 (
            .O(N__22670),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    LocalMux I__2650 (
            .O(N__22667),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    LocalMux I__2649 (
            .O(N__22664),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    IoInMux I__2648 (
            .O(N__22657),
            .I(N__22654));
    LocalMux I__2647 (
            .O(N__22654),
            .I(N__22651));
    Span12Mux_s7_v I__2646 (
            .O(N__22651),
            .I(N__22648));
    Odrv12 I__2645 (
            .O(N__22648),
            .I(s4_phy_c));
    InMux I__2644 (
            .O(N__22645),
            .I(N__22642));
    LocalMux I__2643 (
            .O(N__22642),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0 ));
    InMux I__2642 (
            .O(N__22639),
            .I(bfn_7_17_0_));
    InMux I__2641 (
            .O(N__22636),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_16 ));
    InMux I__2640 (
            .O(N__22633),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_17 ));
    InMux I__2639 (
            .O(N__22630),
            .I(N__22626));
    CascadeMux I__2638 (
            .O(N__22629),
            .I(N__22622));
    LocalMux I__2637 (
            .O(N__22626),
            .I(N__22619));
    InMux I__2636 (
            .O(N__22625),
            .I(N__22616));
    InMux I__2635 (
            .O(N__22622),
            .I(N__22613));
    Span4Mux_h I__2634 (
            .O(N__22619),
            .I(N__22610));
    LocalMux I__2633 (
            .O(N__22616),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    LocalMux I__2632 (
            .O(N__22613),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    Odrv4 I__2631 (
            .O(N__22610),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    CascadeMux I__2630 (
            .O(N__22603),
            .I(N__22600));
    InMux I__2629 (
            .O(N__22600),
            .I(N__22597));
    LocalMux I__2628 (
            .O(N__22597),
            .I(N__22594));
    Odrv4 I__2627 (
            .O(N__22594),
            .I(\phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa ));
    InMux I__2626 (
            .O(N__22591),
            .I(N__22588));
    LocalMux I__2625 (
            .O(N__22588),
            .I(N__22584));
    InMux I__2624 (
            .O(N__22587),
            .I(N__22581));
    Span4Mux_h I__2623 (
            .O(N__22584),
            .I(N__22575));
    LocalMux I__2622 (
            .O(N__22581),
            .I(N__22575));
    InMux I__2621 (
            .O(N__22580),
            .I(N__22572));
    Span4Mux_v I__2620 (
            .O(N__22575),
            .I(N__22569));
    LocalMux I__2619 (
            .O(N__22572),
            .I(N__22566));
    Span4Mux_v I__2618 (
            .O(N__22569),
            .I(N__22563));
    Odrv12 I__2617 (
            .O(N__22566),
            .I(il_min_comp1_D2));
    Odrv4 I__2616 (
            .O(N__22563),
            .I(il_min_comp1_D2));
    InMux I__2615 (
            .O(N__22558),
            .I(N__22553));
    InMux I__2614 (
            .O(N__22557),
            .I(N__22550));
    InMux I__2613 (
            .O(N__22556),
            .I(N__22547));
    LocalMux I__2612 (
            .O(N__22553),
            .I(N__22544));
    LocalMux I__2611 (
            .O(N__22550),
            .I(\phase_controller_inst1.tr_time_passed ));
    LocalMux I__2610 (
            .O(N__22547),
            .I(\phase_controller_inst1.tr_time_passed ));
    Odrv4 I__2609 (
            .O(N__22544),
            .I(\phase_controller_inst1.tr_time_passed ));
    InMux I__2608 (
            .O(N__22537),
            .I(N__22533));
    InMux I__2607 (
            .O(N__22536),
            .I(N__22530));
    LocalMux I__2606 (
            .O(N__22533),
            .I(N__22527));
    LocalMux I__2605 (
            .O(N__22530),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    Odrv4 I__2604 (
            .O(N__22527),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    InMux I__2603 (
            .O(N__22522),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_6 ));
    InMux I__2602 (
            .O(N__22519),
            .I(bfn_7_16_0_));
    InMux I__2601 (
            .O(N__22516),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_8 ));
    InMux I__2600 (
            .O(N__22513),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_9 ));
    InMux I__2599 (
            .O(N__22510),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_10 ));
    InMux I__2598 (
            .O(N__22507),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_11 ));
    InMux I__2597 (
            .O(N__22504),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_12 ));
    InMux I__2596 (
            .O(N__22501),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_13 ));
    InMux I__2595 (
            .O(N__22498),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_14 ));
    CascadeMux I__2594 (
            .O(N__22495),
            .I(\phase_controller_inst2.state_RNI9M3OZ0Z_0_cascade_ ));
    CascadeMux I__2593 (
            .O(N__22492),
            .I(N__22488));
    InMux I__2592 (
            .O(N__22491),
            .I(N__22485));
    InMux I__2591 (
            .O(N__22488),
            .I(N__22482));
    LocalMux I__2590 (
            .O(N__22485),
            .I(N__22479));
    LocalMux I__2589 (
            .O(N__22482),
            .I(N__22476));
    Odrv4 I__2588 (
            .O(N__22479),
            .I(state_ns_i_a3_1));
    Odrv12 I__2587 (
            .O(N__22476),
            .I(state_ns_i_a3_1));
    InMux I__2586 (
            .O(N__22471),
            .I(N__22466));
    InMux I__2585 (
            .O(N__22470),
            .I(N__22463));
    InMux I__2584 (
            .O(N__22469),
            .I(N__22460));
    LocalMux I__2583 (
            .O(N__22466),
            .I(N__22453));
    LocalMux I__2582 (
            .O(N__22463),
            .I(N__22453));
    LocalMux I__2581 (
            .O(N__22460),
            .I(N__22453));
    Odrv12 I__2580 (
            .O(N__22453),
            .I(il_min_comp2_D2));
    CascadeMux I__2579 (
            .O(N__22450),
            .I(N__22447));
    InMux I__2578 (
            .O(N__22447),
            .I(N__22440));
    InMux I__2577 (
            .O(N__22446),
            .I(N__22440));
    InMux I__2576 (
            .O(N__22445),
            .I(N__22437));
    LocalMux I__2575 (
            .O(N__22440),
            .I(\phase_controller_inst2.tr_time_passed ));
    LocalMux I__2574 (
            .O(N__22437),
            .I(\phase_controller_inst2.tr_time_passed ));
    InMux I__2573 (
            .O(N__22432),
            .I(N__22426));
    InMux I__2572 (
            .O(N__22431),
            .I(N__22426));
    LocalMux I__2571 (
            .O(N__22426),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    InMux I__2570 (
            .O(N__22423),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0 ));
    InMux I__2569 (
            .O(N__22420),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_1 ));
    InMux I__2568 (
            .O(N__22417),
            .I(N__22414));
    LocalMux I__2567 (
            .O(N__22414),
            .I(N__22411));
    Odrv4 I__2566 (
            .O(N__22411),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_4 ));
    InMux I__2565 (
            .O(N__22408),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_2 ));
    InMux I__2564 (
            .O(N__22405),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_3 ));
    InMux I__2563 (
            .O(N__22402),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_4 ));
    InMux I__2562 (
            .O(N__22399),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_5 ));
    InMux I__2561 (
            .O(N__22396),
            .I(N__22393));
    LocalMux I__2560 (
            .O(N__22393),
            .I(N__22390));
    Span4Mux_h I__2559 (
            .O(N__22390),
            .I(N__22387));
    Span4Mux_v I__2558 (
            .O(N__22387),
            .I(N__22384));
    Odrv4 I__2557 (
            .O(N__22384),
            .I(il_max_comp2_c));
    InMux I__2556 (
            .O(N__22381),
            .I(N__22378));
    LocalMux I__2555 (
            .O(N__22378),
            .I(N__22375));
    Odrv4 I__2554 (
            .O(N__22375),
            .I(il_max_comp2_D1));
    IoInMux I__2553 (
            .O(N__22372),
            .I(N__22369));
    LocalMux I__2552 (
            .O(N__22369),
            .I(N__22366));
    IoSpan4Mux I__2551 (
            .O(N__22366),
            .I(N__22363));
    Span4Mux_s1_v I__2550 (
            .O(N__22363),
            .I(N__22360));
    Sp12to4 I__2549 (
            .O(N__22360),
            .I(N__22357));
    Span12Mux_s9_v I__2548 (
            .O(N__22357),
            .I(N__22354));
    Odrv12 I__2547 (
            .O(N__22354),
            .I(\delay_measurement_inst.delay_hc_timer.N_302_i ));
    CascadeMux I__2546 (
            .O(N__22351),
            .I(N__22348));
    InMux I__2545 (
            .O(N__22348),
            .I(N__22345));
    LocalMux I__2544 (
            .O(N__22345),
            .I(\phase_controller_inst2.start_timer_tr_0_sqmuxa ));
    InMux I__2543 (
            .O(N__22342),
            .I(N__22339));
    LocalMux I__2542 (
            .O(N__22339),
            .I(N__22336));
    Odrv4 I__2541 (
            .O(N__22336),
            .I(\phase_controller_inst2.state_RNI9M3OZ0Z_0 ));
    InMux I__2540 (
            .O(N__22333),
            .I(N__22329));
    InMux I__2539 (
            .O(N__22332),
            .I(N__22326));
    LocalMux I__2538 (
            .O(N__22329),
            .I(N__22321));
    LocalMux I__2537 (
            .O(N__22326),
            .I(N__22321));
    Span4Mux_s3_v I__2536 (
            .O(N__22321),
            .I(N__22318));
    Span4Mux_h I__2535 (
            .O(N__22318),
            .I(N__22313));
    InMux I__2534 (
            .O(N__22317),
            .I(N__22310));
    InMux I__2533 (
            .O(N__22316),
            .I(N__22307));
    Sp12to4 I__2532 (
            .O(N__22313),
            .I(N__22304));
    LocalMux I__2531 (
            .O(N__22310),
            .I(N__22299));
    LocalMux I__2530 (
            .O(N__22307),
            .I(N__22299));
    Span12Mux_v I__2529 (
            .O(N__22304),
            .I(N__22294));
    Sp12to4 I__2528 (
            .O(N__22299),
            .I(N__22294));
    Span12Mux_v I__2527 (
            .O(N__22294),
            .I(N__22291));
    Span12Mux_h I__2526 (
            .O(N__22291),
            .I(N__22288));
    Odrv12 I__2525 (
            .O(N__22288),
            .I(start_stop_c));
    CascadeMux I__2524 (
            .O(N__22285),
            .I(N__22282));
    InMux I__2523 (
            .O(N__22282),
            .I(N__22279));
    LocalMux I__2522 (
            .O(N__22279),
            .I(\phase_controller_inst1.start_timer_tr_0_sqmuxa ));
    InMux I__2521 (
            .O(N__22276),
            .I(N__22273));
    LocalMux I__2520 (
            .O(N__22273),
            .I(N__22269));
    InMux I__2519 (
            .O(N__22272),
            .I(N__22266));
    Odrv4 I__2518 (
            .O(N__22269),
            .I(\phase_controller_inst1.state_RNI7NN7Z0Z_0 ));
    LocalMux I__2517 (
            .O(N__22266),
            .I(\phase_controller_inst1.state_RNI7NN7Z0Z_0 ));
    InMux I__2516 (
            .O(N__22261),
            .I(N__22254));
    InMux I__2515 (
            .O(N__22260),
            .I(N__22254));
    InMux I__2514 (
            .O(N__22259),
            .I(N__22251));
    LocalMux I__2513 (
            .O(N__22254),
            .I(N__22248));
    LocalMux I__2512 (
            .O(N__22251),
            .I(N__22245));
    Span4Mux_h I__2511 (
            .O(N__22248),
            .I(N__22242));
    Span4Mux_h I__2510 (
            .O(N__22245),
            .I(N__22239));
    Sp12to4 I__2509 (
            .O(N__22242),
            .I(N__22236));
    Span4Mux_v I__2508 (
            .O(N__22239),
            .I(N__22233));
    Span12Mux_v I__2507 (
            .O(N__22236),
            .I(N__22230));
    Span4Mux_v I__2506 (
            .O(N__22233),
            .I(N__22227));
    Odrv12 I__2505 (
            .O(N__22230),
            .I(il_max_comp1_D2));
    Odrv4 I__2504 (
            .O(N__22227),
            .I(il_max_comp1_D2));
    InMux I__2503 (
            .O(N__22222),
            .I(N__22219));
    LocalMux I__2502 (
            .O(N__22219),
            .I(N__22216));
    Odrv12 I__2501 (
            .O(N__22216),
            .I(il_min_comp2_c));
    InMux I__2500 (
            .O(N__22213),
            .I(N__22210));
    LocalMux I__2499 (
            .O(N__22210),
            .I(il_min_comp2_D1));
    CascadeMux I__2498 (
            .O(N__22207),
            .I(N__22204));
    InMux I__2497 (
            .O(N__22204),
            .I(N__22201));
    LocalMux I__2496 (
            .O(N__22201),
            .I(\pwm_generator_inst.thresholdZ0Z_5 ));
    InMux I__2495 (
            .O(N__22198),
            .I(N__22193));
    InMux I__2494 (
            .O(N__22197),
            .I(N__22190));
    InMux I__2493 (
            .O(N__22196),
            .I(N__22187));
    LocalMux I__2492 (
            .O(N__22193),
            .I(N__22182));
    LocalMux I__2491 (
            .O(N__22190),
            .I(N__22182));
    LocalMux I__2490 (
            .O(N__22187),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    Odrv4 I__2489 (
            .O(N__22182),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    InMux I__2488 (
            .O(N__22177),
            .I(N__22174));
    LocalMux I__2487 (
            .O(N__22174),
            .I(\pwm_generator_inst.counter_i_5 ));
    InMux I__2486 (
            .O(N__22171),
            .I(N__22166));
    InMux I__2485 (
            .O(N__22170),
            .I(N__22163));
    InMux I__2484 (
            .O(N__22169),
            .I(N__22160));
    LocalMux I__2483 (
            .O(N__22166),
            .I(N__22155));
    LocalMux I__2482 (
            .O(N__22163),
            .I(N__22155));
    LocalMux I__2481 (
            .O(N__22160),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    Odrv4 I__2480 (
            .O(N__22155),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    CascadeMux I__2479 (
            .O(N__22150),
            .I(N__22147));
    InMux I__2478 (
            .O(N__22147),
            .I(N__22144));
    LocalMux I__2477 (
            .O(N__22144),
            .I(\pwm_generator_inst.thresholdZ0Z_6 ));
    InMux I__2476 (
            .O(N__22141),
            .I(N__22138));
    LocalMux I__2475 (
            .O(N__22138),
            .I(\pwm_generator_inst.counter_i_6 ));
    CascadeMux I__2474 (
            .O(N__22135),
            .I(N__22132));
    InMux I__2473 (
            .O(N__22132),
            .I(N__22129));
    LocalMux I__2472 (
            .O(N__22129),
            .I(\pwm_generator_inst.thresholdZ0Z_7 ));
    InMux I__2471 (
            .O(N__22126),
            .I(N__22121));
    InMux I__2470 (
            .O(N__22125),
            .I(N__22118));
    InMux I__2469 (
            .O(N__22124),
            .I(N__22115));
    LocalMux I__2468 (
            .O(N__22121),
            .I(N__22112));
    LocalMux I__2467 (
            .O(N__22118),
            .I(N__22109));
    LocalMux I__2466 (
            .O(N__22115),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    Odrv4 I__2465 (
            .O(N__22112),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    Odrv4 I__2464 (
            .O(N__22109),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    InMux I__2463 (
            .O(N__22102),
            .I(N__22099));
    LocalMux I__2462 (
            .O(N__22099),
            .I(\pwm_generator_inst.counter_i_7 ));
    CascadeMux I__2461 (
            .O(N__22096),
            .I(N__22093));
    InMux I__2460 (
            .O(N__22093),
            .I(N__22090));
    LocalMux I__2459 (
            .O(N__22090),
            .I(N__22087));
    Span4Mux_h I__2458 (
            .O(N__22087),
            .I(N__22084));
    Odrv4 I__2457 (
            .O(N__22084),
            .I(\pwm_generator_inst.thresholdZ0Z_8 ));
    InMux I__2456 (
            .O(N__22081),
            .I(N__22076));
    InMux I__2455 (
            .O(N__22080),
            .I(N__22073));
    InMux I__2454 (
            .O(N__22079),
            .I(N__22070));
    LocalMux I__2453 (
            .O(N__22076),
            .I(N__22067));
    LocalMux I__2452 (
            .O(N__22073),
            .I(N__22064));
    LocalMux I__2451 (
            .O(N__22070),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    Odrv12 I__2450 (
            .O(N__22067),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    Odrv4 I__2449 (
            .O(N__22064),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    InMux I__2448 (
            .O(N__22057),
            .I(N__22054));
    LocalMux I__2447 (
            .O(N__22054),
            .I(\pwm_generator_inst.counter_i_8 ));
    CascadeMux I__2446 (
            .O(N__22051),
            .I(N__22048));
    InMux I__2445 (
            .O(N__22048),
            .I(N__22045));
    LocalMux I__2444 (
            .O(N__22045),
            .I(\pwm_generator_inst.thresholdZ0Z_9 ));
    InMux I__2443 (
            .O(N__22042),
            .I(N__22037));
    InMux I__2442 (
            .O(N__22041),
            .I(N__22034));
    InMux I__2441 (
            .O(N__22040),
            .I(N__22031));
    LocalMux I__2440 (
            .O(N__22037),
            .I(N__22028));
    LocalMux I__2439 (
            .O(N__22034),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    LocalMux I__2438 (
            .O(N__22031),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    Odrv12 I__2437 (
            .O(N__22028),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    InMux I__2436 (
            .O(N__22021),
            .I(N__22018));
    LocalMux I__2435 (
            .O(N__22018),
            .I(\pwm_generator_inst.counter_i_9 ));
    InMux I__2434 (
            .O(N__22015),
            .I(\pwm_generator_inst.un14_counter_cry_9 ));
    IoInMux I__2433 (
            .O(N__22012),
            .I(N__22009));
    LocalMux I__2432 (
            .O(N__22009),
            .I(N__22006));
    Span4Mux_s1_v I__2431 (
            .O(N__22006),
            .I(N__22003));
    Span4Mux_h I__2430 (
            .O(N__22003),
            .I(N__22000));
    Sp12to4 I__2429 (
            .O(N__22000),
            .I(N__21997));
    Span12Mux_h I__2428 (
            .O(N__21997),
            .I(N__21994));
    Odrv12 I__2427 (
            .O(N__21994),
            .I(pwm_output_c));
    CascadeMux I__2426 (
            .O(N__21991),
            .I(\pwm_generator_inst.un1_counterlto9_2_cascade_ ));
    InMux I__2425 (
            .O(N__21988),
            .I(N__21970));
    InMux I__2424 (
            .O(N__21987),
            .I(N__21970));
    InMux I__2423 (
            .O(N__21986),
            .I(N__21970));
    InMux I__2422 (
            .O(N__21985),
            .I(N__21970));
    InMux I__2421 (
            .O(N__21984),
            .I(N__21961));
    InMux I__2420 (
            .O(N__21983),
            .I(N__21961));
    InMux I__2419 (
            .O(N__21982),
            .I(N__21961));
    InMux I__2418 (
            .O(N__21981),
            .I(N__21961));
    InMux I__2417 (
            .O(N__21980),
            .I(N__21956));
    InMux I__2416 (
            .O(N__21979),
            .I(N__21956));
    LocalMux I__2415 (
            .O(N__21970),
            .I(N__21951));
    LocalMux I__2414 (
            .O(N__21961),
            .I(N__21951));
    LocalMux I__2413 (
            .O(N__21956),
            .I(\pwm_generator_inst.un1_counter_0 ));
    Odrv4 I__2412 (
            .O(N__21951),
            .I(\pwm_generator_inst.un1_counter_0 ));
    CascadeMux I__2411 (
            .O(N__21946),
            .I(\pwm_generator_inst.un1_counterlto2_0_cascade_ ));
    InMux I__2410 (
            .O(N__21943),
            .I(N__21940));
    LocalMux I__2409 (
            .O(N__21940),
            .I(\pwm_generator_inst.un1_counterlt9 ));
    CascadeMux I__2408 (
            .O(N__21937),
            .I(N__21934));
    InMux I__2407 (
            .O(N__21934),
            .I(N__21931));
    LocalMux I__2406 (
            .O(N__21931),
            .I(N__21928));
    Odrv4 I__2405 (
            .O(N__21928),
            .I(\pwm_generator_inst.thresholdZ0Z_0 ));
    InMux I__2404 (
            .O(N__21925),
            .I(N__21920));
    InMux I__2403 (
            .O(N__21924),
            .I(N__21917));
    InMux I__2402 (
            .O(N__21923),
            .I(N__21914));
    LocalMux I__2401 (
            .O(N__21920),
            .I(N__21911));
    LocalMux I__2400 (
            .O(N__21917),
            .I(N__21908));
    LocalMux I__2399 (
            .O(N__21914),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    Odrv12 I__2398 (
            .O(N__21911),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    Odrv4 I__2397 (
            .O(N__21908),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    InMux I__2396 (
            .O(N__21901),
            .I(N__21898));
    LocalMux I__2395 (
            .O(N__21898),
            .I(\pwm_generator_inst.counter_i_0 ));
    CascadeMux I__2394 (
            .O(N__21895),
            .I(N__21892));
    InMux I__2393 (
            .O(N__21892),
            .I(N__21889));
    LocalMux I__2392 (
            .O(N__21889),
            .I(\pwm_generator_inst.thresholdZ0Z_1 ));
    InMux I__2391 (
            .O(N__21886),
            .I(N__21881));
    InMux I__2390 (
            .O(N__21885),
            .I(N__21878));
    InMux I__2389 (
            .O(N__21884),
            .I(N__21875));
    LocalMux I__2388 (
            .O(N__21881),
            .I(N__21872));
    LocalMux I__2387 (
            .O(N__21878),
            .I(N__21869));
    LocalMux I__2386 (
            .O(N__21875),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    Odrv12 I__2385 (
            .O(N__21872),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    Odrv4 I__2384 (
            .O(N__21869),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    InMux I__2383 (
            .O(N__21862),
            .I(N__21859));
    LocalMux I__2382 (
            .O(N__21859),
            .I(\pwm_generator_inst.counter_i_1 ));
    CascadeMux I__2381 (
            .O(N__21856),
            .I(N__21853));
    InMux I__2380 (
            .O(N__21853),
            .I(N__21850));
    LocalMux I__2379 (
            .O(N__21850),
            .I(\pwm_generator_inst.thresholdZ0Z_2 ));
    InMux I__2378 (
            .O(N__21847),
            .I(N__21842));
    InMux I__2377 (
            .O(N__21846),
            .I(N__21839));
    InMux I__2376 (
            .O(N__21845),
            .I(N__21836));
    LocalMux I__2375 (
            .O(N__21842),
            .I(N__21831));
    LocalMux I__2374 (
            .O(N__21839),
            .I(N__21831));
    LocalMux I__2373 (
            .O(N__21836),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    Odrv4 I__2372 (
            .O(N__21831),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    InMux I__2371 (
            .O(N__21826),
            .I(N__21823));
    LocalMux I__2370 (
            .O(N__21823),
            .I(\pwm_generator_inst.counter_i_2 ));
    CascadeMux I__2369 (
            .O(N__21820),
            .I(N__21817));
    InMux I__2368 (
            .O(N__21817),
            .I(N__21814));
    LocalMux I__2367 (
            .O(N__21814),
            .I(\pwm_generator_inst.thresholdZ0Z_3 ));
    InMux I__2366 (
            .O(N__21811),
            .I(N__21806));
    InMux I__2365 (
            .O(N__21810),
            .I(N__21803));
    InMux I__2364 (
            .O(N__21809),
            .I(N__21800));
    LocalMux I__2363 (
            .O(N__21806),
            .I(N__21795));
    LocalMux I__2362 (
            .O(N__21803),
            .I(N__21795));
    LocalMux I__2361 (
            .O(N__21800),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    Odrv4 I__2360 (
            .O(N__21795),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    InMux I__2359 (
            .O(N__21790),
            .I(N__21787));
    LocalMux I__2358 (
            .O(N__21787),
            .I(N__21784));
    Odrv4 I__2357 (
            .O(N__21784),
            .I(\pwm_generator_inst.counter_i_3 ));
    CascadeMux I__2356 (
            .O(N__21781),
            .I(N__21778));
    InMux I__2355 (
            .O(N__21778),
            .I(N__21775));
    LocalMux I__2354 (
            .O(N__21775),
            .I(N__21772));
    Span4Mux_h I__2353 (
            .O(N__21772),
            .I(N__21769));
    Odrv4 I__2352 (
            .O(N__21769),
            .I(\pwm_generator_inst.thresholdZ0Z_4 ));
    InMux I__2351 (
            .O(N__21766),
            .I(N__21761));
    InMux I__2350 (
            .O(N__21765),
            .I(N__21758));
    InMux I__2349 (
            .O(N__21764),
            .I(N__21755));
    LocalMux I__2348 (
            .O(N__21761),
            .I(N__21750));
    LocalMux I__2347 (
            .O(N__21758),
            .I(N__21750));
    LocalMux I__2346 (
            .O(N__21755),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    Odrv4 I__2345 (
            .O(N__21750),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    InMux I__2344 (
            .O(N__21745),
            .I(N__21742));
    LocalMux I__2343 (
            .O(N__21742),
            .I(\pwm_generator_inst.counter_i_4 ));
    InMux I__2342 (
            .O(N__21739),
            .I(\pwm_generator_inst.counter_cry_2 ));
    InMux I__2341 (
            .O(N__21736),
            .I(\pwm_generator_inst.counter_cry_3 ));
    InMux I__2340 (
            .O(N__21733),
            .I(\pwm_generator_inst.counter_cry_4 ));
    InMux I__2339 (
            .O(N__21730),
            .I(\pwm_generator_inst.counter_cry_5 ));
    InMux I__2338 (
            .O(N__21727),
            .I(\pwm_generator_inst.counter_cry_6 ));
    InMux I__2337 (
            .O(N__21724),
            .I(bfn_5_9_0_));
    InMux I__2336 (
            .O(N__21721),
            .I(\pwm_generator_inst.counter_cry_8 ));
    InMux I__2335 (
            .O(N__21718),
            .I(N__21715));
    LocalMux I__2334 (
            .O(N__21715),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_0 ));
    InMux I__2333 (
            .O(N__21712),
            .I(N__21709));
    LocalMux I__2332 (
            .O(N__21709),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_7 ));
    InMux I__2331 (
            .O(N__21706),
            .I(N__21703));
    LocalMux I__2330 (
            .O(N__21703),
            .I(N__21700));
    Odrv4 I__2329 (
            .O(N__21700),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_5 ));
    InMux I__2328 (
            .O(N__21697),
            .I(N__21694));
    LocalMux I__2327 (
            .O(N__21694),
            .I(N__21691));
    Odrv4 I__2326 (
            .O(N__21691),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_2 ));
    InMux I__2325 (
            .O(N__21688),
            .I(N__21685));
    LocalMux I__2324 (
            .O(N__21685),
            .I(N__21682));
    Odrv4 I__2323 (
            .O(N__21682),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_3 ));
    InMux I__2322 (
            .O(N__21679),
            .I(N__21676));
    LocalMux I__2321 (
            .O(N__21676),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_9 ));
    InMux I__2320 (
            .O(N__21673),
            .I(bfn_5_8_0_));
    InMux I__2319 (
            .O(N__21670),
            .I(\pwm_generator_inst.counter_cry_0 ));
    InMux I__2318 (
            .O(N__21667),
            .I(\pwm_generator_inst.counter_cry_1 ));
    InMux I__2317 (
            .O(N__21664),
            .I(N__21661));
    LocalMux I__2316 (
            .O(N__21661),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3 ));
    InMux I__2315 (
            .O(N__21658),
            .I(N__21655));
    LocalMux I__2314 (
            .O(N__21655),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0 ));
    InMux I__2313 (
            .O(N__21652),
            .I(N__21649));
    LocalMux I__2312 (
            .O(N__21649),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7 ));
    InMux I__2311 (
            .O(N__21646),
            .I(N__21643));
    LocalMux I__2310 (
            .O(N__21643),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6 ));
    InMux I__2309 (
            .O(N__21640),
            .I(N__21637));
    LocalMux I__2308 (
            .O(N__21637),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1 ));
    InMux I__2307 (
            .O(N__21634),
            .I(N__21631));
    LocalMux I__2306 (
            .O(N__21631),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5 ));
    CascadeMux I__2305 (
            .O(N__21628),
            .I(N__21621));
    CascadeMux I__2304 (
            .O(N__21627),
            .I(N__21617));
    CascadeMux I__2303 (
            .O(N__21626),
            .I(N__21614));
    InMux I__2302 (
            .O(N__21625),
            .I(N__21589));
    InMux I__2301 (
            .O(N__21624),
            .I(N__21589));
    InMux I__2300 (
            .O(N__21621),
            .I(N__21586));
    InMux I__2299 (
            .O(N__21620),
            .I(N__21583));
    InMux I__2298 (
            .O(N__21617),
            .I(N__21578));
    InMux I__2297 (
            .O(N__21614),
            .I(N__21578));
    InMux I__2296 (
            .O(N__21613),
            .I(N__21569));
    InMux I__2295 (
            .O(N__21612),
            .I(N__21569));
    InMux I__2294 (
            .O(N__21611),
            .I(N__21569));
    InMux I__2293 (
            .O(N__21610),
            .I(N__21569));
    InMux I__2292 (
            .O(N__21609),
            .I(N__21551));
    InMux I__2291 (
            .O(N__21608),
            .I(N__21551));
    InMux I__2290 (
            .O(N__21607),
            .I(N__21551));
    InMux I__2289 (
            .O(N__21606),
            .I(N__21551));
    InMux I__2288 (
            .O(N__21605),
            .I(N__21551));
    InMux I__2287 (
            .O(N__21604),
            .I(N__21551));
    InMux I__2286 (
            .O(N__21603),
            .I(N__21551));
    InMux I__2285 (
            .O(N__21602),
            .I(N__21551));
    InMux I__2284 (
            .O(N__21601),
            .I(N__21548));
    InMux I__2283 (
            .O(N__21600),
            .I(N__21533));
    InMux I__2282 (
            .O(N__21599),
            .I(N__21533));
    InMux I__2281 (
            .O(N__21598),
            .I(N__21533));
    InMux I__2280 (
            .O(N__21597),
            .I(N__21533));
    InMux I__2279 (
            .O(N__21596),
            .I(N__21533));
    InMux I__2278 (
            .O(N__21595),
            .I(N__21533));
    InMux I__2277 (
            .O(N__21594),
            .I(N__21533));
    LocalMux I__2276 (
            .O(N__21589),
            .I(N__21530));
    LocalMux I__2275 (
            .O(N__21586),
            .I(N__21521));
    LocalMux I__2274 (
            .O(N__21583),
            .I(N__21521));
    LocalMux I__2273 (
            .O(N__21578),
            .I(N__21521));
    LocalMux I__2272 (
            .O(N__21569),
            .I(N__21521));
    InMux I__2271 (
            .O(N__21568),
            .I(N__21518));
    LocalMux I__2270 (
            .O(N__21551),
            .I(N__21515));
    LocalMux I__2269 (
            .O(N__21548),
            .I(N__21510));
    LocalMux I__2268 (
            .O(N__21533),
            .I(N__21510));
    Span4Mux_v I__2267 (
            .O(N__21530),
            .I(N__21500));
    Span4Mux_v I__2266 (
            .O(N__21521),
            .I(N__21500));
    LocalMux I__2265 (
            .O(N__21518),
            .I(N__21497));
    Span4Mux_v I__2264 (
            .O(N__21515),
            .I(N__21492));
    Span4Mux_v I__2263 (
            .O(N__21510),
            .I(N__21492));
    InMux I__2262 (
            .O(N__21509),
            .I(N__21487));
    InMux I__2261 (
            .O(N__21508),
            .I(N__21487));
    InMux I__2260 (
            .O(N__21507),
            .I(N__21480));
    InMux I__2259 (
            .O(N__21506),
            .I(N__21480));
    InMux I__2258 (
            .O(N__21505),
            .I(N__21480));
    Odrv4 I__2257 (
            .O(N__21500),
            .I(N_19_1));
    Odrv12 I__2256 (
            .O(N__21497),
            .I(N_19_1));
    Odrv4 I__2255 (
            .O(N__21492),
            .I(N_19_1));
    LocalMux I__2254 (
            .O(N__21487),
            .I(N_19_1));
    LocalMux I__2253 (
            .O(N__21480),
            .I(N_19_1));
    InMux I__2252 (
            .O(N__21469),
            .I(N__21448));
    InMux I__2251 (
            .O(N__21468),
            .I(N__21448));
    InMux I__2250 (
            .O(N__21467),
            .I(N__21448));
    InMux I__2249 (
            .O(N__21466),
            .I(N__21448));
    InMux I__2248 (
            .O(N__21465),
            .I(N__21448));
    InMux I__2247 (
            .O(N__21464),
            .I(N__21448));
    CascadeMux I__2246 (
            .O(N__21463),
            .I(N__21445));
    InMux I__2245 (
            .O(N__21462),
            .I(N__21439));
    InMux I__2244 (
            .O(N__21461),
            .I(N__21439));
    LocalMux I__2243 (
            .O(N__21448),
            .I(N__21436));
    InMux I__2242 (
            .O(N__21445),
            .I(N__21431));
    InMux I__2241 (
            .O(N__21444),
            .I(N__21431));
    LocalMux I__2240 (
            .O(N__21439),
            .I(N__21428));
    Span4Mux_v I__2239 (
            .O(N__21436),
            .I(N__21423));
    LocalMux I__2238 (
            .O(N__21431),
            .I(N__21423));
    Odrv12 I__2237 (
            .O(N__21428),
            .I(\pwm_generator_inst.N_16 ));
    Odrv4 I__2236 (
            .O(N__21423),
            .I(\pwm_generator_inst.N_16 ));
    CascadeMux I__2235 (
            .O(N__21418),
            .I(N__21410));
    CascadeMux I__2234 (
            .O(N__21417),
            .I(N__21407));
    CascadeMux I__2233 (
            .O(N__21416),
            .I(N__21402));
    CascadeMux I__2232 (
            .O(N__21415),
            .I(N__21399));
    CascadeMux I__2231 (
            .O(N__21414),
            .I(N__21396));
    InMux I__2230 (
            .O(N__21413),
            .I(N__21389));
    InMux I__2229 (
            .O(N__21410),
            .I(N__21389));
    InMux I__2228 (
            .O(N__21407),
            .I(N__21376));
    InMux I__2227 (
            .O(N__21406),
            .I(N__21376));
    InMux I__2226 (
            .O(N__21405),
            .I(N__21376));
    InMux I__2225 (
            .O(N__21402),
            .I(N__21376));
    InMux I__2224 (
            .O(N__21399),
            .I(N__21376));
    InMux I__2223 (
            .O(N__21396),
            .I(N__21376));
    InMux I__2222 (
            .O(N__21395),
            .I(N__21371));
    InMux I__2221 (
            .O(N__21394),
            .I(N__21371));
    LocalMux I__2220 (
            .O(N__21389),
            .I(N__21368));
    LocalMux I__2219 (
            .O(N__21376),
            .I(N__21363));
    LocalMux I__2218 (
            .O(N__21371),
            .I(N__21363));
    Span4Mux_v I__2217 (
            .O(N__21368),
            .I(N__21360));
    Span4Mux_v I__2216 (
            .O(N__21363),
            .I(N__21357));
    Odrv4 I__2215 (
            .O(N__21360),
            .I(\pwm_generator_inst.N_17 ));
    Odrv4 I__2214 (
            .O(N__21357),
            .I(\pwm_generator_inst.N_17 ));
    InMux I__2213 (
            .O(N__21352),
            .I(N__21349));
    LocalMux I__2212 (
            .O(N__21349),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2 ));
    InMux I__2211 (
            .O(N__21346),
            .I(N__21343));
    LocalMux I__2210 (
            .O(N__21343),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_1 ));
    InMux I__2209 (
            .O(N__21340),
            .I(N__21337));
    LocalMux I__2208 (
            .O(N__21337),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_6 ));
    InMux I__2207 (
            .O(N__21334),
            .I(N__21331));
    LocalMux I__2206 (
            .O(N__21331),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_7 ));
    InMux I__2205 (
            .O(N__21328),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_6 ));
    CascadeMux I__2204 (
            .O(N__21325),
            .I(N__21322));
    InMux I__2203 (
            .O(N__21322),
            .I(N__21319));
    LocalMux I__2202 (
            .O(N__21319),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_8 ));
    InMux I__2201 (
            .O(N__21316),
            .I(bfn_3_9_0_));
    InMux I__2200 (
            .O(N__21313),
            .I(N__21310));
    LocalMux I__2199 (
            .O(N__21310),
            .I(N__21307));
    Odrv4 I__2198 (
            .O(N__21307),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO ));
    CascadeMux I__2197 (
            .O(N__21304),
            .I(N__21299));
    InMux I__2196 (
            .O(N__21303),
            .I(N__21287));
    InMux I__2195 (
            .O(N__21302),
            .I(N__21284));
    InMux I__2194 (
            .O(N__21299),
            .I(N__21281));
    InMux I__2193 (
            .O(N__21298),
            .I(N__21272));
    InMux I__2192 (
            .O(N__21297),
            .I(N__21272));
    InMux I__2191 (
            .O(N__21296),
            .I(N__21272));
    InMux I__2190 (
            .O(N__21295),
            .I(N__21272));
    InMux I__2189 (
            .O(N__21294),
            .I(N__21263));
    InMux I__2188 (
            .O(N__21293),
            .I(N__21263));
    InMux I__2187 (
            .O(N__21292),
            .I(N__21263));
    InMux I__2186 (
            .O(N__21291),
            .I(N__21263));
    InMux I__2185 (
            .O(N__21290),
            .I(N__21260));
    LocalMux I__2184 (
            .O(N__21287),
            .I(N__21253));
    LocalMux I__2183 (
            .O(N__21284),
            .I(N__21253));
    LocalMux I__2182 (
            .O(N__21281),
            .I(N__21253));
    LocalMux I__2181 (
            .O(N__21272),
            .I(N__21246));
    LocalMux I__2180 (
            .O(N__21263),
            .I(N__21246));
    LocalMux I__2179 (
            .O(N__21260),
            .I(N__21246));
    Span4Mux_v I__2178 (
            .O(N__21253),
            .I(N__21243));
    Span4Mux_v I__2177 (
            .O(N__21246),
            .I(N__21240));
    Odrv4 I__2176 (
            .O(N__21243),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    Odrv4 I__2175 (
            .O(N__21240),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    CascadeMux I__2174 (
            .O(N__21235),
            .I(N__21232));
    InMux I__2173 (
            .O(N__21232),
            .I(N__21229));
    LocalMux I__2172 (
            .O(N__21229),
            .I(N__21226));
    Span4Mux_h I__2171 (
            .O(N__21226),
            .I(N__21223));
    Odrv4 I__2170 (
            .O(N__21223),
            .I(\pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9 ));
    InMux I__2169 (
            .O(N__21220),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_8 ));
    CascadeMux I__2168 (
            .O(N__21217),
            .I(N__21214));
    InMux I__2167 (
            .O(N__21214),
            .I(N__21211));
    LocalMux I__2166 (
            .O(N__21211),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9 ));
    InMux I__2165 (
            .O(N__21208),
            .I(N__21205));
    LocalMux I__2164 (
            .O(N__21205),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8 ));
    InMux I__2163 (
            .O(N__21202),
            .I(N__21199));
    LocalMux I__2162 (
            .O(N__21199),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_8 ));
    InMux I__2161 (
            .O(N__21196),
            .I(N__21193));
    LocalMux I__2160 (
            .O(N__21193),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4 ));
    InMux I__2159 (
            .O(N__21190),
            .I(N__21187));
    LocalMux I__2158 (
            .O(N__21187),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_4 ));
    CascadeMux I__2157 (
            .O(N__21184),
            .I(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ));
    InMux I__2156 (
            .O(N__21181),
            .I(N__21174));
    InMux I__2155 (
            .O(N__21180),
            .I(N__21174));
    InMux I__2154 (
            .O(N__21179),
            .I(N__21171));
    LocalMux I__2153 (
            .O(N__21174),
            .I(N__21168));
    LocalMux I__2152 (
            .O(N__21171),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    Odrv4 I__2151 (
            .O(N__21168),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    InMux I__2150 (
            .O(N__21163),
            .I(N__21160));
    LocalMux I__2149 (
            .O(N__21160),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_0 ));
    InMux I__2148 (
            .O(N__21157),
            .I(N__21154));
    LocalMux I__2147 (
            .O(N__21154),
            .I(N__21151));
    Odrv4 I__2146 (
            .O(N__21151),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_1 ));
    InMux I__2145 (
            .O(N__21148),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_0 ));
    InMux I__2144 (
            .O(N__21145),
            .I(N__21142));
    LocalMux I__2143 (
            .O(N__21142),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_2 ));
    InMux I__2142 (
            .O(N__21139),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_1 ));
    InMux I__2141 (
            .O(N__21136),
            .I(N__21133));
    LocalMux I__2140 (
            .O(N__21133),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_3 ));
    InMux I__2139 (
            .O(N__21130),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_2 ));
    InMux I__2138 (
            .O(N__21127),
            .I(N__21124));
    LocalMux I__2137 (
            .O(N__21124),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_4 ));
    InMux I__2136 (
            .O(N__21121),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_3 ));
    InMux I__2135 (
            .O(N__21118),
            .I(N__21115));
    LocalMux I__2134 (
            .O(N__21115),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_5 ));
    InMux I__2133 (
            .O(N__21112),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_4 ));
    InMux I__2132 (
            .O(N__21109),
            .I(N__21106));
    LocalMux I__2131 (
            .O(N__21106),
            .I(N__21103));
    Odrv4 I__2130 (
            .O(N__21103),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_6 ));
    InMux I__2129 (
            .O(N__21100),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_5 ));
    InMux I__2128 (
            .O(N__21097),
            .I(N__21094));
    LocalMux I__2127 (
            .O(N__21094),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0 ));
    InMux I__2126 (
            .O(N__21091),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ));
    InMux I__2125 (
            .O(N__21088),
            .I(N__21085));
    LocalMux I__2124 (
            .O(N__21085),
            .I(N__21082));
    Span4Mux_v I__2123 (
            .O(N__21082),
            .I(N__21079));
    Odrv4 I__2122 (
            .O(N__21079),
            .I(\pwm_generator_inst.un2_threshold_acc_2_13 ));
    InMux I__2121 (
            .O(N__21076),
            .I(N__21073));
    LocalMux I__2120 (
            .O(N__21073),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0 ));
    InMux I__2119 (
            .O(N__21070),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ));
    CascadeMux I__2118 (
            .O(N__21067),
            .I(N__21064));
    InMux I__2117 (
            .O(N__21064),
            .I(N__21061));
    LocalMux I__2116 (
            .O(N__21061),
            .I(N__21058));
    Span4Mux_h I__2115 (
            .O(N__21058),
            .I(N__21055));
    Odrv4 I__2114 (
            .O(N__21055),
            .I(\pwm_generator_inst.un2_threshold_acc_2_14 ));
    InMux I__2113 (
            .O(N__21052),
            .I(N__21049));
    LocalMux I__2112 (
            .O(N__21049),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0 ));
    InMux I__2111 (
            .O(N__21046),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ));
    InMux I__2110 (
            .O(N__21043),
            .I(N__21040));
    LocalMux I__2109 (
            .O(N__21040),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0 ));
    InMux I__2108 (
            .O(N__21037),
            .I(N__21030));
    CascadeMux I__2107 (
            .O(N__21036),
            .I(N__21027));
    CascadeMux I__2106 (
            .O(N__21035),
            .I(N__21023));
    CascadeMux I__2105 (
            .O(N__21034),
            .I(N__21019));
    InMux I__2104 (
            .O(N__21033),
            .I(N__21015));
    LocalMux I__2103 (
            .O(N__21030),
            .I(N__21012));
    InMux I__2102 (
            .O(N__21027),
            .I(N__20999));
    InMux I__2101 (
            .O(N__21026),
            .I(N__20999));
    InMux I__2100 (
            .O(N__21023),
            .I(N__20999));
    InMux I__2099 (
            .O(N__21022),
            .I(N__20999));
    InMux I__2098 (
            .O(N__21019),
            .I(N__20999));
    InMux I__2097 (
            .O(N__21018),
            .I(N__20999));
    LocalMux I__2096 (
            .O(N__21015),
            .I(N__20992));
    Span4Mux_v I__2095 (
            .O(N__21012),
            .I(N__20992));
    LocalMux I__2094 (
            .O(N__20999),
            .I(N__20992));
    Span4Mux_v I__2093 (
            .O(N__20992),
            .I(N__20989));
    Odrv4 I__2092 (
            .O(N__20989),
            .I(\pwm_generator_inst.un2_threshold_acc_1_25 ));
    InMux I__2091 (
            .O(N__20986),
            .I(N__20983));
    LocalMux I__2090 (
            .O(N__20983),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0 ));
    InMux I__2089 (
            .O(N__20980),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ));
    InMux I__2088 (
            .O(N__20977),
            .I(N__20974));
    LocalMux I__2087 (
            .O(N__20974),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16 ));
    CascadeMux I__2086 (
            .O(N__20971),
            .I(N__20968));
    InMux I__2085 (
            .O(N__20968),
            .I(N__20965));
    LocalMux I__2084 (
            .O(N__20965),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO ));
    InMux I__2083 (
            .O(N__20962),
            .I(bfn_2_13_0_));
    InMux I__2082 (
            .O(N__20959),
            .I(N__20956));
    LocalMux I__2081 (
            .O(N__20956),
            .I(N__20953));
    Odrv4 I__2080 (
            .O(N__20953),
            .I(rgb_drv_RNOZ0));
    InMux I__2079 (
            .O(N__20950),
            .I(N__20947));
    LocalMux I__2078 (
            .O(N__20947),
            .I(N__20944));
    Odrv4 I__2077 (
            .O(N__20944),
            .I(\current_shift_inst.PI_CTRL.N_162 ));
    InMux I__2076 (
            .O(N__20941),
            .I(N__20938));
    LocalMux I__2075 (
            .O(N__20938),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ));
    InMux I__2074 (
            .O(N__20935),
            .I(N__20930));
    InMux I__2073 (
            .O(N__20934),
            .I(N__20927));
    InMux I__2072 (
            .O(N__20933),
            .I(N__20924));
    LocalMux I__2071 (
            .O(N__20930),
            .I(N__20919));
    LocalMux I__2070 (
            .O(N__20927),
            .I(N__20919));
    LocalMux I__2069 (
            .O(N__20924),
            .I(N__20916));
    Odrv4 I__2068 (
            .O(N__20919),
            .I(pwm_duty_input_3));
    Odrv4 I__2067 (
            .O(N__20916),
            .I(pwm_duty_input_3));
    CascadeMux I__2066 (
            .O(N__20911),
            .I(N__20908));
    InMux I__2065 (
            .O(N__20908),
            .I(N__20905));
    LocalMux I__2064 (
            .O(N__20905),
            .I(\pwm_generator_inst.un1_duty_inputlt3 ));
    InMux I__2063 (
            .O(N__20902),
            .I(N__20897));
    InMux I__2062 (
            .O(N__20901),
            .I(N__20894));
    InMux I__2061 (
            .O(N__20900),
            .I(N__20891));
    LocalMux I__2060 (
            .O(N__20897),
            .I(N__20888));
    LocalMux I__2059 (
            .O(N__20894),
            .I(N__20883));
    LocalMux I__2058 (
            .O(N__20891),
            .I(N__20883));
    Span4Mux_s1_h I__2057 (
            .O(N__20888),
            .I(N__20880));
    Odrv4 I__2056 (
            .O(N__20883),
            .I(pwm_duty_input_4));
    Odrv4 I__2055 (
            .O(N__20880),
            .I(pwm_duty_input_4));
    InMux I__2054 (
            .O(N__20875),
            .I(N__20872));
    LocalMux I__2053 (
            .O(N__20872),
            .I(N__20869));
    Span4Mux_v I__2052 (
            .O(N__20869),
            .I(N__20866));
    Odrv4 I__2051 (
            .O(N__20866),
            .I(\pwm_generator_inst.un2_threshold_acc_1_20 ));
    CascadeMux I__2050 (
            .O(N__20863),
            .I(N__20860));
    InMux I__2049 (
            .O(N__20860),
            .I(N__20857));
    LocalMux I__2048 (
            .O(N__20857),
            .I(N__20854));
    Span4Mux_v I__2047 (
            .O(N__20854),
            .I(N__20851));
    Odrv4 I__2046 (
            .O(N__20851),
            .I(\pwm_generator_inst.un2_threshold_acc_2_5 ));
    InMux I__2045 (
            .O(N__20848),
            .I(N__20845));
    LocalMux I__2044 (
            .O(N__20845),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0 ));
    InMux I__2043 (
            .O(N__20842),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ));
    InMux I__2042 (
            .O(N__20839),
            .I(N__20836));
    LocalMux I__2041 (
            .O(N__20836),
            .I(N__20833));
    Span4Mux_v I__2040 (
            .O(N__20833),
            .I(N__20830));
    Odrv4 I__2039 (
            .O(N__20830),
            .I(\pwm_generator_inst.un2_threshold_acc_1_21 ));
    CascadeMux I__2038 (
            .O(N__20827),
            .I(N__20824));
    InMux I__2037 (
            .O(N__20824),
            .I(N__20821));
    LocalMux I__2036 (
            .O(N__20821),
            .I(N__20818));
    Span4Mux_h I__2035 (
            .O(N__20818),
            .I(N__20815));
    Odrv4 I__2034 (
            .O(N__20815),
            .I(\pwm_generator_inst.un2_threshold_acc_2_6 ));
    InMux I__2033 (
            .O(N__20812),
            .I(N__20809));
    LocalMux I__2032 (
            .O(N__20809),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0 ));
    InMux I__2031 (
            .O(N__20806),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ));
    InMux I__2030 (
            .O(N__20803),
            .I(N__20800));
    LocalMux I__2029 (
            .O(N__20800),
            .I(N__20797));
    Span4Mux_v I__2028 (
            .O(N__20797),
            .I(N__20794));
    Odrv4 I__2027 (
            .O(N__20794),
            .I(\pwm_generator_inst.un2_threshold_acc_1_22 ));
    CascadeMux I__2026 (
            .O(N__20791),
            .I(N__20788));
    InMux I__2025 (
            .O(N__20788),
            .I(N__20785));
    LocalMux I__2024 (
            .O(N__20785),
            .I(N__20782));
    Span4Mux_h I__2023 (
            .O(N__20782),
            .I(N__20779));
    Odrv4 I__2022 (
            .O(N__20779),
            .I(\pwm_generator_inst.un2_threshold_acc_2_7 ));
    InMux I__2021 (
            .O(N__20776),
            .I(N__20773));
    LocalMux I__2020 (
            .O(N__20773),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0 ));
    InMux I__2019 (
            .O(N__20770),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ));
    InMux I__2018 (
            .O(N__20767),
            .I(N__20764));
    LocalMux I__2017 (
            .O(N__20764),
            .I(N__20761));
    Span4Mux_h I__2016 (
            .O(N__20761),
            .I(N__20758));
    Span4Mux_v I__2015 (
            .O(N__20758),
            .I(N__20755));
    Odrv4 I__2014 (
            .O(N__20755),
            .I(\pwm_generator_inst.un2_threshold_acc_1_23 ));
    CascadeMux I__2013 (
            .O(N__20752),
            .I(N__20749));
    InMux I__2012 (
            .O(N__20749),
            .I(N__20746));
    LocalMux I__2011 (
            .O(N__20746),
            .I(N__20743));
    Span4Mux_h I__2010 (
            .O(N__20743),
            .I(N__20740));
    Odrv4 I__2009 (
            .O(N__20740),
            .I(\pwm_generator_inst.un2_threshold_acc_2_8 ));
    InMux I__2008 (
            .O(N__20737),
            .I(N__20734));
    LocalMux I__2007 (
            .O(N__20734),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0 ));
    InMux I__2006 (
            .O(N__20731),
            .I(bfn_2_12_0_));
    InMux I__2005 (
            .O(N__20728),
            .I(N__20725));
    LocalMux I__2004 (
            .O(N__20725),
            .I(N__20722));
    Span4Mux_v I__2003 (
            .O(N__20722),
            .I(N__20719));
    Odrv4 I__2002 (
            .O(N__20719),
            .I(\pwm_generator_inst.un2_threshold_acc_1_24 ));
    CascadeMux I__2001 (
            .O(N__20716),
            .I(N__20713));
    InMux I__2000 (
            .O(N__20713),
            .I(N__20710));
    LocalMux I__1999 (
            .O(N__20710),
            .I(N__20707));
    Span4Mux_h I__1998 (
            .O(N__20707),
            .I(N__20704));
    Odrv4 I__1997 (
            .O(N__20704),
            .I(\pwm_generator_inst.un2_threshold_acc_2_9 ));
    InMux I__1996 (
            .O(N__20701),
            .I(N__20698));
    LocalMux I__1995 (
            .O(N__20698),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0 ));
    InMux I__1994 (
            .O(N__20695),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ));
    CascadeMux I__1993 (
            .O(N__20692),
            .I(N__20689));
    InMux I__1992 (
            .O(N__20689),
            .I(N__20686));
    LocalMux I__1991 (
            .O(N__20686),
            .I(N__20683));
    Span4Mux_h I__1990 (
            .O(N__20683),
            .I(N__20680));
    Odrv4 I__1989 (
            .O(N__20680),
            .I(\pwm_generator_inst.un2_threshold_acc_2_10 ));
    InMux I__1988 (
            .O(N__20677),
            .I(N__20674));
    LocalMux I__1987 (
            .O(N__20674),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0 ));
    InMux I__1986 (
            .O(N__20671),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ));
    InMux I__1985 (
            .O(N__20668),
            .I(N__20665));
    LocalMux I__1984 (
            .O(N__20665),
            .I(N__20662));
    Span4Mux_h I__1983 (
            .O(N__20662),
            .I(N__20659));
    Odrv4 I__1982 (
            .O(N__20659),
            .I(\pwm_generator_inst.un2_threshold_acc_2_11 ));
    InMux I__1981 (
            .O(N__20656),
            .I(N__20653));
    LocalMux I__1980 (
            .O(N__20653),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0 ));
    InMux I__1979 (
            .O(N__20650),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ));
    CascadeMux I__1978 (
            .O(N__20647),
            .I(N__20644));
    InMux I__1977 (
            .O(N__20644),
            .I(N__20641));
    LocalMux I__1976 (
            .O(N__20641),
            .I(N__20638));
    Span4Mux_v I__1975 (
            .O(N__20638),
            .I(N__20635));
    Odrv4 I__1974 (
            .O(N__20635),
            .I(\pwm_generator_inst.un2_threshold_acc_2_12 ));
    InMux I__1973 (
            .O(N__20632),
            .I(N__20628));
    InMux I__1972 (
            .O(N__20631),
            .I(N__20625));
    LocalMux I__1971 (
            .O(N__20628),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ));
    LocalMux I__1970 (
            .O(N__20625),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ));
    InMux I__1969 (
            .O(N__20620),
            .I(N__20614));
    InMux I__1968 (
            .O(N__20619),
            .I(N__20614));
    LocalMux I__1967 (
            .O(N__20614),
            .I(N__20611));
    Span4Mux_h I__1966 (
            .O(N__20611),
            .I(N__20608));
    Odrv4 I__1965 (
            .O(N__20608),
            .I(\pwm_generator_inst.O_10 ));
    InMux I__1964 (
            .O(N__20605),
            .I(N__20602));
    LocalMux I__1963 (
            .O(N__20602),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO ));
    CascadeMux I__1962 (
            .O(N__20599),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_10_cascade_ ));
    InMux I__1961 (
            .O(N__20596),
            .I(N__20593));
    LocalMux I__1960 (
            .O(N__20593),
            .I(N__20589));
    InMux I__1959 (
            .O(N__20592),
            .I(N__20586));
    Odrv4 I__1958 (
            .O(N__20589),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ));
    LocalMux I__1957 (
            .O(N__20586),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ));
    InMux I__1956 (
            .O(N__20581),
            .I(N__20577));
    InMux I__1955 (
            .O(N__20580),
            .I(N__20573));
    LocalMux I__1954 (
            .O(N__20577),
            .I(N__20570));
    InMux I__1953 (
            .O(N__20576),
            .I(N__20567));
    LocalMux I__1952 (
            .O(N__20573),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ));
    Odrv4 I__1951 (
            .O(N__20570),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ));
    LocalMux I__1950 (
            .O(N__20567),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ));
    InMux I__1949 (
            .O(N__20560),
            .I(N__20557));
    LocalMux I__1948 (
            .O(N__20557),
            .I(N__20554));
    Span4Mux_h I__1947 (
            .O(N__20554),
            .I(N__20551));
    Odrv4 I__1946 (
            .O(N__20551),
            .I(\pwm_generator_inst.un2_threshold_acc_2_0 ));
    CascadeMux I__1945 (
            .O(N__20548),
            .I(N__20545));
    InMux I__1944 (
            .O(N__20545),
            .I(N__20542));
    LocalMux I__1943 (
            .O(N__20542),
            .I(N__20539));
    Span4Mux_h I__1942 (
            .O(N__20539),
            .I(N__20536));
    Span4Mux_v I__1941 (
            .O(N__20536),
            .I(N__20533));
    Odrv4 I__1940 (
            .O(N__20533),
            .I(\pwm_generator_inst.un2_threshold_acc_1_15 ));
    InMux I__1939 (
            .O(N__20530),
            .I(N__20527));
    LocalMux I__1938 (
            .O(N__20527),
            .I(\pwm_generator_inst.un3_threshold_acc_axbZ0Z_4 ));
    InMux I__1937 (
            .O(N__20524),
            .I(N__20521));
    LocalMux I__1936 (
            .O(N__20521),
            .I(N__20518));
    Span4Mux_v I__1935 (
            .O(N__20518),
            .I(N__20515));
    Odrv4 I__1934 (
            .O(N__20515),
            .I(\pwm_generator_inst.un2_threshold_acc_1_16 ));
    CascadeMux I__1933 (
            .O(N__20512),
            .I(N__20509));
    InMux I__1932 (
            .O(N__20509),
            .I(N__20506));
    LocalMux I__1931 (
            .O(N__20506),
            .I(N__20503));
    Span4Mux_h I__1930 (
            .O(N__20503),
            .I(N__20500));
    Odrv4 I__1929 (
            .O(N__20500),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1 ));
    CascadeMux I__1928 (
            .O(N__20497),
            .I(N__20494));
    InMux I__1927 (
            .O(N__20494),
            .I(N__20491));
    LocalMux I__1926 (
            .O(N__20491),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0 ));
    InMux I__1925 (
            .O(N__20488),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ));
    InMux I__1924 (
            .O(N__20485),
            .I(N__20482));
    LocalMux I__1923 (
            .O(N__20482),
            .I(N__20479));
    Span4Mux_v I__1922 (
            .O(N__20479),
            .I(N__20476));
    Odrv4 I__1921 (
            .O(N__20476),
            .I(\pwm_generator_inst.un2_threshold_acc_1_17 ));
    CascadeMux I__1920 (
            .O(N__20473),
            .I(N__20470));
    InMux I__1919 (
            .O(N__20470),
            .I(N__20467));
    LocalMux I__1918 (
            .O(N__20467),
            .I(N__20464));
    Span4Mux_h I__1917 (
            .O(N__20464),
            .I(N__20461));
    Odrv4 I__1916 (
            .O(N__20461),
            .I(\pwm_generator_inst.un2_threshold_acc_2_2 ));
    InMux I__1915 (
            .O(N__20458),
            .I(N__20455));
    LocalMux I__1914 (
            .O(N__20455),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0 ));
    InMux I__1913 (
            .O(N__20452),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ));
    InMux I__1912 (
            .O(N__20449),
            .I(N__20446));
    LocalMux I__1911 (
            .O(N__20446),
            .I(N__20443));
    Span4Mux_s3_h I__1910 (
            .O(N__20443),
            .I(N__20440));
    Span4Mux_v I__1909 (
            .O(N__20440),
            .I(N__20437));
    Odrv4 I__1908 (
            .O(N__20437),
            .I(\pwm_generator_inst.un2_threshold_acc_1_18 ));
    CascadeMux I__1907 (
            .O(N__20434),
            .I(N__20431));
    InMux I__1906 (
            .O(N__20431),
            .I(N__20428));
    LocalMux I__1905 (
            .O(N__20428),
            .I(N__20425));
    Span4Mux_h I__1904 (
            .O(N__20425),
            .I(N__20422));
    Odrv4 I__1903 (
            .O(N__20422),
            .I(\pwm_generator_inst.un2_threshold_acc_2_3 ));
    InMux I__1902 (
            .O(N__20419),
            .I(N__20416));
    LocalMux I__1901 (
            .O(N__20416),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0 ));
    InMux I__1900 (
            .O(N__20413),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ));
    InMux I__1899 (
            .O(N__20410),
            .I(N__20407));
    LocalMux I__1898 (
            .O(N__20407),
            .I(N__20404));
    Span4Mux_v I__1897 (
            .O(N__20404),
            .I(N__20401));
    Odrv4 I__1896 (
            .O(N__20401),
            .I(\pwm_generator_inst.un2_threshold_acc_1_19 ));
    CascadeMux I__1895 (
            .O(N__20398),
            .I(N__20395));
    InMux I__1894 (
            .O(N__20395),
            .I(N__20392));
    LocalMux I__1893 (
            .O(N__20392),
            .I(N__20389));
    Span4Mux_v I__1892 (
            .O(N__20389),
            .I(N__20386));
    Odrv4 I__1891 (
            .O(N__20386),
            .I(\pwm_generator_inst.un2_threshold_acc_2_4 ));
    InMux I__1890 (
            .O(N__20383),
            .I(N__20380));
    LocalMux I__1889 (
            .O(N__20380),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0 ));
    InMux I__1888 (
            .O(N__20377),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ));
    InMux I__1887 (
            .O(N__20374),
            .I(N__20370));
    InMux I__1886 (
            .O(N__20373),
            .I(N__20367));
    LocalMux I__1885 (
            .O(N__20370),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ));
    LocalMux I__1884 (
            .O(N__20367),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ));
    InMux I__1883 (
            .O(N__20362),
            .I(N__20359));
    LocalMux I__1882 (
            .O(N__20359),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO ));
    CascadeMux I__1881 (
            .O(N__20356),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_14_cascade_ ));
    InMux I__1880 (
            .O(N__20353),
            .I(N__20349));
    InMux I__1879 (
            .O(N__20352),
            .I(N__20346));
    LocalMux I__1878 (
            .O(N__20349),
            .I(N__20341));
    LocalMux I__1877 (
            .O(N__20346),
            .I(N__20341));
    Odrv4 I__1876 (
            .O(N__20341),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ));
    InMux I__1875 (
            .O(N__20338),
            .I(N__20333));
    InMux I__1874 (
            .O(N__20337),
            .I(N__20330));
    InMux I__1873 (
            .O(N__20336),
            .I(N__20327));
    LocalMux I__1872 (
            .O(N__20333),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ));
    LocalMux I__1871 (
            .O(N__20330),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ));
    LocalMux I__1870 (
            .O(N__20327),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ));
    CascadeMux I__1869 (
            .O(N__20320),
            .I(N__20317));
    InMux I__1868 (
            .O(N__20317),
            .I(N__20314));
    LocalMux I__1867 (
            .O(N__20314),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO ));
    InMux I__1866 (
            .O(N__20311),
            .I(N__20308));
    LocalMux I__1865 (
            .O(N__20308),
            .I(N__20304));
    InMux I__1864 (
            .O(N__20307),
            .I(N__20301));
    Odrv4 I__1863 (
            .O(N__20304),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ));
    LocalMux I__1862 (
            .O(N__20301),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ));
    InMux I__1861 (
            .O(N__20296),
            .I(N__20293));
    LocalMux I__1860 (
            .O(N__20293),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO ));
    InMux I__1859 (
            .O(N__20290),
            .I(N__20285));
    InMux I__1858 (
            .O(N__20289),
            .I(N__20280));
    InMux I__1857 (
            .O(N__20288),
            .I(N__20280));
    LocalMux I__1856 (
            .O(N__20285),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ));
    LocalMux I__1855 (
            .O(N__20280),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ));
    CascadeMux I__1854 (
            .O(N__20275),
            .I(N__20272));
    InMux I__1853 (
            .O(N__20272),
            .I(N__20268));
    InMux I__1852 (
            .O(N__20271),
            .I(N__20265));
    LocalMux I__1851 (
            .O(N__20268),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ));
    LocalMux I__1850 (
            .O(N__20265),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ));
    InMux I__1849 (
            .O(N__20260),
            .I(N__20256));
    InMux I__1848 (
            .O(N__20259),
            .I(N__20253));
    LocalMux I__1847 (
            .O(N__20256),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ));
    LocalMux I__1846 (
            .O(N__20253),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ));
    InMux I__1845 (
            .O(N__20248),
            .I(N__20242));
    InMux I__1844 (
            .O(N__20247),
            .I(N__20242));
    LocalMux I__1843 (
            .O(N__20242),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ));
    InMux I__1842 (
            .O(N__20239),
            .I(N__20236));
    LocalMux I__1841 (
            .O(N__20236),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO ));
    CascadeMux I__1840 (
            .O(N__20233),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_ ));
    InMux I__1839 (
            .O(N__20230),
            .I(N__20226));
    InMux I__1838 (
            .O(N__20229),
            .I(N__20223));
    LocalMux I__1837 (
            .O(N__20226),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ));
    LocalMux I__1836 (
            .O(N__20223),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ));
    InMux I__1835 (
            .O(N__20218),
            .I(N__20212));
    InMux I__1834 (
            .O(N__20217),
            .I(N__20212));
    LocalMux I__1833 (
            .O(N__20212),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ));
    InMux I__1832 (
            .O(N__20209),
            .I(N__20206));
    LocalMux I__1831 (
            .O(N__20206),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO ));
    CascadeMux I__1830 (
            .O(N__20203),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_18_cascade_ ));
    InMux I__1829 (
            .O(N__20200),
            .I(N__20197));
    LocalMux I__1828 (
            .O(N__20197),
            .I(\current_shift_inst.PI_CTRL.N_164 ));
    CascadeMux I__1827 (
            .O(N__20194),
            .I(\current_shift_inst.PI_CTRL.N_164_cascade_ ));
    InMux I__1826 (
            .O(N__20191),
            .I(N__20182));
    InMux I__1825 (
            .O(N__20190),
            .I(N__20182));
    InMux I__1824 (
            .O(N__20189),
            .I(N__20182));
    LocalMux I__1823 (
            .O(N__20182),
            .I(\current_shift_inst.PI_CTRL.N_120 ));
    InMux I__1822 (
            .O(N__20179),
            .I(N__20176));
    LocalMux I__1821 (
            .O(N__20176),
            .I(\current_shift_inst.PI_CTRL.N_167 ));
    CascadeMux I__1820 (
            .O(N__20173),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_ ));
    CascadeMux I__1819 (
            .O(N__20170),
            .I(N__20167));
    InMux I__1818 (
            .O(N__20167),
            .I(N__20164));
    LocalMux I__1817 (
            .O(N__20164),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    InMux I__1816 (
            .O(N__20161),
            .I(N__20158));
    LocalMux I__1815 (
            .O(N__20158),
            .I(\current_shift_inst.PI_CTRL.N_168 ));
    CascadeMux I__1814 (
            .O(N__20155),
            .I(\current_shift_inst.PI_CTRL.N_27_cascade_ ));
    InMux I__1813 (
            .O(N__20152),
            .I(N__20148));
    InMux I__1812 (
            .O(N__20151),
            .I(N__20145));
    LocalMux I__1811 (
            .O(N__20148),
            .I(\current_shift_inst.PI_CTRL.N_166 ));
    LocalMux I__1810 (
            .O(N__20145),
            .I(\current_shift_inst.PI_CTRL.N_166 ));
    InMux I__1809 (
            .O(N__20140),
            .I(N__20135));
    InMux I__1808 (
            .O(N__20139),
            .I(N__20132));
    InMux I__1807 (
            .O(N__20138),
            .I(N__20129));
    LocalMux I__1806 (
            .O(N__20135),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ));
    LocalMux I__1805 (
            .O(N__20132),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ));
    LocalMux I__1804 (
            .O(N__20129),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ));
    CascadeMux I__1803 (
            .O(N__20122),
            .I(N__20119));
    InMux I__1802 (
            .O(N__20119),
            .I(N__20116));
    LocalMux I__1801 (
            .O(N__20116),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO ));
    InMux I__1800 (
            .O(N__20113),
            .I(N__20110));
    LocalMux I__1799 (
            .O(N__20110),
            .I(N__20107));
    Span4Mux_h I__1798 (
            .O(N__20107),
            .I(N__20103));
    InMux I__1797 (
            .O(N__20106),
            .I(N__20100));
    Odrv4 I__1796 (
            .O(N__20103),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ));
    LocalMux I__1795 (
            .O(N__20100),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ));
    CascadeMux I__1794 (
            .O(N__20095),
            .I(N__20092));
    InMux I__1793 (
            .O(N__20092),
            .I(N__20089));
    LocalMux I__1792 (
            .O(N__20089),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO ));
    InMux I__1791 (
            .O(N__20086),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_19 ));
    InMux I__1790 (
            .O(N__20083),
            .I(N__20080));
    LocalMux I__1789 (
            .O(N__20080),
            .I(N__20076));
    InMux I__1788 (
            .O(N__20079),
            .I(N__20073));
    Odrv4 I__1787 (
            .O(N__20076),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1_15 ));
    LocalMux I__1786 (
            .O(N__20073),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1_15 ));
    CascadeMux I__1785 (
            .O(N__20068),
            .I(N__20065));
    InMux I__1784 (
            .O(N__20065),
            .I(N__20062));
    LocalMux I__1783 (
            .O(N__20062),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1_16 ));
    InMux I__1782 (
            .O(N__20059),
            .I(N__20056));
    LocalMux I__1781 (
            .O(N__20056),
            .I(N_34_i_i));
    CascadeMux I__1780 (
            .O(N__20053),
            .I(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_ ));
    InMux I__1779 (
            .O(N__20050),
            .I(N__20046));
    InMux I__1778 (
            .O(N__20049),
            .I(N__20043));
    LocalMux I__1777 (
            .O(N__20046),
            .I(N__20040));
    LocalMux I__1776 (
            .O(N__20043),
            .I(pwm_duty_input_0));
    Odrv4 I__1775 (
            .O(N__20040),
            .I(pwm_duty_input_0));
    InMux I__1774 (
            .O(N__20035),
            .I(N__20031));
    InMux I__1773 (
            .O(N__20034),
            .I(N__20028));
    LocalMux I__1772 (
            .O(N__20031),
            .I(N__20025));
    LocalMux I__1771 (
            .O(N__20028),
            .I(pwm_duty_input_1));
    Odrv4 I__1770 (
            .O(N__20025),
            .I(pwm_duty_input_1));
    InMux I__1769 (
            .O(N__20020),
            .I(N__20016));
    InMux I__1768 (
            .O(N__20019),
            .I(N__20013));
    LocalMux I__1767 (
            .O(N__20016),
            .I(N__20010));
    LocalMux I__1766 (
            .O(N__20013),
            .I(pwm_duty_input_2));
    Odrv4 I__1765 (
            .O(N__20010),
            .I(pwm_duty_input_2));
    CascadeMux I__1764 (
            .O(N__20005),
            .I(N__20002));
    InMux I__1763 (
            .O(N__20002),
            .I(N__19995));
    InMux I__1762 (
            .O(N__20001),
            .I(N__19995));
    InMux I__1761 (
            .O(N__20000),
            .I(N__19992));
    LocalMux I__1760 (
            .O(N__19995),
            .I(pwm_duty_input_7));
    LocalMux I__1759 (
            .O(N__19992),
            .I(pwm_duty_input_7));
    InMux I__1758 (
            .O(N__19987),
            .I(N__19984));
    LocalMux I__1757 (
            .O(N__19984),
            .I(N__19979));
    InMux I__1756 (
            .O(N__19983),
            .I(N__19974));
    InMux I__1755 (
            .O(N__19982),
            .I(N__19974));
    Span4Mux_v I__1754 (
            .O(N__19979),
            .I(N__19971));
    LocalMux I__1753 (
            .O(N__19974),
            .I(pwm_duty_input_5));
    Odrv4 I__1752 (
            .O(N__19971),
            .I(pwm_duty_input_5));
    InMux I__1751 (
            .O(N__19966),
            .I(N__19961));
    InMux I__1750 (
            .O(N__19965),
            .I(N__19958));
    InMux I__1749 (
            .O(N__19964),
            .I(N__19955));
    LocalMux I__1748 (
            .O(N__19961),
            .I(N__19952));
    LocalMux I__1747 (
            .O(N__19958),
            .I(pwm_duty_input_8));
    LocalMux I__1746 (
            .O(N__19955),
            .I(pwm_duty_input_8));
    Odrv4 I__1745 (
            .O(N__19952),
            .I(pwm_duty_input_8));
    InMux I__1744 (
            .O(N__19945),
            .I(N__19938));
    InMux I__1743 (
            .O(N__19944),
            .I(N__19938));
    InMux I__1742 (
            .O(N__19943),
            .I(N__19935));
    LocalMux I__1741 (
            .O(N__19938),
            .I(pwm_duty_input_9));
    LocalMux I__1740 (
            .O(N__19935),
            .I(pwm_duty_input_9));
    CascadeMux I__1739 (
            .O(N__19930),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ));
    InMux I__1738 (
            .O(N__19927),
            .I(N__19920));
    InMux I__1737 (
            .O(N__19926),
            .I(N__19920));
    InMux I__1736 (
            .O(N__19925),
            .I(N__19917));
    LocalMux I__1735 (
            .O(N__19920),
            .I(pwm_duty_input_6));
    LocalMux I__1734 (
            .O(N__19917),
            .I(pwm_duty_input_6));
    InMux I__1733 (
            .O(N__19912),
            .I(N__19909));
    LocalMux I__1732 (
            .O(N__19909),
            .I(N__19906));
    Span4Mux_v I__1731 (
            .O(N__19906),
            .I(N__19903));
    Odrv4 I__1730 (
            .O(N__19903),
            .I(\pwm_generator_inst.O_13 ));
    InMux I__1729 (
            .O(N__19900),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_1 ));
    InMux I__1728 (
            .O(N__19897),
            .I(N__19894));
    LocalMux I__1727 (
            .O(N__19894),
            .I(N__19891));
    Span4Mux_v I__1726 (
            .O(N__19891),
            .I(N__19888));
    Odrv4 I__1725 (
            .O(N__19888),
            .I(\pwm_generator_inst.O_14 ));
    InMux I__1724 (
            .O(N__19885),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_2 ));
    InMux I__1723 (
            .O(N__19882),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_3 ));
    InMux I__1722 (
            .O(N__19879),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_4 ));
    InMux I__1721 (
            .O(N__19876),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_5 ));
    InMux I__1720 (
            .O(N__19873),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_6 ));
    InMux I__1719 (
            .O(N__19870),
            .I(bfn_1_11_0_));
    InMux I__1718 (
            .O(N__19867),
            .I(bfn_1_9_0_));
    InMux I__1717 (
            .O(N__19864),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_16 ));
    InMux I__1716 (
            .O(N__19861),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_17 ));
    InMux I__1715 (
            .O(N__19858),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_18 ));
    InMux I__1714 (
            .O(N__19855),
            .I(N__19851));
    InMux I__1713 (
            .O(N__19854),
            .I(N__19848));
    LocalMux I__1712 (
            .O(N__19851),
            .I(N__19843));
    LocalMux I__1711 (
            .O(N__19848),
            .I(N__19843));
    Span4Mux_v I__1710 (
            .O(N__19843),
            .I(N__19840));
    Odrv4 I__1709 (
            .O(N__19840),
            .I(\pwm_generator_inst.un3_threshold_acc ));
    InMux I__1708 (
            .O(N__19837),
            .I(N__19834));
    LocalMux I__1707 (
            .O(N__19834),
            .I(N__19831));
    Span4Mux_v I__1706 (
            .O(N__19831),
            .I(N__19828));
    Odrv4 I__1705 (
            .O(N__19828),
            .I(\pwm_generator_inst.O_12 ));
    InMux I__1704 (
            .O(N__19825),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_0 ));
    InMux I__1703 (
            .O(N__19822),
            .I(N__19819));
    LocalMux I__1702 (
            .O(N__19819),
            .I(N__19816));
    Span4Mux_h I__1701 (
            .O(N__19816),
            .I(N__19813));
    Odrv4 I__1700 (
            .O(N__19813),
            .I(\pwm_generator_inst.O_8 ));
    InMux I__1699 (
            .O(N__19810),
            .I(N__19807));
    LocalMux I__1698 (
            .O(N__19807),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_8 ));
    InMux I__1697 (
            .O(N__19804),
            .I(N__19801));
    LocalMux I__1696 (
            .O(N__19801),
            .I(N__19798));
    Odrv4 I__1695 (
            .O(N__19798),
            .I(\pwm_generator_inst.O_9 ));
    InMux I__1694 (
            .O(N__19795),
            .I(N__19792));
    LocalMux I__1693 (
            .O(N__19792),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_9 ));
    InMux I__1692 (
            .O(N__19789),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_9 ));
    InMux I__1691 (
            .O(N__19786),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_10 ));
    InMux I__1690 (
            .O(N__19783),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_11 ));
    InMux I__1689 (
            .O(N__19780),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_12 ));
    InMux I__1688 (
            .O(N__19777),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_13 ));
    InMux I__1687 (
            .O(N__19774),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_14 ));
    InMux I__1686 (
            .O(N__19771),
            .I(N__19768));
    LocalMux I__1685 (
            .O(N__19768),
            .I(N__19765));
    Span4Mux_h I__1684 (
            .O(N__19765),
            .I(N__19762));
    Odrv4 I__1683 (
            .O(N__19762),
            .I(\pwm_generator_inst.O_0 ));
    InMux I__1682 (
            .O(N__19759),
            .I(N__19756));
    LocalMux I__1681 (
            .O(N__19756),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_0 ));
    InMux I__1680 (
            .O(N__19753),
            .I(N__19750));
    LocalMux I__1679 (
            .O(N__19750),
            .I(N__19747));
    Span4Mux_v I__1678 (
            .O(N__19747),
            .I(N__19744));
    Odrv4 I__1677 (
            .O(N__19744),
            .I(\pwm_generator_inst.O_1 ));
    InMux I__1676 (
            .O(N__19741),
            .I(N__19738));
    LocalMux I__1675 (
            .O(N__19738),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_1 ));
    InMux I__1674 (
            .O(N__19735),
            .I(N__19732));
    LocalMux I__1673 (
            .O(N__19732),
            .I(N__19729));
    Odrv4 I__1672 (
            .O(N__19729),
            .I(\pwm_generator_inst.O_2 ));
    InMux I__1671 (
            .O(N__19726),
            .I(N__19723));
    LocalMux I__1670 (
            .O(N__19723),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_2 ));
    InMux I__1669 (
            .O(N__19720),
            .I(N__19717));
    LocalMux I__1668 (
            .O(N__19717),
            .I(N__19714));
    Odrv4 I__1667 (
            .O(N__19714),
            .I(\pwm_generator_inst.O_3 ));
    InMux I__1666 (
            .O(N__19711),
            .I(N__19708));
    LocalMux I__1665 (
            .O(N__19708),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_3 ));
    InMux I__1664 (
            .O(N__19705),
            .I(N__19702));
    LocalMux I__1663 (
            .O(N__19702),
            .I(N__19699));
    Odrv4 I__1662 (
            .O(N__19699),
            .I(\pwm_generator_inst.O_4 ));
    InMux I__1661 (
            .O(N__19696),
            .I(N__19693));
    LocalMux I__1660 (
            .O(N__19693),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_4 ));
    InMux I__1659 (
            .O(N__19690),
            .I(N__19687));
    LocalMux I__1658 (
            .O(N__19687),
            .I(N__19684));
    Odrv4 I__1657 (
            .O(N__19684),
            .I(\pwm_generator_inst.O_5 ));
    InMux I__1656 (
            .O(N__19681),
            .I(N__19678));
    LocalMux I__1655 (
            .O(N__19678),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_5 ));
    InMux I__1654 (
            .O(N__19675),
            .I(N__19672));
    LocalMux I__1653 (
            .O(N__19672),
            .I(N__19669));
    Span4Mux_h I__1652 (
            .O(N__19669),
            .I(N__19666));
    Odrv4 I__1651 (
            .O(N__19666),
            .I(\pwm_generator_inst.O_6 ));
    InMux I__1650 (
            .O(N__19663),
            .I(N__19660));
    LocalMux I__1649 (
            .O(N__19660),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_6 ));
    InMux I__1648 (
            .O(N__19657),
            .I(N__19654));
    LocalMux I__1647 (
            .O(N__19654),
            .I(N__19651));
    Span4Mux_v I__1646 (
            .O(N__19651),
            .I(N__19648));
    Odrv4 I__1645 (
            .O(N__19648),
            .I(\pwm_generator_inst.O_7 ));
    InMux I__1644 (
            .O(N__19645),
            .I(N__19642));
    LocalMux I__1643 (
            .O(N__19642),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_7 ));
    defparam IN_MUX_bfv_16_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_8_0_));
    defparam IN_MUX_bfv_16_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_9_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un13_integrator_cry_6 ),
            .carryinitout(bfn_16_9_0_));
    defparam IN_MUX_bfv_16_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_10_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un13_integrator_cry_14 ),
            .carryinitout(bfn_16_10_0_));
    defparam IN_MUX_bfv_16_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_11_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un13_integrator_cry_22 ),
            .carryinitout(bfn_16_11_0_));
    defparam IN_MUX_bfv_16_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_12_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un13_integrator_cry_30 ),
            .carryinitout(bfn_16_12_0_));
    defparam IN_MUX_bfv_1_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_10_0_));
    defparam IN_MUX_bfv_1_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_11_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_acc_cry_7 ),
            .carryinitout(bfn_1_11_0_));
    defparam IN_MUX_bfv_1_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_12_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_acc_cry_15 ),
            .carryinitout(bfn_1_12_0_));
    defparam IN_MUX_bfv_7_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_15_0_));
    defparam IN_MUX_bfv_7_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_16_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_7_16_0_));
    defparam IN_MUX_bfv_7_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_17_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_7_17_0_));
    defparam IN_MUX_bfv_10_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_17_0_));
    defparam IN_MUX_bfv_10_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_18_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_10_18_0_));
    defparam IN_MUX_bfv_10_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_19_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_10_19_0_));
    defparam IN_MUX_bfv_11_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_18_0_));
    defparam IN_MUX_bfv_11_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_19_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_11_19_0_));
    defparam IN_MUX_bfv_11_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_20_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_11_20_0_));
    defparam IN_MUX_bfv_8_20_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_20_0_));
    defparam IN_MUX_bfv_8_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_21_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_8_21_0_));
    defparam IN_MUX_bfv_8_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_22_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_8_22_0_));
    defparam IN_MUX_bfv_9_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_22_0_));
    defparam IN_MUX_bfv_9_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_23_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_9_23_0_));
    defparam IN_MUX_bfv_9_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_24_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_9_24_0_));
    defparam IN_MUX_bfv_10_24_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_24_0_));
    defparam IN_MUX_bfv_10_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_25_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_10_25_0_));
    defparam IN_MUX_bfv_10_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_26_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_10_26_0_));
    defparam IN_MUX_bfv_15_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_19_0_));
    defparam IN_MUX_bfv_15_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_20_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .carryinitout(bfn_15_20_0_));
    defparam IN_MUX_bfv_15_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_21_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .carryinitout(bfn_15_21_0_));
    defparam IN_MUX_bfv_15_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_22_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .carryinitout(bfn_15_22_0_));
    defparam IN_MUX_bfv_13_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_17_0_));
    defparam IN_MUX_bfv_13_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_18_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .carryinitout(bfn_13_18_0_));
    defparam IN_MUX_bfv_13_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_19_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .carryinitout(bfn_13_19_0_));
    defparam IN_MUX_bfv_13_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_20_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .carryinitout(bfn_13_20_0_));
    defparam IN_MUX_bfv_15_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_15_0_));
    defparam IN_MUX_bfv_15_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_16_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_7 ),
            .carryinitout(bfn_15_16_0_));
    defparam IN_MUX_bfv_15_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_17_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_15 ),
            .carryinitout(bfn_15_17_0_));
    defparam IN_MUX_bfv_15_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_18_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_23 ),
            .carryinitout(bfn_15_18_0_));
    defparam IN_MUX_bfv_2_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_11_0_));
    defparam IN_MUX_bfv_2_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_12_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7 ),
            .carryinitout(bfn_2_12_0_));
    defparam IN_MUX_bfv_2_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_13_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15 ),
            .carryinitout(bfn_2_13_0_));
    defparam IN_MUX_bfv_1_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_7_0_));
    defparam IN_MUX_bfv_1_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_8_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_acc_1_cry_7 ),
            .carryinitout(bfn_1_8_0_));
    defparam IN_MUX_bfv_1_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_9_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_acc_1_cry_15 ),
            .carryinitout(bfn_1_9_0_));
    defparam IN_MUX_bfv_5_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_11_0_));
    defparam IN_MUX_bfv_5_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_12_0_ (
            .carryinitin(\pwm_generator_inst.un14_counter_cry_7 ),
            .carryinitout(bfn_5_12_0_));
    defparam IN_MUX_bfv_3_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_8_0_));
    defparam IN_MUX_bfv_3_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_9_0_ (
            .carryinitin(\pwm_generator_inst.un19_threshold_acc_cry_7 ),
            .carryinitout(bfn_3_9_0_));
    defparam IN_MUX_bfv_5_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_8_0_));
    defparam IN_MUX_bfv_5_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_9_0_ (
            .carryinitin(\pwm_generator_inst.counter_cry_7 ),
            .carryinitout(bfn_5_9_0_));
    defparam IN_MUX_bfv_9_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_13_0_));
    defparam IN_MUX_bfv_9_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_14_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryinitout(bfn_9_14_0_));
    defparam IN_MUX_bfv_9_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_15_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryinitout(bfn_9_15_0_));
    defparam IN_MUX_bfv_8_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_17_0_));
    defparam IN_MUX_bfv_8_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_18_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryinitout(bfn_8_18_0_));
    defparam IN_MUX_bfv_8_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_19_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryinitout(bfn_8_19_0_));
    defparam IN_MUX_bfv_15_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_11_0_));
    defparam IN_MUX_bfv_15_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_12_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_15_12_0_));
    defparam IN_MUX_bfv_15_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_13_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_15_13_0_));
    defparam IN_MUX_bfv_15_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_14_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_15_14_0_));
    defparam IN_MUX_bfv_17_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_11_0_));
    defparam IN_MUX_bfv_17_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_12_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .carryinitout(bfn_17_12_0_));
    defparam IN_MUX_bfv_17_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_13_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .carryinitout(bfn_17_13_0_));
    defparam IN_MUX_bfv_17_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_14_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .carryinitout(bfn_17_14_0_));
    defparam IN_MUX_bfv_14_26_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_26_0_));
    defparam IN_MUX_bfv_14_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_27_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_14_27_0_));
    defparam IN_MUX_bfv_14_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_28_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_14_28_0_));
    defparam IN_MUX_bfv_14_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_29_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_14_29_0_));
    defparam IN_MUX_bfv_14_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_21_0_));
    defparam IN_MUX_bfv_14_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_22_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .carryinitout(bfn_14_22_0_));
    defparam IN_MUX_bfv_14_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_23_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .carryinitout(bfn_14_23_0_));
    defparam IN_MUX_bfv_14_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_24_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .carryinitout(bfn_14_24_0_));
    defparam IN_MUX_bfv_18_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_18_0_));
    defparam IN_MUX_bfv_18_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_19_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_18_19_0_));
    defparam IN_MUX_bfv_18_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_20_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_18_20_0_));
    defparam IN_MUX_bfv_18_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_21_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_18_21_0_));
    defparam IN_MUX_bfv_17_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_15_0_));
    defparam IN_MUX_bfv_17_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_16_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_8 ),
            .carryinitout(bfn_17_16_0_));
    defparam IN_MUX_bfv_17_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_17_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_16 ),
            .carryinitout(bfn_17_17_0_));
    defparam IN_MUX_bfv_17_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_18_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_24 ),
            .carryinitout(bfn_17_18_0_));
    defparam IN_MUX_bfv_18_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_22_0_));
    defparam IN_MUX_bfv_18_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_23_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_7 ),
            .carryinitout(bfn_18_23_0_));
    defparam IN_MUX_bfv_18_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_24_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_15 ),
            .carryinitout(bfn_18_24_0_));
    defparam IN_MUX_bfv_18_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_25_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_23 ),
            .carryinitout(bfn_18_25_0_));
    defparam IN_MUX_bfv_14_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_15_0_));
    defparam IN_MUX_bfv_14_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_16_0_ (
            .carryinitin(\current_shift_inst.control_input_1_cry_7 ),
            .carryinitout(bfn_14_16_0_));
    defparam IN_MUX_bfv_14_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_17_0_ (
            .carryinitin(\current_shift_inst.control_input_1_cry_15 ),
            .carryinitout(bfn_14_17_0_));
    defparam IN_MUX_bfv_14_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_18_0_ (
            .carryinitin(\current_shift_inst.control_input_1_cry_23 ),
            .carryinitout(bfn_14_18_0_));
    defparam IN_MUX_bfv_14_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_7_0_));
    defparam IN_MUX_bfv_14_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_8_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_7 ),
            .carryinitout(bfn_14_8_0_));
    defparam IN_MUX_bfv_14_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_9_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15 ),
            .carryinitout(bfn_14_9_0_));
    defparam IN_MUX_bfv_14_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_10_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23 ),
            .carryinitout(bfn_14_10_0_));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_8_0_));
    defparam IN_MUX_bfv_9_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_9_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .carryinitout(bfn_9_9_0_));
    defparam IN_MUX_bfv_9_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_10_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .carryinitout(bfn_9_10_0_));
    defparam IN_MUX_bfv_9_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_11_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .carryinitout(bfn_9_11_0_));
    defparam IN_MUX_bfv_13_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_10_0_));
    defparam IN_MUX_bfv_13_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_11_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .carryinitout(bfn_13_11_0_));
    defparam IN_MUX_bfv_13_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_12_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_15 ),
            .carryinitout(bfn_13_12_0_));
    defparam IN_MUX_bfv_13_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_13_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_23 ),
            .carryinitout(bfn_13_13_0_));
    ICE_GB \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_0  (
            .USERSIGNALTOGLOBALBUFFER(N__22372),
            .GLOBALBUFFEROUTPUT(\delay_measurement_inst.delay_hc_timer.N_302_i_g ));
    ICE_GB \current_shift_inst.timer_s1.running_RNII51H_0  (
            .USERSIGNALTOGLOBALBUFFER(N__33295),
            .GLOBALBUFFEROUTPUT(\current_shift_inst.timer_s1.N_180_i_g ));
    ICE_GB \delay_measurement_inst.delay_tr_timer.running_RNICNBI_0  (
            .USERSIGNALTOGLOBALBUFFER(N__39223),
            .GLOBALBUFFEROUTPUT(\delay_measurement_inst.delay_tr_timer.N_304_i_g ));
    defparam osc.CLKHF_DIV="0b10";
    SB_HFOSC osc (
            .CLKHFPU(N__38086),
            .CLKHFEN(N__38087),
            .CLKHF(clk_12mhz));
    defparam rgb_drv.RGB2_CURRENT="0b111111";
    defparam rgb_drv.CURRENT_MODE="0b0";
    defparam rgb_drv.RGB0_CURRENT="0b111111";
    defparam rgb_drv.RGB1_CURRENT="0b111111";
    SB_RGBA_DRV rgb_drv (
            .RGBLEDEN(N__38162),
            .RGB2PWM(N__20059),
            .RGB1(rgb_g),
            .CURREN(N__38163),
            .RGB2(rgb_b),
            .RGB1PWM(N__20959),
            .RGB0PWM(N__49790),
            .RGB0(rgb_r));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_4_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_4_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_4_0 .LUT_INIT=16'b1010111000001110;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_5_LC_1_4_0  (
            .in0(N__24082),
            .in1(N__22820),
            .in2(N__24624),
            .in3(N__22743),
            .lcout(pwm_duty_input_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50278),
            .ce(),
            .sr(N__49667));
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_4_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_4_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_4_6 .LUT_INIT=16'b1010111000001110;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_8_LC_1_4_6  (
            .in0(N__23989),
            .in1(N__22821),
            .in2(N__24625),
            .in3(N__22744),
            .lcout(pwm_duty_input_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50278),
            .ce(),
            .sr(N__49667));
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_5_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_5_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_5_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_1_LC_1_5_0  (
            .in0(_gnd_net_),
            .in1(N__23788),
            .in2(_gnd_net_),
            .in3(N__20190),
            .lcout(pwm_duty_input_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50277),
            .ce(),
            .sr(N__49674));
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_5_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_5_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_5_1 .LUT_INIT=16'b0010001100110011;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_4_LC_1_5_1  (
            .in0(N__24130),
            .in1(N__20950),
            .in2(N__20170),
            .in3(N__22742),
            .lcout(pwm_duty_input_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50277),
            .ce(),
            .sr(N__49674));
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_5_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_5_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_5_3 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_3_LC_1_5_3  (
            .in0(N__23755),
            .in1(N__20200),
            .in2(_gnd_net_),
            .in3(N__20152),
            .lcout(pwm_duty_input_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50277),
            .ce(),
            .sr(N__49674));
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_5_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_5_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_5_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_2_LC_1_5_5  (
            .in0(N__20191),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23773),
            .lcout(pwm_duty_input_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50277),
            .ce(),
            .sr(N__49674));
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_5_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_5_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_5_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_0_LC_1_5_6  (
            .in0(_gnd_net_),
            .in1(N__23803),
            .in2(_gnd_net_),
            .in3(N__20189),
            .lcout(pwm_duty_input_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50277),
            .ce(),
            .sr(N__49674));
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_1  (
            .in0(N__24601),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_19_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50276),
            .ce(),
            .sr(N__49681));
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_6_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_6_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_6_3 .LUT_INIT=16'b1010111000001110;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_6_LC_1_6_3  (
            .in0(N__24049),
            .in1(N__22815),
            .in2(N__24616),
            .in3(N__22745),
            .lcout(pwm_duty_input_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50276),
            .ce(),
            .sr(N__49681));
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_6_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_6_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_6_4 .LUT_INIT=16'b1011101100110000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_9_LC_1_6_4  (
            .in0(N__22747),
            .in1(N__24608),
            .in2(N__22822),
            .in3(N__23956),
            .lcout(pwm_duty_input_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50276),
            .ce(),
            .sr(N__49681));
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_6_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_6_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_6_5 .LUT_INIT=16'b1010111000001110;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_7_LC_1_6_5  (
            .in0(N__24019),
            .in1(N__22816),
            .in2(N__24617),
            .in3(N__22746),
            .lcout(pwm_duty_input_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50276),
            .ce(),
            .sr(N__49681));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_1_7_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_1_7_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_1_7_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_1_7_0  (
            .in0(_gnd_net_),
            .in1(N__19759),
            .in2(_gnd_net_),
            .in3(N__19771),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_0 ),
            .ltout(),
            .carryin(bfn_1_7_0_),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_1_7_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_1_7_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_1_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_1_7_1  (
            .in0(_gnd_net_),
            .in1(N__19741),
            .in2(_gnd_net_),
            .in3(N__19753),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_0 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_1_7_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_1_7_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_1_7_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_1_7_2  (
            .in0(_gnd_net_),
            .in1(N__19726),
            .in2(_gnd_net_),
            .in3(N__19735),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_1 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_1_7_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_1_7_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_1_7_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_1_7_3  (
            .in0(_gnd_net_),
            .in1(N__19711),
            .in2(_gnd_net_),
            .in3(N__19720),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_2 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_1_7_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_1_7_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_1_7_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_1_7_4  (
            .in0(N__19705),
            .in1(N__19696),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_3 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_1_7_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_1_7_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_1_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_1_7_5  (
            .in0(_gnd_net_),
            .in1(N__19681),
            .in2(_gnd_net_),
            .in3(N__19690),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_4 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_1_7_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_1_7_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_1_7_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_1_7_6  (
            .in0(_gnd_net_),
            .in1(N__19663),
            .in2(_gnd_net_),
            .in3(N__19675),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_5 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_1_7_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_1_7_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_1_7_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_1_7_7  (
            .in0(_gnd_net_),
            .in1(N__19645),
            .in2(_gnd_net_),
            .in3(N__19657),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_6 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_1_8_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_1_8_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_1_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_1_8_0  (
            .in0(_gnd_net_),
            .in1(N__19810),
            .in2(_gnd_net_),
            .in3(N__19822),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_8 ),
            .ltout(),
            .carryin(bfn_1_8_0_),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_1_8_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_1_8_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_1_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_1_8_1  (
            .in0(_gnd_net_),
            .in1(N__19795),
            .in2(_gnd_net_),
            .in3(N__19804),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_8 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_1_8_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_1_8_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_1_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_1_8_2  (
            .in0(_gnd_net_),
            .in1(N__20631),
            .in2(_gnd_net_),
            .in3(N__19789),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_9 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_1_8_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_1_8_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_1_8_3 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_1_8_3  (
            .in0(N__21290),
            .in1(N__19855),
            .in2(_gnd_net_),
            .in3(N__19786),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_10 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_1_8_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_1_8_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_1_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_1_8_4  (
            .in0(_gnd_net_),
            .in1(N__20138),
            .in2(_gnd_net_),
            .in3(N__19783),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_11 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_1_8_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_1_8_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_1_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_1_8_5  (
            .in0(_gnd_net_),
            .in1(N__20576),
            .in2(_gnd_net_),
            .in3(N__19780),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_12 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_1_8_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_1_8_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_1_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_1_8_6  (
            .in0(_gnd_net_),
            .in1(N__20373),
            .in2(_gnd_net_),
            .in3(N__19777),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_13 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_1_8_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_1_8_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_1_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_1_8_7  (
            .in0(_gnd_net_),
            .in1(N__20336),
            .in2(_gnd_net_),
            .in3(N__19774),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_14 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_1_9_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_1_9_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_1_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_1_9_0  (
            .in0(_gnd_net_),
            .in1(N__20288),
            .in2(_gnd_net_),
            .in3(N__19867),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_1_9_0_),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_1_9_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_1_9_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_1_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_1_9_1  (
            .in0(_gnd_net_),
            .in1(N__20259),
            .in2(_gnd_net_),
            .in3(N__19864),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_16 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_1_9_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_1_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_1_9_2  (
            .in0(_gnd_net_),
            .in1(N__20229),
            .in2(_gnd_net_),
            .in3(N__19861),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_17 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_1_9_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_1_9_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_1_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_1_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19858),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_1_9_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_1_9_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_1_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_1_9_4  (
            .in0(_gnd_net_),
            .in1(N__20289),
            .in2(_gnd_net_),
            .in3(N__20271),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_1_9_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_1_9_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_1_9_5 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_1_9_5  (
            .in0(_gnd_net_),
            .in1(N__20106),
            .in2(_gnd_net_),
            .in3(N__20140),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_1_9_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_1_9_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_1_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_1_9_6  (
            .in0(N__20338),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20307),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_10_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_10_0  (
            .in0(_gnd_net_),
            .in1(N__19854),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_10_0_),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_10_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_10_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_10_1  (
            .in0(_gnd_net_),
            .in1(N__19837),
            .in2(_gnd_net_),
            .in3(N__19825),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_0 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_10_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_10_2  (
            .in0(_gnd_net_),
            .in1(N__19912),
            .in2(_gnd_net_),
            .in3(N__19900),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_1 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_10_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_10_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_10_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_10_3  (
            .in0(_gnd_net_),
            .in1(N__19897),
            .in2(_gnd_net_),
            .in3(N__19885),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_2 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_10_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_10_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_10_4  (
            .in0(_gnd_net_),
            .in1(N__20530),
            .in2(_gnd_net_),
            .in3(N__19882),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_3 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_10_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_10_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_10_5  (
            .in0(_gnd_net_),
            .in1(N__38339),
            .in2(N__20497),
            .in3(N__19879),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_4 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_10_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_10_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_10_6  (
            .in0(_gnd_net_),
            .in1(N__20458),
            .in2(N__38386),
            .in3(N__19876),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_5 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_10_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_10_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_10_7  (
            .in0(_gnd_net_),
            .in1(N__20419),
            .in2(N__38387),
            .in3(N__19873),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_6 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_11_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(N__20383),
            .in2(_gnd_net_),
            .in3(N__19870),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9 ),
            .ltout(),
            .carryin(bfn_1_11_0_),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_11_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_11_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(N__20848),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_8 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_11_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_11_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(N__20812),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_9 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_11_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_11_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(N__20776),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_10 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_11_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_11_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_11_4  (
            .in0(_gnd_net_),
            .in1(N__20737),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_11 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_11_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_11_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_11_5  (
            .in0(_gnd_net_),
            .in1(N__20701),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_12 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_11_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_11_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_11_6  (
            .in0(_gnd_net_),
            .in1(N__20677),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_13 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_11_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_11_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_11_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_11_7  (
            .in0(_gnd_net_),
            .in1(N__20656),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_14 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_12_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_12_0  (
            .in0(_gnd_net_),
            .in1(N__21097),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_12_0_),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_12_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_12_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_12_1  (
            .in0(_gnd_net_),
            .in1(N__21076),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_16 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_12_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_12_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_12_2  (
            .in0(_gnd_net_),
            .in1(N__21052),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_17 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_12_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_12_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_12_3  (
            .in0(_gnd_net_),
            .in1(N__20986),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_18 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_12_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20086),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_12_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_12_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_12_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_12_5  (
            .in0(N__20079),
            .in1(N__21033),
            .in2(_gnd_net_),
            .in3(N__21601),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_13_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_13_1 .LUT_INIT=16'b1001011000111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_13_1  (
            .in0(N__20083),
            .in1(N__21037),
            .in2(N__20068),
            .in3(N__21568),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_drv_RNO_0_LC_1_30_5.C_ON=1'b0;
    defparam rgb_drv_RNO_0_LC_1_30_5.SEQ_MODE=4'b0000;
    defparam rgb_drv_RNO_0_LC_1_30_5.LUT_INIT=16'b1100110000110011;
    LogicCell40 rgb_drv_RNO_0_LC_1_30_5 (
            .in0(_gnd_net_),
            .in1(N__22333),
            .in2(_gnd_net_),
            .in3(N__49789),
            .lcout(N_34_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_5_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_5_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_5_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_5_0  (
            .in0(N__19983),
            .in1(N__19927),
            .in2(N__20005),
            .in3(N__19945),
            .lcout(),
            .ltout(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_5_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_5_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_5_1 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_5_1  (
            .in0(N__19965),
            .in1(N__20935),
            .in2(N__20053),
            .in3(N__20901),
            .lcout(\pwm_generator_inst.N_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_5_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_5_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_5_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pwm_generator_inst.un1_duty_inputlto2_LC_2_5_2  (
            .in0(N__20049),
            .in1(N__20034),
            .in2(_gnd_net_),
            .in3(N__20019),
            .lcout(\pwm_generator_inst.un1_duty_inputlt3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_5_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_5_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_5_3 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_5_3  (
            .in0(_gnd_net_),
            .in1(N__20001),
            .in2(_gnd_net_),
            .in3(N__19982),
            .lcout(),
            .ltout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_5_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_5_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_5_4 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_5_4  (
            .in0(N__19964),
            .in1(N__19944),
            .in2(N__19930),
            .in3(N__19926),
            .lcout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_2_5_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_2_5_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_2_5_5 .LUT_INIT=16'b0000000000001101;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_2_5_5  (
            .in0(N__24136),
            .in1(N__21181),
            .in2(N__24614),
            .in3(N__22813),
            .lcout(\current_shift_inst.PI_CTRL.N_164 ),
            .ltout(\current_shift_inst.PI_CTRL.N_164_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_2_5_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_2_5_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_2_5_6 .LUT_INIT=16'b1111111111011100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_2_5_6  (
            .in0(N__23751),
            .in1(N__20179),
            .in2(N__20194),
            .in3(N__20151),
            .lcout(\current_shift_inst.PI_CTRL.N_120 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_5_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_5_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_5_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_5_7  (
            .in0(N__24593),
            .in1(N__21180),
            .in2(_gnd_net_),
            .in3(N__22812),
            .lcout(\current_shift_inst.PI_CTRL.N_167 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_6_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_6_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_6_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_6_0  (
            .in0(_gnd_net_),
            .in1(N__24131),
            .in2(_gnd_net_),
            .in3(N__23744),
            .lcout(\current_shift_inst.PI_CTRL.N_168 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_2_6_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_2_6_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_2_6_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_2_6_4  (
            .in0(_gnd_net_),
            .in1(N__24077),
            .in2(_gnd_net_),
            .in3(N__23985),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_6_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_6_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_6_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_6_5  (
            .in0(N__23955),
            .in1(N__24018),
            .in2(N__20173),
            .in3(N__24048),
            .lcout(\current_shift_inst.PI_CTRL.N_27 ),
            .ltout(\current_shift_inst.PI_CTRL.N_27_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_6_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_6_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_6_6 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_6_6  (
            .in0(N__24600),
            .in1(N__20161),
            .in2(N__20155),
            .in3(N__22726),
            .lcout(\current_shift_inst.PI_CTRL.N_166 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_8_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_8_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_8_0 .LUT_INIT=16'b1101011110000010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_8_0  (
            .in0(N__21295),
            .in1(N__20139),
            .in2(N__20122),
            .in3(N__20113),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_8_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_8_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_8_1 .LUT_INIT=16'b1010010111001100;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_8_1  (
            .in0(N__20581),
            .in1(N__20596),
            .in2(N__20095),
            .in3(N__21297),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_2_8_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_2_8_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_2_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_2_8_3  (
            .in0(_gnd_net_),
            .in1(N__20374),
            .in2(_gnd_net_),
            .in3(N__20352),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ),
            .ltout(\pwm_generator_inst.un15_threshold_acc_1_axb_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_8_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_8_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_8_4 .LUT_INIT=16'b1101011110000010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_8_4  (
            .in0(N__21296),
            .in1(N__20362),
            .in2(N__20356),
            .in3(N__20353),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_8_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_8_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_8_6 .LUT_INIT=16'b1101011110000010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_8_6  (
            .in0(N__21298),
            .in1(N__20337),
            .in2(N__20320),
            .in3(N__20311),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_9_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_9_0 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_9_0  (
            .in0(N__20296),
            .in1(N__20290),
            .in2(N__20275),
            .in3(N__21292),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_9_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_9_1  (
            .in0(N__20260),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20247),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ),
            .ltout(\pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_9_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_9_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_9_2 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_9_2  (
            .in0(N__20248),
            .in1(N__20239),
            .in2(N__20233),
            .in3(N__21293),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_9_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_9_3  (
            .in0(N__20230),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20217),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ),
            .ltout(\pwm_generator_inst.un15_threshold_acc_1_axb_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_9_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_9_4 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_9_4  (
            .in0(N__20218),
            .in1(N__20209),
            .in2(N__20203),
            .in3(N__21294),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_2_9_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_2_9_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_2_9_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_2_9_5  (
            .in0(_gnd_net_),
            .in1(N__20632),
            .in2(_gnd_net_),
            .in3(N__20619),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ),
            .ltout(\pwm_generator_inst.un15_threshold_acc_1_axb_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_9_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_9_6 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_9_6  (
            .in0(N__20620),
            .in1(N__20605),
            .in2(N__20599),
            .in3(N__21291),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_9_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_9_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_9_7  (
            .in0(N__20580),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20592),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_axb_4_LC_2_11_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_axb_4_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_axb_4_LC_2_11_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_axb_4_LC_2_11_0  (
            .in0(_gnd_net_),
            .in1(N__20560),
            .in2(N__20548),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un3_threshold_acc_axbZ0Z_4 ),
            .ltout(),
            .carryin(bfn_2_11_0_),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_2_11_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_2_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_2_11_1  (
            .in0(_gnd_net_),
            .in1(N__20524),
            .in2(N__20512),
            .in3(N__20488),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_2_11_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_2_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_2_11_2  (
            .in0(_gnd_net_),
            .in1(N__20485),
            .in2(N__20473),
            .in3(N__20452),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_2_11_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_2_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_2_11_3  (
            .in0(_gnd_net_),
            .in1(N__20449),
            .in2(N__20434),
            .in3(N__20413),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_2_11_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_2_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_2_11_4  (
            .in0(_gnd_net_),
            .in1(N__20410),
            .in2(N__20398),
            .in3(N__20377),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_2_11_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_2_11_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_2_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_2_11_5  (
            .in0(_gnd_net_),
            .in1(N__20875),
            .in2(N__20863),
            .in3(N__20842),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_2_11_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_2_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_2_11_6  (
            .in0(_gnd_net_),
            .in1(N__20839),
            .in2(N__20827),
            .in3(N__20806),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_2_11_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_2_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_2_11_7  (
            .in0(_gnd_net_),
            .in1(N__20803),
            .in2(N__20791),
            .in3(N__20770),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_2_12_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_2_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_2_12_0  (
            .in0(_gnd_net_),
            .in1(N__20767),
            .in2(N__20752),
            .in3(N__20731),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0 ),
            .ltout(),
            .carryin(bfn_2_12_0_),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_2_12_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_2_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_2_12_1  (
            .in0(_gnd_net_),
            .in1(N__20728),
            .in2(N__20716),
            .in3(N__20695),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_2_12_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_2_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_2_12_2  (
            .in0(_gnd_net_),
            .in1(N__21018),
            .in2(N__20692),
            .in3(N__20671),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_2_12_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_2_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_2_12_3  (
            .in0(_gnd_net_),
            .in1(N__20668),
            .in2(N__21034),
            .in3(N__20650),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_2_12_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_2_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_2_12_4  (
            .in0(_gnd_net_),
            .in1(N__21022),
            .in2(N__20647),
            .in3(N__21091),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_2_12_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_2_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_2_12_5  (
            .in0(_gnd_net_),
            .in1(N__21088),
            .in2(N__21035),
            .in3(N__21070),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_2_12_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_2_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_2_12_6  (
            .in0(_gnd_net_),
            .in1(N__21026),
            .in2(N__21067),
            .in3(N__21046),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_2_12_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_2_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_2_12_7  (
            .in0(_gnd_net_),
            .in1(N__21043),
            .in2(N__21036),
            .in3(N__20980),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_2_13_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_2_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_2_13_0  (
            .in0(_gnd_net_),
            .in1(N__20977),
            .in2(N__20971),
            .in3(N__20962),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rgb_drv_RNO_LC_2_30_7.C_ON=1'b0;
    defparam rgb_drv_RNO_LC_2_30_7.SEQ_MODE=4'b0000;
    defparam rgb_drv_RNO_LC_2_30_7.LUT_INIT=16'b0000000011001100;
    LogicCell40 rgb_drv_RNO_LC_2_30_7 (
            .in0(_gnd_net_),
            .in1(N__22332),
            .in2(_gnd_net_),
            .in3(N__49788),
            .lcout(rgb_drv_RNOZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_3_5_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_3_5_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_3_5_3 .LUT_INIT=16'b0000111100000111;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_3_5_3  (
            .in0(N__24135),
            .in1(N__21179),
            .in2(N__24615),
            .in3(N__22814),
            .lcout(\current_shift_inst.PI_CTRL.N_162 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_3_5_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_3_5_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_3_5_7 .LUT_INIT=16'b1010101011111011;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_LC_3_5_7  (
            .in0(N__20941),
            .in1(N__20934),
            .in2(N__20911),
            .in3(N__20900),
            .lcout(\pwm_generator_inst.N_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_6_LC_3_6_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_6_LC_3_6_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_6_LC_3_6_2 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_6_LC_3_6_2  (
            .in0(_gnd_net_),
            .in1(N__23984),
            .in2(_gnd_net_),
            .in3(N__24047),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_3_6_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_3_6_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_3_6_3 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_3_6_3  (
            .in0(N__23948),
            .in1(N__24017),
            .in2(N__21184),
            .in3(N__24078),
            .lcout(\current_shift_inst.PI_CTRL.N_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_3_8_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_3_8_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_3_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_3_8_0  (
            .in0(_gnd_net_),
            .in1(N__21163),
            .in2(N__21304),
            .in3(N__21303),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(bfn_3_8_0_),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_3_8_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_3_8_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_3_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_3_8_1  (
            .in0(_gnd_net_),
            .in1(N__21157),
            .in2(_gnd_net_),
            .in3(N__21148),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_0 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_3_8_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_3_8_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_3_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_3_8_2  (
            .in0(_gnd_net_),
            .in1(N__21145),
            .in2(_gnd_net_),
            .in3(N__21139),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_1 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_3_8_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_3_8_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_3_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_3_8_3  (
            .in0(_gnd_net_),
            .in1(N__21136),
            .in2(_gnd_net_),
            .in3(N__21130),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_2 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_3_8_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_3_8_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_3_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_3_8_4  (
            .in0(_gnd_net_),
            .in1(N__21127),
            .in2(_gnd_net_),
            .in3(N__21121),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_3 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_3_8_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_3_8_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_3_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_3_8_5  (
            .in0(_gnd_net_),
            .in1(N__21118),
            .in2(_gnd_net_),
            .in3(N__21112),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_4 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_3_8_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_3_8_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_3_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_3_8_6  (
            .in0(_gnd_net_),
            .in1(N__21109),
            .in2(_gnd_net_),
            .in3(N__21100),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_5 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_3_8_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_3_8_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_3_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_3_8_7  (
            .in0(_gnd_net_),
            .in1(N__21334),
            .in2(_gnd_net_),
            .in3(N__21328),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_6 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_3_9_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_3_9_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_3_9_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_3_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21325),
            .in3(N__21316),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(bfn_3_9_0_),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_3_9_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_3_9_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_3_9_1 .LUT_INIT=16'b1000011101111000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_3_9_1  (
            .in0(N__21313),
            .in1(N__21302),
            .in2(N__21235),
            .in3(N__21220),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_9_LC_3_10_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_9_LC_3_10_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_9_LC_3_10_0 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_9_LC_3_10_0  (
            .in0(N__21624),
            .in1(N__21413),
            .in2(N__21217),
            .in3(N__21462),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50264),
            .ce(),
            .sr(N__49693));
    defparam \pwm_generator_inst.threshold_ACC_8_LC_3_10_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_8_LC_3_10_1 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_8_LC_3_10_1 .LUT_INIT=16'b1100111111011101;
    LogicCell40 \pwm_generator_inst.threshold_ACC_8_LC_3_10_1  (
            .in0(N__21461),
            .in1(N__21208),
            .in2(N__21418),
            .in3(N__21625),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50264),
            .ce(),
            .sr(N__49693));
    defparam \pwm_generator_inst.threshold_8_LC_3_11_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_8_LC_3_11_6 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_8_LC_3_11_6 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pwm_generator_inst.threshold_8_LC_3_11_6  (
            .in0(_gnd_net_),
            .in1(N__21202),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.thresholdZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50260),
            .ce(),
            .sr(N__49701));
    defparam CONSTANT_ONE_LUT4_LC_3_24_5.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_3_24_5.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_3_24_5.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_3_24_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_4_LC_4_8_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_4_LC_4_8_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_4_LC_4_8_2 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_4_LC_4_8_2  (
            .in0(N__21620),
            .in1(N__21395),
            .in2(N__21463),
            .in3(N__21196),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50269),
            .ce(),
            .sr(N__49675));
    defparam \pwm_generator_inst.threshold_4_LC_4_8_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_4_LC_4_8_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_4_LC_4_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_4_LC_4_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21190),
            .lcout(\pwm_generator_inst.thresholdZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50269),
            .ce(),
            .sr(N__49675));
    defparam \pwm_generator_inst.threshold_ACC_3_LC_4_8_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_3_LC_4_8_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_3_LC_4_8_7 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_3_LC_4_8_7  (
            .in0(N__21394),
            .in1(N__21444),
            .in2(N__21628),
            .in3(N__21664),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50269),
            .ce(),
            .sr(N__49675));
    defparam \pwm_generator_inst.threshold_ACC_0_LC_4_9_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_0_LC_4_9_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_0_LC_4_9_0 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_0_LC_4_9_0  (
            .in0(N__21610),
            .in1(N__21464),
            .in2(N__21414),
            .in3(N__21658),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50265),
            .ce(),
            .sr(N__49682));
    defparam \pwm_generator_inst.threshold_ACC_7_LC_4_9_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_7_LC_4_9_2 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_7_LC_4_9_2 .LUT_INIT=16'b1111111100011011;
    LogicCell40 \pwm_generator_inst.threshold_ACC_7_LC_4_9_2  (
            .in0(N__21613),
            .in1(N__21469),
            .in2(N__21417),
            .in3(N__21652),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50265),
            .ce(),
            .sr(N__49682));
    defparam \pwm_generator_inst.threshold_ACC_6_LC_4_9_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_6_LC_4_9_3 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_6_LC_4_9_3 .LUT_INIT=16'b1111111100110101;
    LogicCell40 \pwm_generator_inst.threshold_ACC_6_LC_4_9_3  (
            .in0(N__21468),
            .in1(N__21406),
            .in2(N__21627),
            .in3(N__21646),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50265),
            .ce(),
            .sr(N__49682));
    defparam \pwm_generator_inst.threshold_ACC_1_LC_4_9_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_1_LC_4_9_4 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_1_LC_4_9_4 .LUT_INIT=16'b1111111100011011;
    LogicCell40 \pwm_generator_inst.threshold_ACC_1_LC_4_9_4  (
            .in0(N__21611),
            .in1(N__21465),
            .in2(N__21415),
            .in3(N__21640),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50265),
            .ce(),
            .sr(N__49682));
    defparam \pwm_generator_inst.threshold_ACC_5_LC_4_9_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_5_LC_4_9_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_5_LC_4_9_5 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_5_LC_4_9_5  (
            .in0(N__21467),
            .in1(N__21405),
            .in2(N__21626),
            .in3(N__21634),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50265),
            .ce(),
            .sr(N__49682));
    defparam \pwm_generator_inst.threshold_ACC_2_LC_4_9_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_2_LC_4_9_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_2_LC_4_9_6 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_2_LC_4_9_6  (
            .in0(N__21612),
            .in1(N__21466),
            .in2(N__21416),
            .in3(N__21352),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50265),
            .ce(),
            .sr(N__49682));
    defparam \pwm_generator_inst.threshold_1_LC_4_10_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_1_LC_4_10_1 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_1_LC_4_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_1_LC_4_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21346),
            .lcout(\pwm_generator_inst.thresholdZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50261),
            .ce(),
            .sr(N__49688));
    defparam \pwm_generator_inst.threshold_6_LC_4_10_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_6_LC_4_10_3 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_6_LC_4_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_6_LC_4_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21340),
            .lcout(\pwm_generator_inst.thresholdZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50261),
            .ce(),
            .sr(N__49688));
    defparam \pwm_generator_inst.threshold_7_LC_4_10_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_7_LC_4_10_5 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_7_LC_4_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_7_LC_4_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21712),
            .lcout(\pwm_generator_inst.thresholdZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50261),
            .ce(),
            .sr(N__49688));
    defparam \pwm_generator_inst.threshold_5_LC_4_11_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_5_LC_4_11_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_5_LC_4_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_5_LC_4_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21706),
            .lcout(\pwm_generator_inst.thresholdZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50254),
            .ce(),
            .sr(N__49694));
    defparam \pwm_generator_inst.threshold_2_LC_4_11_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_2_LC_4_11_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_2_LC_4_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_2_LC_4_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21697),
            .lcout(\pwm_generator_inst.thresholdZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50254),
            .ce(),
            .sr(N__49694));
    defparam \pwm_generator_inst.threshold_3_LC_4_11_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_3_LC_4_11_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_3_LC_4_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_3_LC_4_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21688),
            .lcout(\pwm_generator_inst.thresholdZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50254),
            .ce(),
            .sr(N__49694));
    defparam \pwm_generator_inst.threshold_9_LC_4_11_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_9_LC_4_11_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_9_LC_4_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_9_LC_4_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21679),
            .lcout(\pwm_generator_inst.thresholdZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50254),
            .ce(),
            .sr(N__49694));
    defparam \phase_controller_inst1.state_1_LC_4_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_1_LC_4_17_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_1_LC_4_17_3 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \phase_controller_inst1.state_1_LC_4_17_3  (
            .in0(N__22591),
            .in1(N__22625),
            .in2(N__26051),
            .in3(N__23884),
            .lcout(\phase_controller_inst1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50215),
            .ce(),
            .sr(N__49732));
    defparam \pwm_generator_inst.counter_0_LC_5_8_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_0_LC_5_8_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_0_LC_5_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_0_LC_5_8_0  (
            .in0(N__21985),
            .in1(N__21923),
            .in2(_gnd_net_),
            .in3(N__21673),
            .lcout(\pwm_generator_inst.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_5_8_0_),
            .carryout(\pwm_generator_inst.counter_cry_0 ),
            .clk(N__50266),
            .ce(),
            .sr(N__49668));
    defparam \pwm_generator_inst.counter_1_LC_5_8_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_1_LC_5_8_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_1_LC_5_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_1_LC_5_8_1  (
            .in0(N__21981),
            .in1(N__21884),
            .in2(_gnd_net_),
            .in3(N__21670),
            .lcout(\pwm_generator_inst.counterZ0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_0 ),
            .carryout(\pwm_generator_inst.counter_cry_1 ),
            .clk(N__50266),
            .ce(),
            .sr(N__49668));
    defparam \pwm_generator_inst.counter_2_LC_5_8_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_2_LC_5_8_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_2_LC_5_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_2_LC_5_8_2  (
            .in0(N__21986),
            .in1(N__21845),
            .in2(_gnd_net_),
            .in3(N__21667),
            .lcout(\pwm_generator_inst.counterZ0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_1 ),
            .carryout(\pwm_generator_inst.counter_cry_2 ),
            .clk(N__50266),
            .ce(),
            .sr(N__49668));
    defparam \pwm_generator_inst.counter_3_LC_5_8_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_3_LC_5_8_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_3_LC_5_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_3_LC_5_8_3  (
            .in0(N__21982),
            .in1(N__21809),
            .in2(_gnd_net_),
            .in3(N__21739),
            .lcout(\pwm_generator_inst.counterZ0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_2 ),
            .carryout(\pwm_generator_inst.counter_cry_3 ),
            .clk(N__50266),
            .ce(),
            .sr(N__49668));
    defparam \pwm_generator_inst.counter_4_LC_5_8_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_4_LC_5_8_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_4_LC_5_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_4_LC_5_8_4  (
            .in0(N__21987),
            .in1(N__21764),
            .in2(_gnd_net_),
            .in3(N__21736),
            .lcout(\pwm_generator_inst.counterZ0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_3 ),
            .carryout(\pwm_generator_inst.counter_cry_4 ),
            .clk(N__50266),
            .ce(),
            .sr(N__49668));
    defparam \pwm_generator_inst.counter_5_LC_5_8_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_5_LC_5_8_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_5_LC_5_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_5_LC_5_8_5  (
            .in0(N__21983),
            .in1(N__22196),
            .in2(_gnd_net_),
            .in3(N__21733),
            .lcout(\pwm_generator_inst.counterZ0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_4 ),
            .carryout(\pwm_generator_inst.counter_cry_5 ),
            .clk(N__50266),
            .ce(),
            .sr(N__49668));
    defparam \pwm_generator_inst.counter_6_LC_5_8_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_6_LC_5_8_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_6_LC_5_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_6_LC_5_8_6  (
            .in0(N__21988),
            .in1(N__22169),
            .in2(_gnd_net_),
            .in3(N__21730),
            .lcout(\pwm_generator_inst.counterZ0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_5 ),
            .carryout(\pwm_generator_inst.counter_cry_6 ),
            .clk(N__50266),
            .ce(),
            .sr(N__49668));
    defparam \pwm_generator_inst.counter_7_LC_5_8_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_7_LC_5_8_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_7_LC_5_8_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_7_LC_5_8_7  (
            .in0(N__21984),
            .in1(N__22124),
            .in2(_gnd_net_),
            .in3(N__21727),
            .lcout(\pwm_generator_inst.counterZ0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_6 ),
            .carryout(\pwm_generator_inst.counter_cry_7 ),
            .clk(N__50266),
            .ce(),
            .sr(N__49668));
    defparam \pwm_generator_inst.counter_8_LC_5_9_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_8_LC_5_9_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_8_LC_5_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_8_LC_5_9_0  (
            .in0(N__21980),
            .in1(N__22079),
            .in2(_gnd_net_),
            .in3(N__21724),
            .lcout(\pwm_generator_inst.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_5_9_0_),
            .carryout(\pwm_generator_inst.counter_cry_8 ),
            .clk(N__50262),
            .ce(),
            .sr(N__49676));
    defparam \pwm_generator_inst.counter_9_LC_5_9_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_9_LC_5_9_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_9_LC_5_9_1 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \pwm_generator_inst.counter_9_LC_5_9_1  (
            .in0(N__22041),
            .in1(N__21979),
            .in2(_gnd_net_),
            .in3(N__21721),
            .lcout(\pwm_generator_inst.counterZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50262),
            .ce(),
            .sr(N__49676));
    defparam \pwm_generator_inst.threshold_0_LC_5_9_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_0_LC_5_9_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_0_LC_5_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_0_LC_5_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21718),
            .lcout(\pwm_generator_inst.thresholdZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50262),
            .ce(),
            .sr(N__49676));
    defparam \pwm_generator_inst.counter_RNITBL3_9_LC_5_10_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNITBL3_9_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNITBL3_9_LC_5_10_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNITBL3_9_LC_5_10_2  (
            .in0(N__22198),
            .in1(N__22040),
            .in2(_gnd_net_),
            .in3(N__22080),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlto9_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIFA6C_6_LC_5_10_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIFA6C_6_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIFA6C_6_LC_5_10_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \pwm_generator_inst.counter_RNIFA6C_6_LC_5_10_3  (
            .in0(N__22126),
            .in1(N__22171),
            .in2(N__21991),
            .in3(N__21943),
            .lcout(\pwm_generator_inst.un1_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIRPD2_0_LC_5_10_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIRPD2_0_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIRPD2_0_LC_5_10_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIRPD2_0_LC_5_10_6  (
            .in0(_gnd_net_),
            .in1(N__21885),
            .in2(_gnd_net_),
            .in3(N__21924),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlto2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIBO26_2_LC_5_10_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIBO26_2_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIBO26_2_LC_5_10_7 .LUT_INIT=16'b0000000000010011;
    LogicCell40 \pwm_generator_inst.counter_RNIBO26_2_LC_5_10_7  (
            .in0(N__21847),
            .in1(N__21766),
            .in2(N__21946),
            .in3(N__21811),
            .lcout(\pwm_generator_inst.un1_counterlt9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_5_11_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_5_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_5_11_0  (
            .in0(_gnd_net_),
            .in1(N__21901),
            .in2(N__21937),
            .in3(N__21925),
            .lcout(\pwm_generator_inst.counter_i_0 ),
            .ltout(),
            .carryin(bfn_5_11_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_5_11_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_5_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_5_11_1  (
            .in0(_gnd_net_),
            .in1(N__21862),
            .in2(N__21895),
            .in3(N__21886),
            .lcout(\pwm_generator_inst.counter_i_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_0 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_5_11_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_5_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_5_11_2  (
            .in0(_gnd_net_),
            .in1(N__21826),
            .in2(N__21856),
            .in3(N__21846),
            .lcout(\pwm_generator_inst.counter_i_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_1 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_5_11_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_5_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_5_11_3  (
            .in0(_gnd_net_),
            .in1(N__21790),
            .in2(N__21820),
            .in3(N__21810),
            .lcout(\pwm_generator_inst.counter_i_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_2 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_5_11_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_5_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_5_11_4  (
            .in0(_gnd_net_),
            .in1(N__21745),
            .in2(N__21781),
            .in3(N__21765),
            .lcout(\pwm_generator_inst.counter_i_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_3 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_5_11_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_5_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_5_11_5  (
            .in0(_gnd_net_),
            .in1(N__22177),
            .in2(N__22207),
            .in3(N__22197),
            .lcout(\pwm_generator_inst.counter_i_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_4 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_5_11_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_5_11_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_5_11_6  (
            .in0(N__22170),
            .in1(N__22141),
            .in2(N__22150),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_5 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_5_11_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_5_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_5_11_7  (
            .in0(_gnd_net_),
            .in1(N__22102),
            .in2(N__22135),
            .in3(N__22125),
            .lcout(\pwm_generator_inst.counter_i_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_6 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_5_12_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_5_12_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_5_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_5_12_0  (
            .in0(_gnd_net_),
            .in1(N__22057),
            .in2(N__22096),
            .in3(N__22081),
            .lcout(\pwm_generator_inst.counter_i_8 ),
            .ltout(),
            .carryin(bfn_5_12_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_5_12_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_5_12_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_5_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_5_12_1  (
            .in0(_gnd_net_),
            .in1(N__22021),
            .in2(N__22051),
            .in3(N__22042),
            .lcout(\pwm_generator_inst.counter_i_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_8 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.pwm_out_LC_5_12_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.pwm_out_LC_5_12_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.pwm_out_LC_5_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.pwm_out_LC_5_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22015),
            .lcout(pwm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50242),
            .ce(),
            .sr(N__49695));
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_5_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_5_13_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_1_LC_5_13_5  (
            .in0(_gnd_net_),
            .in1(N__32122),
            .in2(_gnd_net_),
            .in3(N__22259),
            .lcout(\phase_controller_inst1.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_ns_i_a3_1_LC_5_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_ns_i_a3_1_LC_5_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_ns_i_a3_1_LC_5_14_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.state_ns_i_a3_1_LC_5_14_5  (
            .in0(N__22316),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25109),
            .lcout(state_ns_i_a3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_4_LC_5_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_4_LC_5_15_2 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst1.state_4_LC_5_15_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.state_4_LC_5_15_2  (
            .in0(_gnd_net_),
            .in1(N__22317),
            .in2(_gnd_net_),
            .in3(N__25110),
            .lcout(phase_controller_inst1_state_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50225),
            .ce(),
            .sr(N__49711));
    defparam \phase_controller_inst1.state_2_LC_5_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_2_LC_5_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_2_LC_5_16_6 .LUT_INIT=16'b1000100011111000;
    LogicCell40 \phase_controller_inst1.state_2_LC_5_16_6  (
            .in0(N__32120),
            .in1(N__22261),
            .in2(N__22629),
            .in3(N__23880),
            .lcout(\phase_controller_inst1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50216),
            .ce(),
            .sr(N__49719));
    defparam \phase_controller_inst1.state_3_LC_5_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_3_LC_5_16_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_3_LC_5_16_7 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \phase_controller_inst1.state_3_LC_5_16_7  (
            .in0(N__22260),
            .in1(N__32121),
            .in2(N__22492),
            .in3(N__22276),
            .lcout(state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50216),
            .ce(),
            .sr(N__49719));
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_5_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_5_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_5_17_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_tr_RNO_0_LC_5_17_3  (
            .in0(_gnd_net_),
            .in1(N__26041),
            .in2(_gnd_net_),
            .in3(N__22587),
            .lcout(\phase_controller_inst1.start_timer_tr_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_tr_LC_5_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_LC_5_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_tr_LC_5_18_5 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \phase_controller_inst1.start_timer_tr_LC_5_18_5  (
            .in0(N__25132),
            .in1(N__25324),
            .in2(N__22285),
            .in3(N__22272),
            .lcout(\phase_controller_inst1.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50204),
            .ce(),
            .sr(N__49733));
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_5_19_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_5_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_5_19_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.state_RNI7NN7_0_LC_5_19_1  (
            .in0(_gnd_net_),
            .in1(N__22558),
            .in2(_gnd_net_),
            .in3(N__22537),
            .lcout(\phase_controller_inst1.state_RNI7NN7Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MAX_D2_LC_7_3_7.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_7_3_7.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_7_3_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MAX_D2_LC_7_3_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22840),
            .lcout(il_max_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50275),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MIN_D1_LC_7_4_7.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MIN_D1_LC_7_4_7.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MIN_D1_LC_7_4_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MIN_D1_LC_7_4_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22222),
            .lcout(il_min_comp2_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50273),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MIN_D2_LC_7_5_1.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MIN_D2_LC_7_5_1.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MIN_D2_LC_7_5_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MIN_D2_LC_7_5_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22213),
            .lcout(il_min_comp2_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50270),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MAX_D1_LC_7_5_2.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MAX_D1_LC_7_5_2.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MAX_D1_LC_7_5_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MAX_D1_LC_7_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22396),
            .lcout(il_max_comp2_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50270),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MAX_D2_LC_7_8_1.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MAX_D2_LC_7_8_1.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MAX_D2_LC_7_8_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MAX_D2_LC_7_8_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22381),
            .lcout(il_max_comp2_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50255),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MIN_D2_LC_7_9_3.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_7_9_3.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_7_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MIN_D2_LC_7_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23815),
            .lcout(il_min_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50250),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_1_LC_7_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_1_LC_7_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_1_LC_7_10_5 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \phase_controller_inst2.state_1_LC_7_10_5  (
            .in0(N__22470),
            .in1(N__28033),
            .in2(N__22685),
            .in3(N__27999),
            .lcout(\phase_controller_inst2.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50243),
            .ce(),
            .sr(N__49669));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_7_11_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_7_11_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_7_11_2  (
            .in0(_gnd_net_),
            .in1(N__26386),
            .in2(_gnd_net_),
            .in3(N__30498),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_302_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_7_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_7_11_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.start_timer_tr_RNO_0_LC_7_11_6  (
            .in0(N__22675),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22469),
            .lcout(\phase_controller_inst2.start_timer_tr_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_tr_LC_7_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_LC_7_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_tr_LC_7_12_7 .LUT_INIT=16'b1111000011110010;
    LogicCell40 \phase_controller_inst2.start_timer_tr_LC_7_12_7  (
            .in0(N__29907),
            .in1(N__25133),
            .in2(N__22351),
            .in3(N__22342),
            .lcout(\phase_controller_inst2.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50231),
            .ce(),
            .sr(N__49683));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_7_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_7_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_7_13_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_7_13_2  (
            .in0(N__29701),
            .in1(N__29815),
            .in2(N__29959),
            .in3(N__22417),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50226),
            .ce(),
            .sr(N__49689));
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_7_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_7_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_7_14_3 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_inst2.stoper_tr.time_passed_LC_7_14_3  (
            .in0(N__22446),
            .in1(N__23035),
            .in2(N__22900),
            .in3(N__29860),
            .lcout(\phase_controller_inst2.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50217),
            .ce(),
            .sr(N__49696));
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_7_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_7_14_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.state_RNI9M3O_0_LC_7_14_5  (
            .in0(_gnd_net_),
            .in1(N__22445),
            .in2(_gnd_net_),
            .in3(N__22431),
            .lcout(\phase_controller_inst2.state_RNI9M3OZ0Z_0 ),
            .ltout(\phase_controller_inst2.state_RNI9M3OZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_3_LC_7_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_3_LC_7_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_3_LC_7_14_6 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \phase_controller_inst2.state_3_LC_7_14_6  (
            .in0(N__26095),
            .in1(N__25730),
            .in2(N__22495),
            .in3(N__22491),
            .lcout(\phase_controller_inst2.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50217),
            .ce(),
            .sr(N__49696));
    defparam \phase_controller_inst2.state_0_LC_7_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_0_LC_7_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_0_LC_7_14_7 .LUT_INIT=16'b1010111000001100;
    LogicCell40 \phase_controller_inst2.state_0_LC_7_14_7  (
            .in0(N__22471),
            .in1(N__22432),
            .in2(N__22450),
            .in3(N__22686),
            .lcout(\phase_controller_inst2.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50217),
            .ce(),
            .sr(N__49696));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_7_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_7_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(N__23050),
            .in2(N__24535),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_15_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_LC_7_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_LC_7_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_LC_7_15_1  (
            .in0(_gnd_net_),
            .in1(N__24505),
            .in2(_gnd_net_),
            .in3(N__22423),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_3_LC_7_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_3_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_3_LC_7_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_3_LC_7_15_2  (
            .in0(_gnd_net_),
            .in1(N__23041),
            .in2(N__24484),
            .in3(N__22420),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_4_LC_7_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_4_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_4_LC_7_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_4_LC_7_15_3  (
            .in0(_gnd_net_),
            .in1(N__24460),
            .in2(_gnd_net_),
            .in3(N__22408),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_5_LC_7_15_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_5_LC_7_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_5_LC_7_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_5_LC_7_15_4  (
            .in0(_gnd_net_),
            .in1(N__24850),
            .in2(_gnd_net_),
            .in3(N__22405),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_6_LC_7_15_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_6_LC_7_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_6_LC_7_15_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_6_LC_7_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24817),
            .in3(N__22402),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_7_LC_7_15_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_7_LC_7_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_7_LC_7_15_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_7_LC_7_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24793),
            .in3(N__22399),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_8_LC_7_15_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_8_LC_7_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_8_LC_7_15_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_8_LC_7_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24769),
            .in3(N__22522),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_9_LC_7_16_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_9_LC_7_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_9_LC_7_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_9_LC_7_16_0  (
            .in0(_gnd_net_),
            .in1(N__24744),
            .in2(_gnd_net_),
            .in3(N__22519),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_9 ),
            .ltout(),
            .carryin(bfn_7_16_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_10_LC_7_16_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_10_LC_7_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_10_LC_7_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_10_LC_7_16_1  (
            .in0(_gnd_net_),
            .in1(N__24724),
            .in2(_gnd_net_),
            .in3(N__22516),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_11_LC_7_16_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_11_LC_7_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_11_LC_7_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_11_LC_7_16_2  (
            .in0(_gnd_net_),
            .in1(N__24706),
            .in2(_gnd_net_),
            .in3(N__22513),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_12_LC_7_16_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_12_LC_7_16_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_12_LC_7_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_12_LC_7_16_3  (
            .in0(_gnd_net_),
            .in1(N__24688),
            .in2(_gnd_net_),
            .in3(N__22510),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_13_LC_7_16_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_13_LC_7_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_13_LC_7_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_13_LC_7_16_4  (
            .in0(_gnd_net_),
            .in1(N__24985),
            .in2(_gnd_net_),
            .in3(N__22507),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_14_LC_7_16_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_14_LC_7_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_14_LC_7_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_14_LC_7_16_5  (
            .in0(_gnd_net_),
            .in1(N__24967),
            .in2(_gnd_net_),
            .in3(N__22504),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_15_LC_7_16_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_15_LC_7_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_15_LC_7_16_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_15_LC_7_16_6  (
            .in0(_gnd_net_),
            .in1(N__24949),
            .in2(_gnd_net_),
            .in3(N__22501),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_16_LC_7_16_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_16_LC_7_16_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_16_LC_7_16_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_16_LC_7_16_7  (
            .in0(_gnd_net_),
            .in1(N__24927),
            .in2(_gnd_net_),
            .in3(N__22498),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_17_LC_7_17_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_17_LC_7_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_17_LC_7_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_17_LC_7_17_0  (
            .in0(_gnd_net_),
            .in1(N__24907),
            .in2(_gnd_net_),
            .in3(N__22639),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_17 ),
            .ltout(),
            .carryin(bfn_7_17_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_18_LC_7_17_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_18_LC_7_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_18_LC_7_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_18_LC_7_17_1  (
            .in0(_gnd_net_),
            .in1(N__24889),
            .in2(_gnd_net_),
            .in3(N__22636),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_19_LC_7_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_19_LC_7_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_19_LC_7_17_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_19_LC_7_17_2  (
            .in0(_gnd_net_),
            .in1(N__24871),
            .in2(_gnd_net_),
            .in3(N__22633),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_7_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_7_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_7_17_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_0_LC_7_17_3  (
            .in0(_gnd_net_),
            .in1(N__22630),
            .in2(_gnd_net_),
            .in3(N__23873),
            .lcout(\phase_controller_inst1.start_timer_hc_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_7_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_7_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_7_17_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_7_17_6  (
            .in0(N__25373),
            .in1(N__25633),
            .in2(_gnd_net_),
            .in3(N__25515),
            .lcout(\phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_7_17_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_7_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_7_17_7 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_7_17_7  (
            .in0(N__25516),
            .in1(_gnd_net_),
            .in2(N__25660),
            .in3(N__25374),
            .lcout(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_7_18_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_7_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_7_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_16_LC_7_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28081),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50189),
            .ce(N__25176),
            .sr(N__49720));
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_7_19_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_7_19_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_7_19_3 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_LC_7_19_3  (
            .in0(N__22557),
            .in1(N__25783),
            .in2(N__22603),
            .in3(N__25814),
            .lcout(\phase_controller_inst1.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50183),
            .ce(),
            .sr(N__49727));
    defparam \phase_controller_inst1.state_0_LC_7_19_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_0_LC_7_19_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_0_LC_7_19_5 .LUT_INIT=16'b1011001110100000;
    LogicCell40 \phase_controller_inst1.state_0_LC_7_19_5  (
            .in0(N__22580),
            .in1(N__22556),
            .in2(N__26062),
            .in3(N__22536),
            .lcout(\phase_controller_inst1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50183),
            .ce(),
            .sr(N__49727));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_7_19_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_7_19_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_7_19_6 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_7_19_6  (
            .in0(N__25658),
            .in1(N__25385),
            .in2(N__23653),
            .in3(N__25551),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50183),
            .ce(),
            .sr(N__49727));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_7_19_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_7_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_7_19_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_7_19_7  (
            .in0(N__25550),
            .in1(N__25659),
            .in2(N__25427),
            .in3(N__22645),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50183),
            .ce(),
            .sr(N__49727));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_7_20_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_7_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_7_20_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_7_20_1  (
            .in0(N__25778),
            .in1(N__23375),
            .in2(_gnd_net_),
            .in3(N__25808),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_7_20_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_7_20_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_7_20_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_7_20_2  (
            .in0(N__25652),
            .in1(N__25532),
            .in2(N__25434),
            .in3(N__23503),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50178),
            .ce(),
            .sr(N__49734));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_7_20_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_7_20_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_7_20_3 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_7_20_3  (
            .in0(N__25529),
            .in1(N__25417),
            .in2(N__23479),
            .in3(N__25655),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50178),
            .ce(),
            .sr(N__49734));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_7_20_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_7_20_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_7_20_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_7_20_4  (
            .in0(N__25653),
            .in1(N__25533),
            .in2(N__25435),
            .in3(N__23449),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50178),
            .ce(),
            .sr(N__49734));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_7_20_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_7_20_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_7_20_5 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_7_20_5  (
            .in0(N__25530),
            .in1(N__25418),
            .in2(N__23425),
            .in3(N__25656),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50178),
            .ce(),
            .sr(N__49734));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_7_20_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_7_20_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_7_20_6 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_7_20_6  (
            .in0(N__25654),
            .in1(N__25534),
            .in2(N__25436),
            .in3(N__23707),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50178),
            .ce(),
            .sr(N__49734));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_7_20_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_7_20_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_7_20_7 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_7_20_7  (
            .in0(N__25531),
            .in1(N__25419),
            .in2(N__23683),
            .in3(N__25657),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50178),
            .ce(),
            .sr(N__49734));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_7_21_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_7_21_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_7_21_0 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_7_21_0  (
            .in0(N__25509),
            .in1(N__25641),
            .in2(N__25428),
            .in3(N__23620),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50173),
            .ce(),
            .sr(N__49737));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_7_21_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_7_21_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_7_21_1 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_7_21_1  (
            .in0(N__25637),
            .in1(N__25386),
            .in2(N__25552),
            .in3(N__23596),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50173),
            .ce(),
            .sr(N__49737));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_7_21_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_7_21_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_7_21_2 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_7_21_2  (
            .in0(N__25510),
            .in1(N__25642),
            .in2(N__25429),
            .in3(N__23569),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50173),
            .ce(),
            .sr(N__49737));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_7_21_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_7_21_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_7_21_3 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_7_21_3  (
            .in0(N__25638),
            .in1(N__25387),
            .in2(N__25553),
            .in3(N__23335),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50173),
            .ce(),
            .sr(N__49737));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_7_21_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_7_21_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_7_21_4 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_7_21_4  (
            .in0(N__25511),
            .in1(N__25643),
            .in2(N__25430),
            .in3(N__23305),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50173),
            .ce(),
            .sr(N__49737));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_7_21_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_7_21_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_7_21_5 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_7_21_5  (
            .in0(N__25639),
            .in1(N__25388),
            .in2(N__25554),
            .in3(N__23278),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50173),
            .ce(),
            .sr(N__49737));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_7_21_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_7_21_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_7_21_6 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_7_21_6  (
            .in0(N__25512),
            .in1(N__25644),
            .in2(N__25431),
            .in3(N__23563),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50173),
            .ce(),
            .sr(N__49737));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_7_21_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_7_21_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_7_21_7 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_7_21_7  (
            .in0(N__25640),
            .in1(N__25389),
            .in2(N__25555),
            .in3(N__23536),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50173),
            .ce(),
            .sr(N__49737));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_0_LC_7_22_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_0_LC_7_22_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_0_LC_7_22_2 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_0_LC_7_22_2  (
            .in0(N__25815),
            .in1(N__25631),
            .in2(N__25432),
            .in3(N__25513),
            .lcout(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50167),
            .ce(N__36399),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_1_LC_7_22_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_1_LC_7_22_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_1_LC_7_22_4 .LUT_INIT=16'b0001000111000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_1_LC_7_22_4  (
            .in0(N__25816),
            .in1(N__25632),
            .in2(N__25433),
            .in3(N__25514),
            .lcout(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50167),
            .ce(N__36399),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.S2_LC_7_23_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.S2_LC_7_23_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S2_LC_7_23_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S2_LC_7_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22690),
            .lcout(s4_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50163),
            .ce(),
            .sr(N__49740));
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_3_2.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_3_2.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_3_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MAX_D1_LC_8_3_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22849),
            .lcout(il_max_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50274),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQJB4_15_LC_8_8_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQJB4_15_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQJB4_15_LC_8_8_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIQJB4_15_LC_8_8_1  (
            .in0(N__24187),
            .in1(N__24208),
            .in2(N__24169),
            .in3(N__24223),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_10_LC_8_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_10_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_10_LC_8_8_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_10_LC_8_8_5  (
            .in0(_gnd_net_),
            .in1(N__24669),
            .in2(_gnd_net_),
            .in3(N__23919),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI5IJ5_27_LC_8_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI5IJ5_27_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI5IJ5_27_LC_8_8_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI5IJ5_27_LC_8_8_6  (
            .in0(N__24324),
            .in1(N__24649),
            .in2(N__22834),
            .in3(N__24301),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_8_8_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_8_8_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_8_8_7  (
            .in0(N__22756),
            .in1(N__22831),
            .in2(N__22825),
            .in3(N__22888),
            .lcout(\current_shift_inst.PI_CTRL.N_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA3B4_11_LC_8_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA3B4_11_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA3B4_11_LC_8_9_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIA3B4_11_LC_8_9_0  (
            .in0(N__24262),
            .in1(N__24276),
            .in2(N__24238),
            .in3(N__23904),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_10_LC_8_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_10_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_10_LC_8_9_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_10_LC_8_9_1  (
            .in0(N__24277),
            .in1(N__24670),
            .in2(N__23926),
            .in3(N__24391),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_8_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_8_9_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_8_9_2  (
            .in0(N__22696),
            .in1(N__22867),
            .in2(N__22750),
            .in3(N__22861),
            .lcout(\current_shift_inst.PI_CTRL.N_118 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIKHF4_11_LC_8_9_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIKHF4_11_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIKHF4_11_LC_8_9_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIKHF4_11_LC_8_9_3  (
            .in0(N__23905),
            .in1(N__24297),
            .in2(N__24325),
            .in3(N__24645),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIBB4_13_LC_8_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIBB4_13_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIBB4_13_LC_8_9_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIIBB4_13_LC_8_9_5  (
            .in0(N__24222),
            .in1(N__24234),
            .in2(N__24207),
            .in3(N__24261),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNITR72_25_LC_8_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNITR72_25_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNITR72_25_LC_8_9_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNITR72_25_LC_8_9_6  (
            .in0(_gnd_net_),
            .in1(N__24343),
            .in2(_gnd_net_),
            .in3(N__24361),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI5VT8_23_LC_8_9_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI5VT8_23_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI5VT8_23_LC_8_9_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI5VT8_23_LC_8_9_7  (
            .in0(N__24379),
            .in1(N__24390),
            .in2(N__22891),
            .in3(N__22882),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFBE4_19_LC_8_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFBE4_19_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFBE4_19_LC_8_10_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIFBE4_19_LC_8_10_1  (
            .in0(N__24435),
            .in1(N__24147),
            .in2(N__24408),
            .in3(N__24424),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_19_LC_8_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_19_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_19_LC_8_10_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_19_LC_8_10_4  (
            .in0(N__24148),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24436),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIBVN8_17_LC_8_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIBVN8_17_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIBVN8_17_LC_8_10_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIBVN8_17_LC_8_10_5  (
            .in0(N__24186),
            .in1(N__24165),
            .in2(N__22876),
            .in3(N__22873),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVBJ5_22_LC_8_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVBJ5_22_LC_8_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVBJ5_22_LC_8_10_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIVBJ5_22_LC_8_10_7  (
            .in0(N__24342),
            .in1(N__24360),
            .in2(N__24409),
            .in3(N__22855),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINL72_21_LC_8_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINL72_21_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINL72_21_LC_8_11_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNINL72_21_LC_8_11_4  (
            .in0(_gnd_net_),
            .in1(N__24375),
            .in2(_gnd_net_),
            .in3(N__24423),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_8_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_8_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_8_12_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_11_LC_8_12_0  (
            .in0(_gnd_net_),
            .in1(N__26464),
            .in2(_gnd_net_),
            .in3(N__28186),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50227),
            .ce(N__25192),
            .sr(N__49677));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_8_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_8_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_8_13_0 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_8_13_0  (
            .in0(N__29696),
            .in1(N__29910),
            .in2(N__22966),
            .in3(N__29814),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50218),
            .ce(),
            .sr(N__49684));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_8_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_8_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_8_13_1 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_8_13_1  (
            .in0(N__29809),
            .in1(N__29698),
            .in2(N__29956),
            .in3(N__22951),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50218),
            .ce(),
            .sr(N__49684));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_8_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_8_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_8_13_2 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_8_13_2  (
            .in0(N__29694),
            .in1(N__29908),
            .in2(N__23017),
            .in3(N__29812),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50218),
            .ce(),
            .sr(N__49684));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_8_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_8_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_8_13_3 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_8_13_3  (
            .in0(N__29808),
            .in1(N__29697),
            .in2(N__29955),
            .in3(N__22942),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50218),
            .ce(),
            .sr(N__49684));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_8_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_8_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_8_13_5 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_8_13_5  (
            .in0(N__29811),
            .in1(N__29700),
            .in2(N__29958),
            .in3(N__22933),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50218),
            .ce(),
            .sr(N__49684));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_8_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_8_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_8_13_6 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_8_13_6  (
            .in0(N__29695),
            .in1(N__29909),
            .in2(N__22924),
            .in3(N__29813),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50218),
            .ce(),
            .sr(N__49684));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_8_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_8_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_8_13_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_8_13_7  (
            .in0(N__29810),
            .in1(N__29699),
            .in2(N__29957),
            .in3(N__22909),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50218),
            .ce(),
            .sr(N__49684));
    defparam \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_8_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_8_14_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_8_14_0  (
            .in0(N__29754),
            .in1(N__29927),
            .in2(_gnd_net_),
            .in3(N__29659),
            .lcout(\phase_controller_inst2.stoper_tr.time_passed_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.stoper_state_RNIH19L_0_LC_8_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.stoper_state_RNIH19L_0_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.stoper_state_RNIH19L_0_LC_8_14_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \phase_controller_inst2.stoper_tr.stoper_state_RNIH19L_0_LC_8_14_1  (
            .in0(N__29926),
            .in1(N__29658),
            .in2(_gnd_net_),
            .in3(N__29753),
            .lcout(\phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_8_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_8_14_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_8_14_4  (
            .in0(_gnd_net_),
            .in1(N__23033),
            .in2(_gnd_net_),
            .in3(N__29835),
            .lcout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.stoper_state_RNID9EC_0_LC_8_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.stoper_state_RNID9EC_0_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.stoper_state_RNID9EC_0_LC_8_14_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.stoper_state_RNID9EC_0_LC_8_14_5  (
            .in0(_gnd_net_),
            .in1(N__29657),
            .in2(_gnd_net_),
            .in3(N__29752),
            .lcout(\phase_controller_inst2.stoper_tr.time_passed11 ),
            .ltout(\phase_controller_inst2.stoper_tr.time_passed11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNIF9HJ_LC_8_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNIF9HJ_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNIF9HJ_LC_8_14_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNIF9HJ_LC_8_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23044),
            .in3(N__29836),
            .lcout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNIF9HJZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_1_LC_8_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_1_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_1_LC_8_15_1 .LUT_INIT=16'b0110110001101100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_1_LC_8_15_1  (
            .in0(N__23034),
            .in1(N__24534),
            .in2(N__29848),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_8_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_8_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_8_15_2 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_8_15_2  (
            .in0(N__29651),
            .in1(N__29981),
            .in2(N__23005),
            .in3(N__29805),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50205),
            .ce(),
            .sr(N__49697));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_8_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_8_15_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_8_15_3 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_8_15_3  (
            .in0(N__29802),
            .in1(N__29654),
            .in2(N__29991),
            .in3(N__22996),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50205),
            .ce(),
            .sr(N__49697));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_8_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_8_15_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_8_15_4 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_8_15_4  (
            .in0(N__29652),
            .in1(N__29982),
            .in2(N__22990),
            .in3(N__29806),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50205),
            .ce(),
            .sr(N__49697));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_8_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_8_15_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_8_15_5 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_8_15_5  (
            .in0(N__29803),
            .in1(N__29655),
            .in2(N__29992),
            .in3(N__22981),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50205),
            .ce(),
            .sr(N__49697));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_8_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_8_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_8_15_6 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_8_15_6  (
            .in0(N__29653),
            .in1(N__29983),
            .in2(N__22975),
            .in3(N__29807),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50205),
            .ce(),
            .sr(N__49697));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_8_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_8_15_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_8_15_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_8_15_7  (
            .in0(N__29804),
            .in1(N__29656),
            .in2(N__29993),
            .in3(N__23125),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50205),
            .ce(),
            .sr(N__49697));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_8_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_8_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_8_16_0 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_8_16_0  (
            .in0(N__29797),
            .in1(N__29963),
            .in2(N__23119),
            .in3(N__29691),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50196),
            .ce(),
            .sr(N__49702));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_8_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_8_16_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_8_16_1 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_8_16_1  (
            .in0(N__29690),
            .in1(N__29801),
            .in2(N__29990),
            .in3(N__23110),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50196),
            .ce(),
            .sr(N__49702));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_8_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_8_16_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_8_16_2 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_8_16_2  (
            .in0(N__29798),
            .in1(N__29964),
            .in2(N__23104),
            .in3(N__29692),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50196),
            .ce(),
            .sr(N__49702));
    defparam \phase_controller_inst1.start_timer_hc_LC_8_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_LC_8_16_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_hc_LC_8_16_3 .LUT_INIT=16'b1010101010111010;
    LogicCell40 \phase_controller_inst1.start_timer_hc_LC_8_16_3  (
            .in0(N__23095),
            .in1(N__25134),
            .in2(N__30989),
            .in3(N__23083),
            .lcout(\phase_controller_inst1.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50196),
            .ce(),
            .sr(N__49702));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_8_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_8_16_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_8_16_4 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_8_16_4  (
            .in0(N__29799),
            .in1(N__29965),
            .in2(N__23077),
            .in3(N__29693),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50196),
            .ce(),
            .sr(N__49702));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_8_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_8_16_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_8_16_7 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_8_16_7  (
            .in0(N__29689),
            .in1(N__29800),
            .in2(N__29989),
            .in3(N__23068),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50196),
            .ce(),
            .sr(N__49702));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_8_17_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_8_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_8_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_8_17_0  (
            .in0(_gnd_net_),
            .in1(N__23062),
            .in2(N__25066),
            .in3(N__23376),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_8_17_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_8_17_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_8_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_8_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_8_17_1  (
            .in0(_gnd_net_),
            .in1(N__23056),
            .in2(N__25027),
            .in3(N__23353),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_8_17_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_8_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_8_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_8_17_2  (
            .in0(_gnd_net_),
            .in1(N__23194),
            .in2(N__25057),
            .in3(N__23326),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_8_17_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_8_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_8_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_8_17_3  (
            .in0(_gnd_net_),
            .in1(N__23188),
            .in2(N__25219),
            .in3(N__23296),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_8_17_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_8_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_8_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_8_17_4  (
            .in0(_gnd_net_),
            .in1(N__23182),
            .in2(N__25249),
            .in3(N__23268),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_8_17_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_8_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_8_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_8_17_5  (
            .in0(_gnd_net_),
            .in1(N__23176),
            .in2(N__25231),
            .in3(N__23553),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_8_17_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_8_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_8_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_8_17_6  (
            .in0(_gnd_net_),
            .in1(N__25033),
            .in2(N__23170),
            .in3(N__25705),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_8_17_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_8_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_8_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_8_17_7  (
            .in0(_gnd_net_),
            .in1(N__23161),
            .in2(N__25264),
            .in3(N__25680),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_8_18_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_8_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_8_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_8_18_0  (
            .in0(_gnd_net_),
            .in1(N__23155),
            .in2(N__25048),
            .in3(N__25275),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_8_18_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_8_18_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_8_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_8_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_8_18_1  (
            .in0(_gnd_net_),
            .in1(N__23149),
            .in2(N__25201),
            .in3(N__23518),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_8_18_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_8_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_8_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_8_18_2  (
            .in0(_gnd_net_),
            .in1(N__23131),
            .in2(N__23143),
            .in3(N__23494),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_8_18_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_8_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_8_18_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_8_18_3  (
            .in0(N__23466),
            .in1(N__23251),
            .in2(N__25240),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_8_18_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_8_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_8_18_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_8_18_4  (
            .in0(_gnd_net_),
            .in1(N__23245),
            .in2(N__25210),
            .in3(N__23440),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_8_18_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_8_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_8_18_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_8_18_5  (
            .in0(N__23722),
            .in1(N__23239),
            .in2(N__25015),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_8_18_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_8_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_8_18_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_8_18_6  (
            .in0(N__23698),
            .in1(N__23233),
            .in2(N__25000),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_8_18_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_8_18_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_8_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_8_18_7  (
            .in0(_gnd_net_),
            .in1(N__23218),
            .in2(N__23227),
            .in3(N__23664),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_8_19_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_8_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_8_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_8_19_0  (
            .in0(_gnd_net_),
            .in1(N__23212),
            .in2(N__23404),
            .in3(N__23635),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_8_19_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_8_19_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_8_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_8_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_8_19_1  (
            .in0(_gnd_net_),
            .in1(N__23206),
            .in2(N__23395),
            .in3(N__23611),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_8_19_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_8_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_8_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_8_19_2  (
            .in0(_gnd_net_),
            .in1(N__23200),
            .in2(N__23386),
            .in3(N__23587),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_8_19_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_8_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_8_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_8_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23407),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_8_19_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_8_19_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_8_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_17_LC_8_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29461),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50179),
            .ce(N__25191),
            .sr(N__49721));
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_8_19_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_8_19_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_8_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_18_LC_8_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29418),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50179),
            .ce(N__25191),
            .sr(N__49721));
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_8_19_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_8_19_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_8_19_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_19_LC_8_19_6  (
            .in0(N__29333),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50179),
            .ce(N__25191),
            .sr(N__49721));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_8_20_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_8_20_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_8_20_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_8_20_0  (
            .in0(_gnd_net_),
            .in1(N__25822),
            .in2(N__23377),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_20_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_8_20_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_8_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_8_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_8_20_1  (
            .in0(_gnd_net_),
            .in1(N__23349),
            .in2(_gnd_net_),
            .in3(N__23329),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_8_20_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_8_20_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_8_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_8_20_2  (
            .in0(_gnd_net_),
            .in1(N__25750),
            .in2(N__23325),
            .in3(N__23299),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_8_20_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_8_20_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_8_20_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_8_20_3  (
            .in0(_gnd_net_),
            .in1(N__23292),
            .in2(_gnd_net_),
            .in3(N__23272),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_8_20_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_8_20_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_8_20_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_8_20_4  (
            .in0(_gnd_net_),
            .in1(N__23269),
            .in2(_gnd_net_),
            .in3(N__23557),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_8_20_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_8_20_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_8_20_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_8_20_5  (
            .in0(_gnd_net_),
            .in1(N__23554),
            .in2(_gnd_net_),
            .in3(N__23530),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_8_20_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_8_20_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_8_20_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_8_20_6  (
            .in0(_gnd_net_),
            .in1(N__25704),
            .in2(_gnd_net_),
            .in3(N__23527),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_8_20_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_8_20_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_8_20_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_8_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25681),
            .in3(N__23524),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_8_21_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_8_21_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_8_21_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_8_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25282),
            .in3(N__23521),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9 ),
            .ltout(),
            .carryin(bfn_8_21_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_8_21_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_8_21_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_8_21_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_8_21_1  (
            .in0(_gnd_net_),
            .in1(N__23517),
            .in2(_gnd_net_),
            .in3(N__23497),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_8_21_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_8_21_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_8_21_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_8_21_2  (
            .in0(_gnd_net_),
            .in1(N__23493),
            .in2(_gnd_net_),
            .in3(N__23470),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_8_21_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_8_21_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_8_21_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_8_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23467),
            .in3(N__23443),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_8_21_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_8_21_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_8_21_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_8_21_4  (
            .in0(_gnd_net_),
            .in1(N__23439),
            .in2(_gnd_net_),
            .in3(N__23410),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_8_21_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_8_21_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_8_21_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_8_21_5  (
            .in0(_gnd_net_),
            .in1(N__23721),
            .in2(_gnd_net_),
            .in3(N__23701),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_8_21_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_8_21_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_8_21_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_8_21_6  (
            .in0(_gnd_net_),
            .in1(N__23697),
            .in2(_gnd_net_),
            .in3(N__23671),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_8_21_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_8_21_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_8_21_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_8_21_7  (
            .in0(_gnd_net_),
            .in1(N__23668),
            .in2(_gnd_net_),
            .in3(N__23638),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_8_22_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_8_22_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_8_22_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_8_22_0  (
            .in0(_gnd_net_),
            .in1(N__23634),
            .in2(_gnd_net_),
            .in3(N__23614),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17 ),
            .ltout(),
            .carryin(bfn_8_22_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_8_22_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_8_22_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_8_22_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_8_22_1  (
            .in0(_gnd_net_),
            .in1(N__23610),
            .in2(_gnd_net_),
            .in3(N__23590),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_8_22_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_8_22_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_8_22_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_8_22_2  (
            .in0(_gnd_net_),
            .in1(N__23586),
            .in2(_gnd_net_),
            .in3(N__23572),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_8_22_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_8_22_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_8_22_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_8_22_3  (
            .in0(_gnd_net_),
            .in1(N__25587),
            .in2(_gnd_net_),
            .in3(N__25476),
            .lcout(\phase_controller_inst1.stoper_tr.time_passed11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_8_23_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_8_23_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_8_23_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_8_23_6  (
            .in0(N__30972),
            .in1(N__30896),
            .in2(_gnd_net_),
            .in3(N__30770),
            .lcout(\phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_8_24_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_8_24_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_8_24_6 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_LC_8_24_6  (
            .in0(N__23864),
            .in1(N__28831),
            .in2(N__23893),
            .in3(N__25977),
            .lcout(\phase_controller_inst1.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50155),
            .ce(),
            .sr(N__49741));
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_8_30_4.C_ON=1'b0;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_8_30_4.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_8_30_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_8_30_4 (
            .in0(N__23848),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_clk_12mhz_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.stop_timer_hc_LC_9_6_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_hc_LC_9_6_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.stop_timer_hc_LC_9_6_2 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \delay_measurement_inst.stop_timer_hc_LC_9_6_2  (
            .in0(N__27364),
            .in1(N__26179),
            .in2(N__49792),
            .in3(N__27397),
            .lcout(\delay_measurement_inst.stop_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50256),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MIN_D1_LC_9_6_5.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_9_6_5.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_9_6_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MIN_D1_LC_9_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23824),
            .lcout(il_min_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50256),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_9_7_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_9_7_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_9_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_14_LC_9_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43873),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50251),
            .ce(),
            .sr(N__49640));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_9_8_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_9_8_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_9_8_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_0_LC_9_8_0  (
            .in0(_gnd_net_),
            .in1(N__39436),
            .in2(N__26188),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ),
            .ltout(),
            .carryin(bfn_9_8_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ),
            .clk(N__50244),
            .ce(),
            .sr(N__49647));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_9_8_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_9_8_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_9_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_LC_9_8_1  (
            .in0(_gnd_net_),
            .in1(N__36530),
            .in2(N__26146),
            .in3(N__23776),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .clk(N__50244),
            .ce(),
            .sr(N__49647));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_9_8_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_9_8_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_9_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_2_LC_9_8_2  (
            .in0(_gnd_net_),
            .in1(N__26128),
            .in2(N__39403),
            .in3(N__23758),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .clk(N__50244),
            .ce(),
            .sr(N__49647));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_9_8_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_9_8_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_9_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_3_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(N__40882),
            .in2(N__28996),
            .in3(N__23725),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .clk(N__50244),
            .ce(),
            .sr(N__49647));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_9_8_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_9_8_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_9_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_4_LC_9_8_4  (
            .in0(_gnd_net_),
            .in1(N__39360),
            .in2(N__26161),
            .in3(N__24085),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .clk(N__50244),
            .ce(),
            .sr(N__49647));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_9_8_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_9_8_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_9_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_5_LC_9_8_5  (
            .in0(_gnd_net_),
            .in1(N__26152),
            .in2(N__43477),
            .in3(N__24052),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .clk(N__50244),
            .ce(),
            .sr(N__49647));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_9_8_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_9_8_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_9_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_6_LC_9_8_6  (
            .in0(_gnd_net_),
            .in1(N__43535),
            .in2(N__26137),
            .in3(N__24022),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .clk(N__50244),
            .ce(),
            .sr(N__49647));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_9_8_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_9_8_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_9_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_7_LC_9_8_7  (
            .in0(_gnd_net_),
            .in1(N__44202),
            .in2(N__28954),
            .in3(N__23992),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .clk(N__50244),
            .ce(),
            .sr(N__49647));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_9_9_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_9_9_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_9_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_8_LC_9_9_0  (
            .in0(_gnd_net_),
            .in1(N__43636),
            .in2(N__26269),
            .in3(N__23959),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ),
            .ltout(),
            .carryin(bfn_9_9_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .clk(N__50237),
            .ce(),
            .sr(N__49652));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_9_9_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_9_9_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_9_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_9_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(N__43591),
            .in2(N__26236),
            .in3(N__23929),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .clk(N__50237),
            .ce(),
            .sr(N__49652));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_9_9_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_9_9_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_9_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_10_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(N__43801),
            .in2(N__27583),
            .in3(N__23908),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .clk(N__50237),
            .ce(),
            .sr(N__49652));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_9_9_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_9_9_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_9_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_11_LC_9_9_3  (
            .in0(_gnd_net_),
            .in1(N__41739),
            .in2(N__27673),
            .in3(N__23896),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .clk(N__50237),
            .ce(),
            .sr(N__49652));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_9_9_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_9_9_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_9_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_12_LC_9_9_4  (
            .in0(_gnd_net_),
            .in1(N__41670),
            .in2(N__26257),
            .in3(N__24265),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .clk(N__50237),
            .ce(),
            .sr(N__49652));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_9_9_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_9_9_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_9_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_13_LC_9_9_5  (
            .in0(_gnd_net_),
            .in1(N__44139),
            .in2(N__26245),
            .in3(N__24253),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .clk(N__50237),
            .ce(),
            .sr(N__49652));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_9_9_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_9_9_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_9_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_14_LC_9_9_6  (
            .in0(_gnd_net_),
            .in1(N__41523),
            .in2(N__24250),
            .in3(N__24226),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .clk(N__50237),
            .ce(),
            .sr(N__49652));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_9_9_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_9_9_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_9_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_15_LC_9_9_7  (
            .in0(_gnd_net_),
            .in1(N__26122),
            .in2(N__36927),
            .in3(N__24211),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .clk(N__50237),
            .ce(),
            .sr(N__49652));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_9_10_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_9_10_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_9_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_16_LC_9_10_0  (
            .in0(_gnd_net_),
            .in1(N__37116),
            .in2(N__27514),
            .in3(N__24190),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ),
            .ltout(),
            .carryin(bfn_9_10_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .clk(N__50232),
            .ce(),
            .sr(N__49656));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_9_10_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_9_10_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_9_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_17_LC_9_10_1  (
            .in0(_gnd_net_),
            .in1(N__27604),
            .in2(N__41800),
            .in3(N__24172),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .clk(N__50232),
            .ce(),
            .sr(N__49656));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_9_10_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_9_10_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_9_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_18_LC_9_10_2  (
            .in0(_gnd_net_),
            .in1(N__40206),
            .in2(N__26116),
            .in3(N__24151),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .clk(N__50232),
            .ce(),
            .sr(N__49656));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_9_10_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_9_10_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_9_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_19_LC_9_10_3  (
            .in0(_gnd_net_),
            .in1(N__40149),
            .in2(N__27619),
            .in3(N__24139),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .clk(N__50232),
            .ce(),
            .sr(N__49656));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_9_10_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_9_10_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_9_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_20_LC_9_10_4  (
            .in0(_gnd_net_),
            .in1(N__40269),
            .in2(N__27595),
            .in3(N__24427),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .clk(N__50232),
            .ce(),
            .sr(N__49656));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_9_10_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_9_10_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_9_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_21_LC_9_10_5  (
            .in0(_gnd_net_),
            .in1(N__41458),
            .in2(N__27730),
            .in3(N__24412),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .clk(N__50232),
            .ce(),
            .sr(N__49656));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_9_10_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_9_10_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_9_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_22_LC_9_10_6  (
            .in0(_gnd_net_),
            .in1(N__39491),
            .in2(N__27526),
            .in3(N__24394),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .clk(N__50232),
            .ce(),
            .sr(N__49656));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_9_10_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_9_10_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_9_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_23_LC_9_10_7  (
            .in0(_gnd_net_),
            .in1(N__26224),
            .in2(N__44461),
            .in3(N__24382),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .clk(N__50232),
            .ce(),
            .sr(N__49656));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_9_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_9_11_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_9_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_24_LC_9_11_0  (
            .in0(_gnd_net_),
            .in1(N__44573),
            .in2(N__27742),
            .in3(N__24364),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ),
            .ltout(),
            .carryin(bfn_9_11_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .clk(N__50228),
            .ce(),
            .sr(N__49662));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_9_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_9_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_9_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_25_LC_9_11_1  (
            .in0(_gnd_net_),
            .in1(N__41344),
            .in2(N__27658),
            .in3(N__24346),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .clk(N__50228),
            .ce(),
            .sr(N__49662));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_9_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_9_11_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_9_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_26_LC_9_11_2  (
            .in0(_gnd_net_),
            .in1(N__44653),
            .in2(N__26216),
            .in3(N__24328),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .clk(N__50228),
            .ce(),
            .sr(N__49662));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_9_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_9_11_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_9_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_27_LC_9_11_3  (
            .in0(_gnd_net_),
            .in1(N__26207),
            .in2(N__36832),
            .in3(N__24304),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .clk(N__50228),
            .ce(),
            .sr(N__49662));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_9_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_9_11_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_9_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_28_LC_9_11_4  (
            .in0(_gnd_net_),
            .in1(N__44521),
            .in2(N__26217),
            .in3(N__24280),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .clk(N__50228),
            .ce(),
            .sr(N__49662));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_9_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_9_11_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_9_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_29_LC_9_11_5  (
            .in0(_gnd_net_),
            .in1(N__26211),
            .in2(N__39996),
            .in3(N__24652),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .clk(N__50228),
            .ce(),
            .sr(N__49662));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_9_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_9_11_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_9_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_30_LC_9_11_6  (
            .in0(_gnd_net_),
            .in1(N__32191),
            .in2(N__26218),
            .in3(N__24631),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ),
            .clk(N__50228),
            .ce(),
            .sr(N__49662));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_9_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_9_11_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_9_11_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_31_LC_9_11_7  (
            .in0(N__44913),
            .in1(N__26215),
            .in2(_gnd_net_),
            .in3(N__24628),
            .lcout(\current_shift_inst.PI_CTRL.un8_enablelto31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50228),
            .ce(),
            .sr(N__49662));
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_9_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_9_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_9_12_2 .LUT_INIT=16'b0101010100010001;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_6_LC_9_12_2  (
            .in0(N__26680),
            .in1(N__26759),
            .in2(_gnd_net_),
            .in3(N__27828),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50219),
            .ce(N__33917),
            .sr(N__49670));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_9_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_9_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_9_13_0  (
            .in0(_gnd_net_),
            .in1(N__24511),
            .in2(N__26311),
            .in3(N__24524),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_9_13_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_9_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_9_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_9_13_1  (
            .in0(_gnd_net_),
            .in1(N__24490),
            .in2(N__26302),
            .in3(N__24501),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_9_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_9_13_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_9_13_2  (
            .in0(N__24477),
            .in1(N__24466),
            .in2(N__26281),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_9_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_9_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_9_13_3  (
            .in0(_gnd_net_),
            .in1(N__24442),
            .in2(N__26344),
            .in3(N__24459),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_9_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_9_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_9_13_4  (
            .in0(_gnd_net_),
            .in1(N__24835),
            .in2(N__26353),
            .in3(N__24846),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_9_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_9_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_9_13_5  (
            .in0(_gnd_net_),
            .in1(N__24799),
            .in2(N__24829),
            .in3(N__24810),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_9_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_9_13_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_9_13_6  (
            .in0(_gnd_net_),
            .in1(N__24775),
            .in2(N__26323),
            .in3(N__24786),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_9_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_9_13_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_9_13_7  (
            .in0(N__24762),
            .in1(N__24751),
            .in2(N__26335),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_9_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_9_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_9_14_0  (
            .in0(_gnd_net_),
            .in1(N__24730),
            .in2(N__26530),
            .in3(N__24745),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_9_14_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_9_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_9_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(N__24712),
            .in2(N__26476),
            .in3(N__24723),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_9_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_9_14_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(N__24694),
            .in2(N__26488),
            .in3(N__24705),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_9_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_9_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(N__24676),
            .in2(N__26509),
            .in3(N__24687),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_9_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_9_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_9_14_4  (
            .in0(_gnd_net_),
            .in1(N__24973),
            .in2(N__26497),
            .in3(N__24984),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_9_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_9_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_9_14_5  (
            .in0(_gnd_net_),
            .in1(N__24955),
            .in2(N__26410),
            .in3(N__24966),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_9_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_9_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(N__24937),
            .in2(N__33943),
            .in3(N__24948),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_9_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_9_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_9_14_7  (
            .in0(_gnd_net_),
            .in1(N__24913),
            .in2(N__26293),
            .in3(N__24931),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_9_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_9_15_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_9_15_0  (
            .in0(_gnd_net_),
            .in1(N__24895),
            .in2(N__26518),
            .in3(N__24906),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_9_15_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_9_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_9_15_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_9_15_1  (
            .in0(N__24888),
            .in1(N__24877),
            .in2(N__25084),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_9_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_9_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(N__24859),
            .in2(N__25075),
            .in3(N__24870),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_9_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_9_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24853),
            .lcout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_9_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_9_15_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_9_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_18_LC_9_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29419),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50197),
            .ce(N__33925),
            .sr(N__49690));
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_9_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_9_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_9_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_19_LC_9_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29334),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50197),
            .ce(N__33925),
            .sr(N__49690));
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_9_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_9_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_9_16_0 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_1_LC_9_16_0  (
            .in0(N__26717),
            .in1(N__26639),
            .in2(N__27799),
            .in3(N__26555),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50190),
            .ce(N__25189),
            .sr(N__49698));
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_9_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_9_16_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_9_16_1 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_3_LC_9_16_1  (
            .in0(N__26638),
            .in1(N__26715),
            .in2(N__27886),
            .in3(N__26577),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50190),
            .ce(N__25189),
            .sr(N__49698));
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_9_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_9_16_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_9_16_2 .LUT_INIT=16'b1111010011110101;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_9_LC_9_16_2  (
            .in0(N__26446),
            .in1(N__34047),
            .in2(N__27919),
            .in3(N__28108),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50190),
            .ce(N__25189),
            .sr(N__49698));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_9_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_9_16_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_9_16_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_LC_9_16_3  (
            .in0(_gnd_net_),
            .in1(N__26716),
            .in2(_gnd_net_),
            .in3(N__27568),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50190),
            .ce(N__25189),
            .sr(N__49698));
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_9_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_9_16_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_9_16_4 .LUT_INIT=16'b0000000011100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_2_LC_9_16_4  (
            .in0(N__26718),
            .in1(N__26640),
            .in2(N__27856),
            .in3(N__26556),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50190),
            .ce(N__25189),
            .sr(N__49698));
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_9_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_9_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_9_16_5 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_14_LC_9_16_5  (
            .in0(N__34046),
            .in1(N__33983),
            .in2(_gnd_net_),
            .in3(N__27775),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50190),
            .ce(N__25189),
            .sr(N__49698));
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_9_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_9_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_9_16_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_15_LC_9_16_6  (
            .in0(N__33984),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34048),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50190),
            .ce(N__25189),
            .sr(N__49698));
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_9_17_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_9_17_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_9_17_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_8_LC_9_17_0  (
            .in0(N__26731),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27715),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50184),
            .ce(N__25190),
            .sr(N__49703));
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_9_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_9_17_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_9_17_2 .LUT_INIT=16'b1111101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_5_LC_9_17_2  (
            .in0(N__26729),
            .in1(_gnd_net_),
            .in2(N__26670),
            .in3(N__27646),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50184),
            .ce(N__25190),
            .sr(N__49703));
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_9_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_9_17_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_9_17_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_12_LC_9_17_3  (
            .in0(_gnd_net_),
            .in1(N__26459),
            .in2(_gnd_net_),
            .in3(N__28210),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50184),
            .ce(N__25190),
            .sr(N__49703));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_9_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_9_17_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_9_17_4 .LUT_INIT=16'b0000111100000101;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_LC_9_17_4  (
            .in0(N__26730),
            .in1(_gnd_net_),
            .in2(N__26671),
            .in3(N__27829),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50184),
            .ce(N__25190),
            .sr(N__49703));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_9_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_9_17_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_9_17_5 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_LC_9_17_5  (
            .in0(N__27949),
            .in1(N__26648),
            .in2(_gnd_net_),
            .in3(N__26728),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50184),
            .ce(N__25190),
            .sr(N__49703));
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_9_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_9_17_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_9_17_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_13_LC_9_17_6  (
            .in0(N__26460),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28162),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50184),
            .ce(N__25190),
            .sr(N__49703));
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_9_17_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_9_17_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_9_17_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_10_LC_9_17_7  (
            .in0(_gnd_net_),
            .in1(N__26458),
            .in2(_gnd_net_),
            .in3(N__28135),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50184),
            .ce(N__25190),
            .sr(N__49703));
    defparam \phase_controller_inst2.start_timer_hc_RNO_1_LC_9_18_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_RNO_1_LC_9_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_hc_RNO_1_LC_9_18_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.start_timer_hc_RNO_1_LC_9_18_0  (
            .in0(_gnd_net_),
            .in1(N__26096),
            .in2(_gnd_net_),
            .in3(N__25737),
            .lcout(),
            .ltout(\phase_controller_inst2.start_timer_hc_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_hc_LC_9_18_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_LC_9_18_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_hc_LC_9_18_1 .LUT_INIT=16'b1111000011110010;
    LogicCell40 \phase_controller_inst2.start_timer_hc_LC_9_18_1  (
            .in0(N__30260),
            .in1(N__27961),
            .in2(N__25138),
            .in3(N__25135),
            .lcout(\phase_controller_inst2.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50180),
            .ce(),
            .sr(N__49705));
    defparam \phase_controller_inst2.state_2_LC_9_18_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_2_LC_9_18_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_2_LC_9_18_3 .LUT_INIT=16'b1101010111000000;
    LogicCell40 \phase_controller_inst2.state_2_LC_9_18_3  (
            .in0(N__28000),
            .in1(N__25738),
            .in2(N__26103),
            .in3(N__28019),
            .lcout(\phase_controller_inst2.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50180),
            .ce(),
            .sr(N__49705));
    defparam \phase_controller_inst2.stoper_hc.stoper_state_RNINF2L_0_LC_9_18_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.stoper_state_RNINF2L_0_LC_9_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.stoper_state_RNINF2L_0_LC_9_18_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.stoper_state_RNINF2L_0_LC_9_18_4  (
            .in0(N__30186),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30447),
            .lcout(\phase_controller_inst2.stoper_hc.time_passed11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_9_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_9_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_9_18_6 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_9_18_6  (
            .in0(N__30187),
            .in1(N__30261),
            .in2(N__28651),
            .in3(N__30448),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50180),
            .ce(),
            .sr(N__49705));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_9_19_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_9_19_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_9_19_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_9_19_0  (
            .in0(N__25661),
            .in1(N__25548),
            .in2(N__25437),
            .in3(N__25711),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50174),
            .ce(),
            .sr(N__49712));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_9_19_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_9_19_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_9_19_1 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_9_19_1  (
            .in0(N__25547),
            .in1(N__25420),
            .in2(N__25690),
            .in3(N__25663),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50174),
            .ce(),
            .sr(N__49712));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_9_19_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_9_19_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_9_19_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_9_19_2  (
            .in0(N__25662),
            .in1(N__25549),
            .in2(N__25438),
            .in3(N__25291),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50174),
            .ce(),
            .sr(N__49712));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_9_19_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_9_19_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_9_19_5 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_9_19_5  (
            .in0(N__30184),
            .in1(N__30437),
            .in2(N__30308),
            .in3(N__26866),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50174),
            .ce(),
            .sr(N__49712));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_3_LC_9_19_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_3_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_3_LC_9_19_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_3_LC_9_19_6  (
            .in0(N__29456),
            .in1(N__29417),
            .in2(N__29335),
            .in3(N__28080),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_9_19_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_9_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_9_19_7 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_9_19_7  (
            .in0(N__30183),
            .in1(N__30436),
            .in2(N__30307),
            .in3(N__28285),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50174),
            .ce(),
            .sr(N__49712));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_0_LC_9_20_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_0_LC_9_20_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_0_LC_9_20_0 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_0_LC_9_20_0  (
            .in0(N__30843),
            .in1(N__30717),
            .in2(N__31077),
            .in3(N__25983),
            .lcout(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50168),
            .ce(N__36410),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_1_LC_9_20_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_1_LC_9_20_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_1_LC_9_20_1 .LUT_INIT=16'b0000110001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_1_LC_9_20_1  (
            .in0(N__25984),
            .in1(N__31022),
            .in2(N__30757),
            .in3(N__30844),
            .lcout(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50168),
            .ce(N__36410),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_9_20_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_9_20_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_9_20_6  (
            .in0(_gnd_net_),
            .in1(N__25774),
            .in2(_gnd_net_),
            .in3(N__25806),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_9_20_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_9_20_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_9_20_7 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_9_20_7  (
            .in0(N__25807),
            .in1(_gnd_net_),
            .in2(N__25782),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_9_21_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_9_21_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_9_21_0 .LUT_INIT=16'b1111110011111000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_1_LC_9_21_0  (
            .in0(N__30549),
            .in1(N__31748),
            .in2(N__31522),
            .in3(N__32983),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50164),
            .ce(N__31594),
            .sr(N__49728));
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_9_21_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_9_21_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_9_21_3 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_5_LC_9_21_3  (
            .in0(N__31751),
            .in1(_gnd_net_),
            .in2(N__31521),
            .in3(N__31165),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50164),
            .ce(N__31594),
            .sr(N__49728));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_9_21_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_9_21_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_9_21_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_LC_9_21_4  (
            .in0(N__32839),
            .in1(N__31750),
            .in2(_gnd_net_),
            .in3(N__31493),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50164),
            .ce(N__31594),
            .sr(N__49728));
    defparam \phase_controller_inst1.stoper_hc.target_time_0_LC_9_21_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_0_LC_9_21_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_0_LC_9_21_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_0_LC_9_21_5  (
            .in0(N__31747),
            .in1(N__30551),
            .in2(N__31520),
            .in3(N__33076),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50164),
            .ce(N__31594),
            .sr(N__49728));
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_9_21_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_9_21_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_9_21_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_2_LC_9_21_6  (
            .in0(N__30550),
            .in1(N__31749),
            .in2(N__32796),
            .in3(N__31492),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50164),
            .ce(N__31594),
            .sr(N__49728));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_9_22_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_9_22_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_9_22_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_9_22_0  (
            .in0(_gnd_net_),
            .in1(N__25744),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_22_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_9_22_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_9_22_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_9_22_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_9_22_1  (
            .in0(_gnd_net_),
            .in1(N__25897),
            .in2(N__25906),
            .in3(N__27128),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_9_22_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_9_22_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_9_22_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_9_22_2  (
            .in0(_gnd_net_),
            .in1(N__25882),
            .in2(N__25891),
            .in3(N__27114),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_9_22_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_9_22_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_9_22_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_9_22_3  (
            .in0(_gnd_net_),
            .in1(N__25876),
            .in2(N__28924),
            .in3(N__27084),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_9_22_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_9_22_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_9_22_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_9_22_4  (
            .in0(_gnd_net_),
            .in1(N__25861),
            .in2(N__25870),
            .in3(N__27063),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_9_22_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_9_22_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_9_22_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_9_22_5  (
            .in0(_gnd_net_),
            .in1(N__25846),
            .in2(N__25855),
            .in3(N__27042),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_9_22_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_9_22_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_9_22_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_9_22_6  (
            .in0(_gnd_net_),
            .in1(N__25840),
            .in2(N__28696),
            .in3(N__27021),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_9_22_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_9_22_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_9_22_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_9_22_7  (
            .in0(_gnd_net_),
            .in1(N__25834),
            .in2(N__28684),
            .in3(N__27000),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_9_23_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_9_23_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_9_23_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_9_23_0  (
            .in0(_gnd_net_),
            .in1(N__25828),
            .in2(N__28867),
            .in3(N__27342),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(bfn_9_23_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_9_23_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_9_23_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_9_23_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_9_23_1  (
            .in0(N__27318),
            .in1(N__25954),
            .in2(N__30655),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_9_23_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_9_23_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_9_23_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_9_23_2  (
            .in0(_gnd_net_),
            .in1(N__25948),
            .in2(N__28843),
            .in3(N__27291),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_9_23_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_9_23_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_9_23_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_9_23_3  (
            .in0(_gnd_net_),
            .in1(N__25942),
            .in2(N__31768),
            .in3(N__27268),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_9_23_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_9_23_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_9_23_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_9_23_4  (
            .in0(N__27244),
            .in1(N__25936),
            .in2(N__30640),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_9_23_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_9_23_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_9_23_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_9_23_5  (
            .in0(_gnd_net_),
            .in1(N__25930),
            .in2(N__28897),
            .in3(N__27220),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_9_23_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_9_23_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_9_23_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_9_23_6  (
            .in0(_gnd_net_),
            .in1(N__25924),
            .in2(N__28855),
            .in3(N__27196),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_9_23_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_9_23_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_9_23_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_9_23_7  (
            .in0(_gnd_net_),
            .in1(N__25918),
            .in2(N__28909),
            .in3(N__27172),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_9_24_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_9_24_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_9_24_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_9_24_0  (
            .in0(_gnd_net_),
            .in1(N__25912),
            .in2(N__28711),
            .in3(N__27501),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_16 ),
            .ltout(),
            .carryin(bfn_9_24_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_9_24_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_9_24_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_9_24_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_9_24_1  (
            .in0(_gnd_net_),
            .in1(N__26005),
            .in2(N__31609),
            .in3(N__27480),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_17 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_9_24_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_9_24_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_9_24_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_9_24_2  (
            .in0(_gnd_net_),
            .in1(N__25999),
            .in2(N__28939),
            .in3(N__27459),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_9_24_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_9_24_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_9_24_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_9_24_3  (
            .in0(_gnd_net_),
            .in1(N__25993),
            .in2(N__28882),
            .in3(N__27439),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_9_24_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_9_24_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_9_24_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_9_24_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25987),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_9_24_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_9_24_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_9_24_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_9_24_5  (
            .in0(N__28829),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25975),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_9_24_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_9_24_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_9_24_6 .LUT_INIT=16'b0101101011110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_9_24_6  (
            .in0(N__25976),
            .in1(_gnd_net_),
            .in2(N__27142),
            .in3(N__28830),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_9_24_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_9_24_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_9_24_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_9_24_7  (
            .in0(N__28828),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25974),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_9_25_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_9_25_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_9_25_0 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_9_25_0  (
            .in0(N__30794),
            .in1(N__30908),
            .in2(N__31104),
            .in3(N__27448),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50147),
            .ce(),
            .sr(N__49742));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_9_25_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_9_25_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_9_25_1 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_9_25_1  (
            .in0(N__30904),
            .in1(N__30798),
            .in2(N__31100),
            .in3(N__27469),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50147),
            .ce(),
            .sr(N__49742));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_9_25_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_9_25_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_9_25_2 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_9_25_2  (
            .in0(N__30792),
            .in1(N__30906),
            .in2(N__31102),
            .in3(N__27181),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50147),
            .ce(),
            .sr(N__49742));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_9_25_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_9_25_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_9_25_3 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_9_25_3  (
            .in0(N__30903),
            .in1(N__30797),
            .in2(N__31099),
            .in3(N__27490),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50147),
            .ce(),
            .sr(N__49742));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_9_25_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_9_25_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_9_25_4 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_9_25_4  (
            .in0(N__30793),
            .in1(N__30907),
            .in2(N__31103),
            .in3(N__27157),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50147),
            .ce(),
            .sr(N__49742));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_9_25_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_9_25_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_9_25_5 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_9_25_5  (
            .in0(N__30901),
            .in1(N__30795),
            .in2(N__31097),
            .in3(N__27229),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50147),
            .ce(),
            .sr(N__49742));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_9_25_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_9_25_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_9_25_6 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_9_25_6  (
            .in0(N__30791),
            .in1(N__30905),
            .in2(N__31101),
            .in3(N__27253),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50147),
            .ce(),
            .sr(N__49742));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_9_25_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_9_25_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_9_25_7 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_9_25_7  (
            .in0(N__30902),
            .in1(N__30796),
            .in2(N__31098),
            .in3(N__27205),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50147),
            .ce(),
            .sr(N__49742));
    defparam \phase_controller_inst2.S1_LC_9_26_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.S1_LC_9_26_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S1_LC_9_26_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S1_LC_9_26_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26107),
            .lcout(s3_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50142),
            .ce(),
            .sr(N__49745));
    defparam \phase_controller_inst1.S2_LC_9_26_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.S2_LC_9_26_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S2_LC_9_26_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S2_LC_9_26_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26061),
            .lcout(s2_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50142),
            .ce(),
            .sr(N__49745));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_9_26_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_9_26_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_9_26_7 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_9_26_7  (
            .in0(N__30909),
            .in1(N__30799),
            .in2(N__31094),
            .in3(N__27421),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50142),
            .ce(),
            .sr(N__49745));
    defparam \delay_measurement_inst.hc_state_0_LC_10_6_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.hc_state_0_LC_10_6_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.hc_state_0_LC_10_6_5 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \delay_measurement_inst.hc_state_0_LC_10_6_5  (
            .in0(N__27359),
            .in1(N__26177),
            .in2(_gnd_net_),
            .in3(N__27385),
            .lcout(\delay_measurement_inst.hc_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50245),
            .ce(N__36411),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_10_7_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_10_7_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_10_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_0_LC_10_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33265),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50238),
            .ce(),
            .sr(N__49628));
    defparam \delay_measurement_inst.start_timer_hc_LC_10_7_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_hc_LC_10_7_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.start_timer_hc_LC_10_7_6 .LUT_INIT=16'b1101110100100010;
    LogicCell40 \delay_measurement_inst.start_timer_hc_LC_10_7_6  (
            .in0(N__27393),
            .in1(N__27363),
            .in2(_gnd_net_),
            .in3(N__26178),
            .lcout(\delay_measurement_inst.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50238),
            .ce(),
            .sr(N__49628));
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_10_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_10_8_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_10_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_4_LC_10_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36205),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50233),
            .ce(),
            .sr(N__49636));
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_10_8_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_10_8_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_10_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_5_LC_10_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36241),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50233),
            .ce(),
            .sr(N__49636));
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_10_8_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_10_8_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_10_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_1_LC_10_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33241),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50233),
            .ce(),
            .sr(N__49636));
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_10_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_10_8_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_10_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_6_LC_10_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36277),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50233),
            .ce(),
            .sr(N__49636));
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_10_8_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_10_8_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_10_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_2_LC_10_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33451),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50233),
            .ce(),
            .sr(N__49636));
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_10_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_10_9_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_10_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_15_LC_10_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36862),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50229),
            .ce(),
            .sr(N__49641));
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_10_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_10_9_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_10_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_18_LC_10_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41572),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50229),
            .ce(),
            .sr(N__49641));
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_10_9_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_10_9_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_10_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_8_LC_10_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36169),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50229),
            .ce(),
            .sr(N__49641));
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_10_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_10_9_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_10_9_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_12_LC_10_9_5  (
            .in0(_gnd_net_),
            .in1(N__36570),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50229),
            .ce(),
            .sr(N__49641));
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_10_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_10_9_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_10_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_13_LC_10_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36321),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50229),
            .ce(),
            .sr(N__49641));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_10_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_10_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_10_10_3  (
            .in0(_gnd_net_),
            .in1(N__37064),
            .in2(_gnd_net_),
            .in3(N__44019),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_10_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_10_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_10_10_5  (
            .in0(N__37199),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44018),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_10_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_10_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_10_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_9_LC_10_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36642),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50209),
            .ce(),
            .sr(N__49653));
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_10_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_10_11_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_10_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_23_LC_10_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36739),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50209),
            .ce(),
            .sr(N__49653));
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_10_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_10_11_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_10_11_4 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_LC_10_11_4  (
            .in0(N__26401),
            .in1(N__26385),
            .in2(_gnd_net_),
            .in3(N__30497),
            .lcout(\delay_measurement_inst.delay_hc_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50209),
            .ce(),
            .sr(N__49653));
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_10_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_10_11_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_10_11_5 .LUT_INIT=16'b0011000011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_30_LC_10_11_5  (
            .in0(N__45117),
            .in1(N__45279),
            .in2(N__44917),
            .in3(N__40012),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50209),
            .ce(),
            .sr(N__49653));
    defparam \current_shift_inst.PI_CTRL.prop_term_26_LC_10_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_26_LC_10_11_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_26_LC_10_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_26_LC_10_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44078),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50209),
            .ce(),
            .sr(N__49653));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_10_12_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_10_12_0 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_10_12_0  (
            .in0(N__26400),
            .in1(N__26384),
            .in2(_gnd_net_),
            .in3(N__30496),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_303_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_10_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_10_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_10_13_0 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_5_LC_10_13_0  (
            .in0(N__26750),
            .in1(N__26674),
            .in2(_gnd_net_),
            .in3(N__27635),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50199),
            .ce(N__33928),
            .sr(N__49663));
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_10_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_10_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_10_13_1 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_4_LC_10_13_1  (
            .in0(N__26673),
            .in1(N__27941),
            .in2(_gnd_net_),
            .in3(N__26749),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50199),
            .ce(N__33928),
            .sr(N__49663));
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_10_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_10_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_10_13_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_8_LC_10_13_2  (
            .in0(N__26754),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27706),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50199),
            .ce(N__33928),
            .sr(N__49663));
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_10_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_10_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_10_13_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_7_LC_10_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26760),
            .in3(N__27566),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50199),
            .ce(N__33928),
            .sr(N__49663));
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_10_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_10_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_10_13_5 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_1_LC_10_13_5  (
            .in0(N__26675),
            .in1(N__26755),
            .in2(N__27792),
            .in3(N__26562),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50199),
            .ce(N__33928),
            .sr(N__49663));
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_10_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_10_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_10_13_6 .LUT_INIT=16'b0100010001000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_2_LC_10_13_6  (
            .in0(N__26563),
            .in1(N__27848),
            .in2(N__26761),
            .in3(N__26676),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50199),
            .ce(N__33928),
            .sr(N__49663));
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_10_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_10_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_10_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_16_LC_10_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28067),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50191),
            .ce(N__33921),
            .sr(N__49671));
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_10_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_10_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_10_14_1 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_3_LC_10_14_1  (
            .in0(N__26672),
            .in1(N__26732),
            .in2(N__27881),
            .in3(N__26581),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50191),
            .ce(N__33921),
            .sr(N__49671));
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_10_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_10_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_10_14_2 .LUT_INIT=16'b1100111011001111;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_9_LC_10_14_2  (
            .in0(N__34025),
            .in1(N__27908),
            .in2(N__26457),
            .in3(N__28101),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50191),
            .ce(N__33921),
            .sr(N__49671));
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_10_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_10_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_10_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_17_LC_10_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29457),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50191),
            .ce(N__33921),
            .sr(N__49671));
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_10_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_10_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_10_14_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_12_LC_10_14_4  (
            .in0(N__26441),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28203),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50191),
            .ce(N__33921),
            .sr(N__49671));
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_10_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_10_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_10_14_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_13_LC_10_14_5  (
            .in0(_gnd_net_),
            .in1(N__26442),
            .in2(_gnd_net_),
            .in3(N__28154),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50191),
            .ce(N__33921),
            .sr(N__49671));
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_10_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_10_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_10_14_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_11_LC_10_14_6  (
            .in0(N__26440),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28179),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50191),
            .ce(N__33921),
            .sr(N__49671));
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_10_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_10_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_10_14_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_10_LC_10_14_7  (
            .in0(_gnd_net_),
            .in1(N__26439),
            .in2(_gnd_net_),
            .in3(N__28127),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50191),
            .ce(N__33921),
            .sr(N__49671));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_9_LC_10_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_9_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_9_LC_10_15_1 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_9_LC_10_15_1  (
            .in0(N__33966),
            .in1(N__34021),
            .in2(_gnd_net_),
            .in3(N__27765),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_10_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_10_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_10_15_6 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_14_LC_10_15_6  (
            .in0(N__27766),
            .in1(N__34026),
            .in2(_gnd_net_),
            .in3(N__33967),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50185),
            .ce(N__33926),
            .sr(N__49678));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4_3_LC_10_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4_3_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4_3_LC_10_16_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4_3_LC_10_16_0  (
            .in0(N__27770),
            .in1(N__27642),
            .in2(N__34043),
            .in3(N__27948),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_9_LC_10_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_9_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_9_LC_10_16_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_9_LC_10_16_1  (
            .in0(_gnd_net_),
            .in1(N__28099),
            .in2(_gnd_net_),
            .in3(N__27915),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_6_LC_10_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_6_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_6_LC_10_16_2 .LUT_INIT=16'b1111111100110001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_6_LC_10_16_2  (
            .in0(N__27771),
            .in1(N__34045),
            .in2(N__26764),
            .in3(N__33968),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1_6_LC_10_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1_6_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1_6_LC_10_16_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1_6_LC_10_16_3  (
            .in0(N__27821),
            .in1(N__27711),
            .in2(_gnd_net_),
            .in3(N__27562),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0_6_LC_10_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0_6_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0_6_LC_10_16_4 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0_6_LC_10_16_4  (
            .in0(N__28100),
            .in1(_gnd_net_),
            .in2(N__26683),
            .in3(N__34044),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_LC_10_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_LC_10_16_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_LC_10_16_5  (
            .in0(N__26614),
            .in1(N__26602),
            .in2(N__26596),
            .in3(N__26587),
            .lcout(\phase_controller_inst1.stoper_tr.N_248 ),
            .ltout(\phase_controller_inst1.stoper_tr.N_248_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a3_1_LC_10_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a3_1_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a3_1_LC_10_16_6 .LUT_INIT=16'b0101000011110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a3_1_LC_10_16_6  (
            .in0(N__27849),
            .in1(_gnd_net_),
            .in2(N__26566),
            .in3(N__27882),
            .lcout(\phase_controller_inst1.stoper_tr.N_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_c_LC_10_17_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_c_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_c_LC_10_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_c_LC_10_17_0  (
            .in0(_gnd_net_),
            .in1(N__26929),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_17_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_10_17_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_10_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_10_17_1  (
            .in0(_gnd_net_),
            .in1(N__26542),
            .in2(N__28768),
            .in3(N__28260),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_10_17_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_10_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_10_17_2  (
            .in0(_gnd_net_),
            .in1(N__26536),
            .in2(N__28738),
            .in3(N__28236),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_10_17_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_10_17_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_10_17_3  (
            .in0(N__28461),
            .in1(N__26812),
            .in2(N__28753),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_10_17_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_10_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_10_17_4  (
            .in0(_gnd_net_),
            .in1(N__26806),
            .in2(N__29587),
            .in3(N__28440),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_10_17_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_10_17_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_10_17_5  (
            .in0(N__28416),
            .in1(N__26800),
            .in2(N__26905),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_10_17_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_10_17_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_10_17_6  (
            .in0(N__28395),
            .in1(N__26794),
            .in2(N__26956),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_10_17_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_10_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_10_17_7  (
            .in0(_gnd_net_),
            .in1(N__26788),
            .in2(N__26890),
            .in3(N__28371),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_10_18_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_10_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_10_18_0  (
            .in0(_gnd_net_),
            .in1(N__26782),
            .in2(N__29548),
            .in3(N__28350),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(bfn_10_18_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_10_18_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_10_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_10_18_1  (
            .in0(_gnd_net_),
            .in1(N__26776),
            .in2(N__29536),
            .in3(N__28323),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_10_18_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_10_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_10_18_2  (
            .in0(_gnd_net_),
            .in1(N__26770),
            .in2(N__30463),
            .in3(N__28296),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_10_18_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_10_18_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_10_18_3  (
            .in0(_gnd_net_),
            .in1(N__26860),
            .in2(N__30628),
            .in3(N__28662),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_10_18_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_10_18_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_10_18_4  (
            .in0(N__28633),
            .in1(N__26854),
            .in2(N__29512),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_10_18_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_10_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_10_18_5  (
            .in0(_gnd_net_),
            .in1(N__26848),
            .in2(N__26980),
            .in3(N__28609),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_10_18_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_10_18_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_10_18_6  (
            .in0(N__28582),
            .in1(N__26842),
            .in2(N__26917),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_10_18_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_10_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_10_18_7  (
            .in0(_gnd_net_),
            .in1(N__26836),
            .in2(N__29524),
            .in3(N__28558),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_10_19_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_10_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_10_19_0  (
            .in0(_gnd_net_),
            .in1(N__26830),
            .in2(N__28723),
            .in3(N__28530),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_16 ),
            .ltout(),
            .carryin(bfn_10_19_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_10_19_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_10_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_10_19_1  (
            .in0(_gnd_net_),
            .in1(N__26824),
            .in2(N__29572),
            .in3(N__28509),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_17 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_10_19_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_10_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_10_19_2  (
            .in0(_gnd_net_),
            .in1(N__26818),
            .in2(N__26941),
            .in3(N__28485),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_10_19_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_10_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_10_19_3  (
            .in0(_gnd_net_),
            .in1(N__26875),
            .in2(N__28780),
            .in3(N__28806),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_10_19_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_10_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_10_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26869),
            .lcout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_10_19_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_10_19_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_10_19_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_10_19_5  (
            .in0(_gnd_net_),
            .in1(N__30061),
            .in2(_gnd_net_),
            .in3(N__30019),
            .lcout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_LC_10_19_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_LC_10_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_LC_10_19_6 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_LC_10_19_6  (
            .in0(N__30020),
            .in1(N__30065),
            .in2(_gnd_net_),
            .in3(N__28259),
            .lcout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.stoper_state_RNI0RST_0_LC_10_19_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.stoper_state_RNI0RST_0_LC_10_19_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.stoper_state_RNI0RST_0_LC_10_19_7 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.stoper_state_RNI0RST_0_LC_10_19_7  (
            .in0(N__30239),
            .in1(N__30148),
            .in2(_gnd_net_),
            .in3(N__30435),
            .lcout(\phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_10_20_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_10_20_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_10_20_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_10_20_0  (
            .in0(N__30188),
            .in1(N__30443),
            .in2(N__30323),
            .in3(N__28618),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50161),
            .ce(),
            .sr(N__49706));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_10_20_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_10_20_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_10_20_1 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_10_20_1  (
            .in0(N__30439),
            .in1(N__30291),
            .in2(N__28594),
            .in3(N__30192),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50161),
            .ce(),
            .sr(N__49706));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_10_20_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_10_20_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_10_20_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_10_20_2  (
            .in0(N__30189),
            .in1(N__30444),
            .in2(N__30324),
            .in3(N__28567),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50161),
            .ce(),
            .sr(N__49706));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_10_20_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_10_20_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_10_20_3 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_10_20_3  (
            .in0(N__30440),
            .in1(N__30292),
            .in2(N__28543),
            .in3(N__30193),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50161),
            .ce(),
            .sr(N__49706));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_10_20_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_10_20_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_10_20_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_10_20_4  (
            .in0(N__30190),
            .in1(N__30445),
            .in2(N__30325),
            .in3(N__28519),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50161),
            .ce(),
            .sr(N__49706));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_10_20_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_10_20_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_10_20_5 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_10_20_5  (
            .in0(N__30441),
            .in1(N__30293),
            .in2(N__28498),
            .in3(N__30194),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50161),
            .ce(),
            .sr(N__49706));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_10_20_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_10_20_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_10_20_6 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_10_20_6  (
            .in0(N__30191),
            .in1(N__30446),
            .in2(N__30326),
            .in3(N__28474),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50161),
            .ce(),
            .sr(N__49706));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_10_20_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_10_20_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_10_20_7 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_10_20_7  (
            .in0(N__30442),
            .in1(N__30294),
            .in2(N__28792),
            .in3(N__30195),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50161),
            .ce(),
            .sr(N__49706));
    defparam \phase_controller_inst2.stoper_hc.target_timeZ0Z_6_LC_10_21_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_timeZ0Z_6_LC_10_21_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_timeZ0Z_6_LC_10_21_0 .LUT_INIT=16'b0100010001010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_timeZ0Z_6_LC_10_21_0  (
            .in0(N__31497),
            .in1(N__31903),
            .in2(_gnd_net_),
            .in3(N__31740),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ1Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50157),
            .ce(N__30595),
            .sr(N__49713));
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_10_21_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_10_21_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_10_21_1 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_18_LC_10_21_1  (
            .in0(N__31744),
            .in1(N__31501),
            .in2(_gnd_net_),
            .in3(N__31246),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50157),
            .ce(N__30595),
            .sr(N__49713));
    defparam \phase_controller_inst2.stoper_hc.target_time_0_LC_10_21_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_0_LC_10_21_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_0_LC_10_21_2 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_0_LC_10_21_2  (
            .in0(N__30552),
            .in1(N__31741),
            .in2(N__31523),
            .in3(N__33075),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50157),
            .ce(N__30595),
            .sr(N__49713));
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_10_21_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_10_21_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_10_21_3 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_14_LC_10_21_3  (
            .in0(N__31743),
            .in1(N__31500),
            .in2(_gnd_net_),
            .in3(N__31957),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50157),
            .ce(N__30595),
            .sr(N__49713));
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_10_21_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_10_21_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_10_21_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_5_LC_10_21_5  (
            .in0(N__31745),
            .in1(N__31502),
            .in2(_gnd_net_),
            .in3(N__31164),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50157),
            .ce(N__30595),
            .sr(N__49713));
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_10_21_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_10_21_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_10_21_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_7_LC_10_21_6  (
            .in0(N__31498),
            .in1(N__32673),
            .in2(_gnd_net_),
            .in3(N__31746),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50157),
            .ce(N__30595),
            .sr(N__49713));
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_10_21_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_10_21_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_10_21_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_13_LC_10_21_7  (
            .in0(N__31742),
            .in1(N__31499),
            .in2(_gnd_net_),
            .in3(N__31852),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50157),
            .ce(N__30595),
            .sr(N__49713));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_10_22_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_10_22_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_10_22_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_10_22_0  (
            .in0(N__30893),
            .in1(N__30768),
            .in2(N__31096),
            .in3(N__27307),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50152),
            .ce(),
            .sr(N__49722));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_10_22_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_10_22_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_10_22_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_10_22_2  (
            .in0(N__30892),
            .in1(N__30767),
            .in2(N__31095),
            .in3(N__26968),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50152),
            .ce(),
            .sr(N__49722));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_10_23_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_10_23_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_10_23_0 .LUT_INIT=16'b1100100010001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_10_23_0  (
            .in0(N__30759),
            .in1(N__27103),
            .in2(N__30925),
            .in3(N__31093),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50148),
            .ce(),
            .sr(N__49729));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_10_23_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_10_23_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_10_23_1 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_10_23_1  (
            .in0(N__30899),
            .in1(N__30765),
            .in2(N__31107),
            .in3(N__27052),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50148),
            .ce(),
            .sr(N__49729));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_10_23_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_10_23_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_10_23_2 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_10_23_2  (
            .in0(N__30762),
            .in1(N__31080),
            .in2(N__30924),
            .in3(N__27331),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50148),
            .ce(),
            .sr(N__49729));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_10_23_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_10_23_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_10_23_3 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_10_23_3  (
            .in0(N__30897),
            .in1(N__30763),
            .in2(N__31105),
            .in3(N__27280),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50148),
            .ce(),
            .sr(N__49729));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_10_23_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_10_23_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_10_23_4 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_10_23_4  (
            .in0(N__30761),
            .in1(N__31079),
            .in2(N__30923),
            .in3(N__26989),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50148),
            .ce(),
            .sr(N__49729));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_10_23_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_10_23_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_10_23_5 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_10_23_5  (
            .in0(N__30900),
            .in1(N__30766),
            .in2(N__31108),
            .in3(N__27010),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50148),
            .ce(),
            .sr(N__49729));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_10_23_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_10_23_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_10_23_6 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_10_23_6  (
            .in0(N__30760),
            .in1(N__31078),
            .in2(N__30922),
            .in3(N__27031),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50148),
            .ce(),
            .sr(N__49729));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_10_23_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_10_23_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_10_23_7 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_10_23_7  (
            .in0(N__30898),
            .in1(N__30764),
            .in2(N__31106),
            .in3(N__27073),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50148),
            .ce(),
            .sr(N__49729));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_10_24_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_10_24_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_10_24_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_10_24_0  (
            .in0(_gnd_net_),
            .in1(N__27148),
            .in2(N__27141),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_24_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_10_24_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_10_24_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_10_24_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_10_24_1  (
            .in0(_gnd_net_),
            .in1(N__27115),
            .in2(_gnd_net_),
            .in3(N__27097),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_10_24_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_10_24_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_10_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_10_24_2  (
            .in0(_gnd_net_),
            .in1(N__27094),
            .in2(N__27088),
            .in3(N__27067),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_10_24_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_10_24_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_10_24_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_10_24_3  (
            .in0(_gnd_net_),
            .in1(N__27064),
            .in2(_gnd_net_),
            .in3(N__27046),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_10_24_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_10_24_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_10_24_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_10_24_4  (
            .in0(_gnd_net_),
            .in1(N__27043),
            .in2(_gnd_net_),
            .in3(N__27025),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_10_24_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_10_24_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_10_24_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_10_24_5  (
            .in0(_gnd_net_),
            .in1(N__27022),
            .in2(_gnd_net_),
            .in3(N__27004),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_10_24_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_10_24_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_10_24_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_10_24_6  (
            .in0(_gnd_net_),
            .in1(N__27001),
            .in2(_gnd_net_),
            .in3(N__26983),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_10_24_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_10_24_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_10_24_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_10_24_7  (
            .in0(_gnd_net_),
            .in1(N__27343),
            .in2(_gnd_net_),
            .in3(N__27325),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_10_25_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_10_25_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_10_25_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_10_25_0  (
            .in0(_gnd_net_),
            .in1(N__27322),
            .in2(_gnd_net_),
            .in3(N__27298),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_10_25_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_10_25_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_10_25_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_10_25_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_10_25_1  (
            .in0(_gnd_net_),
            .in1(N__27295),
            .in2(_gnd_net_),
            .in3(N__27271),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_10_25_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_10_25_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_10_25_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_10_25_2  (
            .in0(_gnd_net_),
            .in1(N__27267),
            .in2(_gnd_net_),
            .in3(N__27247),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_10_25_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_10_25_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_10_25_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_10_25_3  (
            .in0(_gnd_net_),
            .in1(N__27243),
            .in2(_gnd_net_),
            .in3(N__27223),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_10_25_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_10_25_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_10_25_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_10_25_4  (
            .in0(_gnd_net_),
            .in1(N__27219),
            .in2(_gnd_net_),
            .in3(N__27199),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_10_25_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_10_25_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_10_25_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_10_25_5  (
            .in0(_gnd_net_),
            .in1(N__27195),
            .in2(_gnd_net_),
            .in3(N__27175),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_10_25_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_10_25_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_10_25_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_10_25_6  (
            .in0(_gnd_net_),
            .in1(N__27171),
            .in2(_gnd_net_),
            .in3(N__27151),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_10_25_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_10_25_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_10_25_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_10_25_7  (
            .in0(_gnd_net_),
            .in1(N__27502),
            .in2(_gnd_net_),
            .in3(N__27484),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_10_26_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_10_26_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_10_26_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_10_26_0  (
            .in0(_gnd_net_),
            .in1(N__27481),
            .in2(_gnd_net_),
            .in3(N__27463),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(bfn_10_26_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_10_26_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_10_26_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_10_26_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_10_26_1  (
            .in0(_gnd_net_),
            .in1(N__27460),
            .in2(_gnd_net_),
            .in3(N__27442),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_10_26_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_10_26_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_10_26_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_10_26_2  (
            .in0(_gnd_net_),
            .in1(N__27438),
            .in2(_gnd_net_),
            .in3(N__27424),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam reset_ibuf_gb_io_RNI79U7_LC_10_28_5.C_ON=1'b0;
    defparam reset_ibuf_gb_io_RNI79U7_LC_10_28_5.SEQ_MODE=4'b0000;
    defparam reset_ibuf_gb_io_RNI79U7_LC_10_28_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 reset_ibuf_gb_io_RNI79U7_LC_10_28_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49787),
            .lcout(red_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_DELAY_HC2_LC_11_5_3.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_HC2_LC_11_5_3.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_HC2_LC_11_5_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_DELAY_HC2_LC_11_5_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27403),
            .lcout(delay_hc_d2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50246),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_DELAY_HC1_LC_11_5_4.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_HC1_LC_11_5_4.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_HC1_LC_11_5_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_DELAY_HC1_LC_11_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27415),
            .lcout(delay_hc_d1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50246),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.prev_hc_sig_LC_11_6_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.prev_hc_sig_LC_11_6_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.prev_hc_sig_LC_11_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.prev_hc_sig_LC_11_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27392),
            .lcout(\delay_measurement_inst.prev_hc_sigZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50239),
            .ce(),
            .sr(N__49621));
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_11_7_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_11_7_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_11_7_5 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_LC_11_7_5  (
            .in0(N__45067),
            .in1(N__45211),
            .in2(_gnd_net_),
            .in3(N__39241),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50234),
            .ce(),
            .sr(N__49623));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_11_8_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_11_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33766),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIIOJ3_19_LC_11_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIIOJ3_19_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIIOJ3_19_LC_11_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIIOJ3_19_LC_11_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36950),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_11_9_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_11_9_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_11_9_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_19_LC_11_9_3  (
            .in0(N__36951),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50221),
            .ce(),
            .sr(N__49637));
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_11_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_11_10_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_11_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_17_LC_11_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44266),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50210),
            .ce(),
            .sr(N__49642));
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_11_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_11_10_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_11_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_20_LC_11_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37147),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50210),
            .ce(),
            .sr(N__49642));
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_11_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_11_10_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_11_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_10_LC_11_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36610),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50210),
            .ce(),
            .sr(N__49642));
    defparam \delay_measurement_inst.delay_tr_reg_7_LC_11_10_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_7_LC_11_10_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_7_LC_11_10_3 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_7_LC_11_10_3  (
            .in0(N__29248),
            .in1(N__29028),
            .in2(N__27567),
            .in3(N__37432),
            .lcout(measured_delay_tr_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50210),
            .ce(),
            .sr(N__49642));
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_11_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_11_10_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_11_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_22_LC_11_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36451),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50210),
            .ce(),
            .sr(N__49642));
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_11_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_11_10_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_11_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_16_LC_11_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36772),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50210),
            .ce(),
            .sr(N__49642));
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_11_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_11_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_11_10_7 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_LC_11_10_7  (
            .in0(N__27988),
            .in1(N__30076),
            .in2(N__28045),
            .in3(N__30040),
            .lcout(\phase_controller_inst2.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50210),
            .ce(),
            .sr(N__49642));
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_11_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_11_11_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_11_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_24_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40330),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50206),
            .ce(),
            .sr(N__49648));
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_11_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_11_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_11_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_21_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41842),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50206),
            .ce(),
            .sr(N__49648));
    defparam \delay_measurement_inst.delay_tr_reg_8_LC_11_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_8_LC_11_11_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_8_LC_11_11_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_8_LC_11_11_4  (
            .in0(N__37404),
            .in1(N__29029),
            .in2(N__27710),
            .in3(N__29247),
            .lcout(measured_delay_tr_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50206),
            .ce(),
            .sr(N__49648));
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_11_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_11_11_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_11_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_11_LC_11_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36487),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50206),
            .ce(),
            .sr(N__49648));
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_11_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_11_11_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_11_11_6 .LUT_INIT=16'b0011000011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_29_LC_11_11_6  (
            .in0(N__45116),
            .in1(N__45280),
            .in2(N__44916),
            .in3(N__40039),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50206),
            .ce(),
            .sr(N__49648));
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_11_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_11_11_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_11_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_25_LC_11_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41392),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50206),
            .ce(),
            .sr(N__49648));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_30_LC_11_12_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_30_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_30_LC_11_12_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_30_LC_11_12_0  (
            .in0(N__29470),
            .in1(N__44344),
            .in2(N__37756),
            .in3(N__33688),
            .lcout(\delay_measurement_inst.N_325 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_esr_5_LC_11_12_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_5_LC_11_12_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_5_LC_11_12_2 .LUT_INIT=16'b1100010011000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_5_LC_11_12_2  (
            .in0(N__37486),
            .in1(N__36973),
            .in2(N__29054),
            .in3(N__29215),
            .lcout(measured_delay_tr_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50200),
            .ce(N__29288),
            .sr(N__49654));
    defparam \delay_measurement_inst.delay_tr_reg_esr_4_LC_11_12_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_4_LC_11_12_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_4_LC_11_12_6 .LUT_INIT=16'b1100010011000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_4_LC_11_12_6  (
            .in0(N__37485),
            .in1(N__36994),
            .in2(N__29053),
            .in3(N__29214),
            .lcout(measured_delay_tr_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50200),
            .ce(N__29288),
            .sr(N__49654));
    defparam \delay_measurement_inst.delay_tr_reg_esr_9_LC_11_13_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_9_LC_11_13_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_9_LC_11_13_0 .LUT_INIT=16'b0000111100000010;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_9_LC_11_13_0  (
            .in0(N__29496),
            .in1(N__37927),
            .in2(N__29107),
            .in3(N__37371),
            .lcout(measured_delay_tr_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50192),
            .ce(N__29287),
            .sr(N__49660));
    defparam \delay_measurement_inst.delay_tr_reg_esr_10_LC_11_13_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_10_LC_11_13_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_10_LC_11_13_3 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_10_LC_11_13_3  (
            .in0(N__37926),
            .in1(N__29497),
            .in2(_gnd_net_),
            .in3(N__37327),
            .lcout(measured_delay_tr_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50192),
            .ce(N__29287),
            .sr(N__49660));
    defparam \delay_measurement_inst.delay_tr_reg_ess_3_LC_11_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_ess_3_LC_11_13_4 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_tr_reg_ess_3_LC_11_13_4 .LUT_INIT=16'b1111000000100000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_ess_3_LC_11_13_4  (
            .in0(N__29213),
            .in1(N__37483),
            .in2(N__37039),
            .in3(N__29052),
            .lcout(measured_delay_tr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50192),
            .ce(N__29287),
            .sr(N__49660));
    defparam \delay_measurement_inst.delay_tr_reg_esr_2_LC_11_13_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_2_LC_11_13_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_2_LC_11_13_5 .LUT_INIT=16'b1100010011000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_2_LC_11_13_5  (
            .in0(N__37481),
            .in1(N__44311),
            .in2(N__29055),
            .in3(N__29210),
            .lcout(measured_delay_tr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50192),
            .ce(N__29287),
            .sr(N__49660));
    defparam \delay_measurement_inst.delay_tr_reg_esr_6_LC_11_13_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_6_LC_11_13_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_6_LC_11_13_6 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_6_LC_11_13_6  (
            .in0(N__29211),
            .in1(N__29051),
            .in2(_gnd_net_),
            .in3(N__37484),
            .lcout(measured_delay_tr_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50192),
            .ce(N__29287),
            .sr(N__49660));
    defparam \delay_measurement_inst.delay_tr_reg_ess_1_LC_11_13_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_ess_1_LC_11_13_7 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_tr_reg_ess_1_LC_11_13_7 .LUT_INIT=16'b1100010011000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_ess_1_LC_11_13_7  (
            .in0(N__37482),
            .in1(N__50305),
            .in2(N__29056),
            .in3(N__29212),
            .lcout(measured_delay_tr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50192),
            .ce(N__29287),
            .sr(N__49660));
    defparam \delay_measurement_inst.delay_tr_reg_esr_13_LC_11_14_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_13_LC_11_14_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_13_LC_11_14_0 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_13_LC_11_14_0  (
            .in0(N__29487),
            .in1(N__37910),
            .in2(_gnd_net_),
            .in3(N__37258),
            .lcout(measured_delay_tr_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50186),
            .ce(N__29289),
            .sr(N__49664));
    defparam \delay_measurement_inst.delay_tr_reg_esr_15_LC_11_14_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_15_LC_11_14_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_15_LC_11_14_1 .LUT_INIT=16'b1111010000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_15_LC_11_14_1  (
            .in0(N__29375),
            .in1(N__29166),
            .in2(N__37931),
            .in3(N__37693),
            .lcout(measured_delay_tr_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50186),
            .ce(N__29289),
            .sr(N__49664));
    defparam \delay_measurement_inst.delay_tr_reg_esr_14_LC_11_14_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_14_LC_11_14_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_14_LC_11_14_2 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_14_LC_11_14_2  (
            .in0(N__29488),
            .in1(N__37911),
            .in2(_gnd_net_),
            .in3(N__37738),
            .lcout(measured_delay_tr_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50186),
            .ce(N__29289),
            .sr(N__49664));
    defparam \delay_measurement_inst.delay_tr_reg_esr_16_LC_11_14_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_16_LC_11_14_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_16_LC_11_14_4 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_16_LC_11_14_4  (
            .in0(N__37651),
            .in1(N__37912),
            .in2(_gnd_net_),
            .in3(N__29374),
            .lcout(measured_delay_tr_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50186),
            .ce(N__29289),
            .sr(N__49664));
    defparam \delay_measurement_inst.delay_tr_reg_esr_11_LC_11_14_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_11_LC_11_14_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_11_LC_11_14_5 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_11_LC_11_14_5  (
            .in0(N__37908),
            .in1(N__29489),
            .in2(_gnd_net_),
            .in3(N__37303),
            .lcout(measured_delay_tr_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50186),
            .ce(N__29289),
            .sr(N__49664));
    defparam \delay_measurement_inst.delay_tr_reg_esr_12_LC_11_14_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_12_LC_11_14_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_12_LC_11_14_7 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_12_LC_11_14_7  (
            .in0(N__37909),
            .in1(N__29490),
            .in2(_gnd_net_),
            .in3(N__37282),
            .lcout(measured_delay_tr_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50186),
            .ce(N__29289),
            .sr(N__49664));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_6_LC_11_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_6_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_6_LC_11_15_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_6_LC_11_15_0  (
            .in0(N__28202),
            .in1(N__28178),
            .in2(N__28158),
            .in3(N__28131),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_11_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_11_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34444),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_o2_15_LC_11_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_o2_15_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_o2_15_LC_11_15_6 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_i_o2_15_LC_11_15_6  (
            .in0(N__29407),
            .in1(N__29443),
            .in2(N__29329),
            .in3(N__28066),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_11_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_11_16_5 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_11_16_5  (
            .in0(N__30166),
            .in1(N__30309),
            .in2(_gnd_net_),
            .in3(N__30438),
            .lcout(\phase_controller_inst2.stoper_hc.time_passed_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_11_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_11_16_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_11_16_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.start_timer_hc_RNO_0_LC_11_16_7  (
            .in0(_gnd_net_),
            .in1(N__28029),
            .in2(_gnd_net_),
            .in3(N__27989),
            .lcout(\phase_controller_inst2.start_timer_hc_RNO_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_11_17_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_11_17_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_11_17_0 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_11_17_0  (
            .in0(N__30315),
            .in1(N__30182),
            .in2(N__28225),
            .in3(N__30429),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50170),
            .ce(),
            .sr(N__49685));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_11_17_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_11_17_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_11_17_1 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_11_17_1  (
            .in0(N__30422),
            .in1(N__30319),
            .in2(N__30196),
            .in3(N__28450),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50170),
            .ce(),
            .sr(N__49685));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_11_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_11_17_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_11_17_2 .LUT_INIT=16'b1110000011010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_11_17_2  (
            .in0(N__30316),
            .in1(N__30426),
            .in2(N__28429),
            .in3(N__30179),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50170),
            .ce(),
            .sr(N__49685));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_11_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_11_17_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_11_17_3 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_11_17_3  (
            .in0(N__30423),
            .in1(N__30320),
            .in2(N__30197),
            .in3(N__28405),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50170),
            .ce(),
            .sr(N__49685));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_11_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_11_17_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_11_17_4 .LUT_INIT=16'b1110000011010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_11_17_4  (
            .in0(N__30317),
            .in1(N__30427),
            .in2(N__28384),
            .in3(N__30180),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50170),
            .ce(),
            .sr(N__49685));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_11_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_11_17_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_11_17_5 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_11_17_5  (
            .in0(N__30424),
            .in1(N__30321),
            .in2(N__30198),
            .in3(N__28360),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50170),
            .ce(),
            .sr(N__49685));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_11_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_11_17_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_11_17_6 .LUT_INIT=16'b1110000011010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_11_17_6  (
            .in0(N__30318),
            .in1(N__30428),
            .in2(N__28339),
            .in3(N__30181),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50170),
            .ce(),
            .sr(N__49685));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_11_17_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_11_17_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_11_17_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_11_17_7  (
            .in0(N__30425),
            .in1(N__30322),
            .in2(N__30199),
            .in3(N__28312),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50170),
            .ce(),
            .sr(N__49685));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_11_18_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_11_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_11_18_0  (
            .in0(_gnd_net_),
            .in1(N__28273),
            .in2(N__28267),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_18_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_2_LC_11_18_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_2_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_2_LC_11_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_2_LC_11_18_1  (
            .in0(_gnd_net_),
            .in1(N__28237),
            .in2(_gnd_net_),
            .in3(N__28213),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_3_LC_11_18_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_3_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_3_LC_11_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_3_LC_11_18_2  (
            .in0(_gnd_net_),
            .in1(N__30001),
            .in2(N__28465),
            .in3(N__28444),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_4_LC_11_18_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_4_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_4_LC_11_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_4_LC_11_18_3  (
            .in0(_gnd_net_),
            .in1(N__28441),
            .in2(_gnd_net_),
            .in3(N__28420),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_5_LC_11_18_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_5_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_5_LC_11_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_5_LC_11_18_4  (
            .in0(_gnd_net_),
            .in1(N__28417),
            .in2(_gnd_net_),
            .in3(N__28399),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_6_LC_11_18_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_6_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_6_LC_11_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_6_LC_11_18_5  (
            .in0(_gnd_net_),
            .in1(N__28396),
            .in2(_gnd_net_),
            .in3(N__28375),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_7_LC_11_18_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_7_LC_11_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_7_LC_11_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_7_LC_11_18_6  (
            .in0(_gnd_net_),
            .in1(N__28372),
            .in2(_gnd_net_),
            .in3(N__28354),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_8_LC_11_18_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_8_LC_11_18_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_8_LC_11_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_8_LC_11_18_7  (
            .in0(_gnd_net_),
            .in1(N__28351),
            .in2(_gnd_net_),
            .in3(N__28330),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_9_LC_11_19_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_9_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_9_LC_11_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_9_LC_11_19_0  (
            .in0(_gnd_net_),
            .in1(N__28327),
            .in2(_gnd_net_),
            .in3(N__28303),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_9 ),
            .ltout(),
            .carryin(bfn_11_19_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_10_LC_11_19_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_10_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_10_LC_11_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_10_LC_11_19_1  (
            .in0(_gnd_net_),
            .in1(N__28300),
            .in2(_gnd_net_),
            .in3(N__28276),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_11_LC_11_19_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_11_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_11_LC_11_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_11_LC_11_19_2  (
            .in0(_gnd_net_),
            .in1(N__28669),
            .in2(_gnd_net_),
            .in3(N__28636),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_12_LC_11_19_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_12_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_12_LC_11_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_12_LC_11_19_3  (
            .in0(_gnd_net_),
            .in1(N__28632),
            .in2(_gnd_net_),
            .in3(N__28612),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_13_LC_11_19_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_13_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_13_LC_11_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_13_LC_11_19_4  (
            .in0(_gnd_net_),
            .in1(N__28608),
            .in2(_gnd_net_),
            .in3(N__28585),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_14_LC_11_19_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_14_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_14_LC_11_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_14_LC_11_19_5  (
            .in0(_gnd_net_),
            .in1(N__28581),
            .in2(_gnd_net_),
            .in3(N__28561),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_15_LC_11_19_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_15_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_15_LC_11_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_15_LC_11_19_6  (
            .in0(_gnd_net_),
            .in1(N__28557),
            .in2(_gnd_net_),
            .in3(N__28534),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_16_LC_11_19_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_16_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_16_LC_11_19_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_16_LC_11_19_7  (
            .in0(_gnd_net_),
            .in1(N__28531),
            .in2(_gnd_net_),
            .in3(N__28513),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_17_LC_11_20_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_17_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_17_LC_11_20_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_17_LC_11_20_0  (
            .in0(_gnd_net_),
            .in1(N__28510),
            .in2(_gnd_net_),
            .in3(N__28489),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_17 ),
            .ltout(),
            .carryin(bfn_11_20_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_18_LC_11_20_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_18_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_18_LC_11_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_18_LC_11_20_1  (
            .in0(_gnd_net_),
            .in1(N__28486),
            .in2(_gnd_net_),
            .in3(N__28468),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_19_LC_11_20_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_19_LC_11_20_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_19_LC_11_20_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_19_LC_11_20_2  (
            .in0(_gnd_net_),
            .in1(N__28807),
            .in2(_gnd_net_),
            .in3(N__28795),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_11_21_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_11_21_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_11_21_0 .LUT_INIT=16'b0001000100110011;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_19_LC_11_21_0  (
            .in0(N__38779),
            .in1(N__31512),
            .in2(_gnd_net_),
            .in3(N__32731),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50153),
            .ce(N__30612),
            .sr(N__49707));
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_11_21_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_11_21_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_11_21_1 .LUT_INIT=16'b1111111011110000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_1_LC_11_21_1  (
            .in0(N__30543),
            .in1(N__32982),
            .in2(N__31524),
            .in3(N__31666),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50153),
            .ce(N__30612),
            .sr(N__49707));
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_11_21_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_11_21_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_11_21_3 .LUT_INIT=16'b1111111011110000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_3_LC_11_21_3  (
            .in0(N__30544),
            .in1(N__31327),
            .in2(N__31525),
            .in3(N__31668),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50153),
            .ce(N__30612),
            .sr(N__49707));
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_11_21_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_11_21_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_11_21_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_2_LC_11_21_4  (
            .in0(N__31667),
            .in1(N__31513),
            .in2(N__32797),
            .in3(N__30545),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50153),
            .ce(N__30612),
            .sr(N__49707));
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_11_21_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_11_21_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_11_21_5 .LUT_INIT=16'b0100010001010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_16_LC_11_21_5  (
            .in0(N__31511),
            .in1(N__33026),
            .in2(_gnd_net_),
            .in3(N__31665),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50153),
            .ce(N__30612),
            .sr(N__49707));
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_11_22_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_11_22_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_11_22_0 .LUT_INIT=16'b0100010001010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_16_LC_11_22_0  (
            .in0(N__31507),
            .in1(N__33027),
            .in2(_gnd_net_),
            .in3(N__31716),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50149),
            .ce(N__31582),
            .sr(N__49714));
    defparam \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_11_22_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_11_22_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_11_22_2 .LUT_INIT=16'b0100010001010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_11_22_2  (
            .in0(N__31506),
            .in1(N__31897),
            .in2(_gnd_net_),
            .in3(N__31715),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ1Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50149),
            .ce(N__31582),
            .sr(N__49714));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_11_22_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_11_22_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_11_22_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_LC_11_22_3  (
            .in0(N__31719),
            .in1(N__31510),
            .in2(_gnd_net_),
            .in3(N__32674),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50149),
            .ce(N__31582),
            .sr(N__49714));
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_11_22_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_11_22_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_11_22_6 .LUT_INIT=16'b0100010001010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_18_LC_11_22_6  (
            .in0(N__31508),
            .in1(N__31244),
            .in2(_gnd_net_),
            .in3(N__31717),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50149),
            .ce(N__31582),
            .sr(N__49714));
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_11_22_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_11_22_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_11_22_7 .LUT_INIT=16'b1110111011101100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_3_LC_11_22_7  (
            .in0(N__31718),
            .in1(N__31509),
            .in2(N__30553),
            .in3(N__31325),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50149),
            .ce(N__31582),
            .sr(N__49714));
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_11_23_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_11_23_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_11_23_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_15_LC_11_23_0  (
            .in0(N__31738),
            .in1(N__31395),
            .in2(_gnd_net_),
            .in3(N__32893),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50143),
            .ce(N__31584),
            .sr(N__49723));
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_11_23_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_11_23_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_11_23_1 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_13_LC_11_23_1  (
            .in0(N__31851),
            .in1(_gnd_net_),
            .in2(N__31440),
            .in3(N__31736),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50143),
            .ce(N__31584),
            .sr(N__49723));
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_11_23_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_11_23_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_11_23_2 .LUT_INIT=16'b0001000100110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_19_LC_11_23_2  (
            .in0(N__38778),
            .in1(N__31394),
            .in2(_gnd_net_),
            .in3(N__32730),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50143),
            .ce(N__31584),
            .sr(N__49723));
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_11_23_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_11_23_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_11_23_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_8_LC_11_23_4  (
            .in0(N__31739),
            .in1(N__31396),
            .in2(_gnd_net_),
            .in3(N__32947),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50143),
            .ce(N__31584),
            .sr(N__49723));
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_11_23_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_11_23_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_11_23_6 .LUT_INIT=16'b0000000011110101;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_14_LC_11_23_6  (
            .in0(N__31737),
            .in1(_gnd_net_),
            .in2(N__31953),
            .in3(N__31400),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50143),
            .ce(N__31584),
            .sr(N__49723));
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_11_23_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_11_23_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_11_23_7 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_10_LC_11_23_7  (
            .in0(N__31393),
            .in1(N__31551),
            .in2(_gnd_net_),
            .in3(N__31735),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50143),
            .ce(N__31584),
            .sr(N__49723));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_11_24_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_11_24_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_11_24_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_11_24_6  (
            .in0(_gnd_net_),
            .in1(N__30758),
            .in2(_gnd_net_),
            .in3(N__30894),
            .lcout(\phase_controller_inst1.stoper_hc.time_passed11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_26_LC_11_28_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_26_LC_11_28_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_26_LC_11_28_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_26_LC_11_28_3  (
            .in0(N__31782),
            .in1(N__41213),
            .in2(_gnd_net_),
            .in3(N__41046),
            .lcout(measured_delay_hc_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50129),
            .ce(),
            .sr(N__49743));
    defparam \phase_controller_inst1.S1_LC_11_29_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.S1_LC_11_29_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S1_LC_11_29_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S1_LC_11_29_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32155),
            .lcout(s1_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50128),
            .ce(),
            .sr(N__49746));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_12_6_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_12_6_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_12_6_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_12_6_1  (
            .in0(N__44201),
            .in1(N__43527),
            .in2(N__43589),
            .in3(N__43470),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_12_6_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_12_6_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_12_6_2 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_12_6_2  (
            .in0(N__43632),
            .in1(N__39343),
            .in2(N__28978),
            .in3(N__40877),
            .lcout(\current_shift_inst.PI_CTRL.N_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFI5U3_10_LC_12_7_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFI5U3_10_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFI5U3_10_LC_12_7_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIFI5U3_10_LC_12_7_1  (
            .in0(N__43797),
            .in1(N__40205),
            .in2(N__32059),
            .in3(N__28975),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGGAM_28_LC_12_7_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGGAM_28_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGGAM_28_LC_12_7_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIGGAM_28_LC_12_7_2  (
            .in0(N__44652),
            .in1(N__41339),
            .in2(N__44520),
            .in3(N__41446),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNINKHC1_30_LC_12_7_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNINKHC1_30_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNINKHC1_30_LC_12_7_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNINKHC1_30_LC_12_7_5  (
            .in0(N__36820),
            .in1(N__29071),
            .in2(N__32212),
            .in3(N__29080),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_10_LC_12_7_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_10_LC_12_7_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_10_LC_12_7_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI24CN6_10_LC_12_7_6  (
            .in0(N__29140),
            .in1(N__28969),
            .in2(N__28963),
            .in3(N__28960),
            .lcout(\current_shift_inst.PI_CTRL.N_74 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_12_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_12_8_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_12_8_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_7_LC_12_8_0  (
            .in0(N__36678),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50220),
            .ce(),
            .sr(N__49624));
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_12_8_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_12_8_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_12_8_2 .LUT_INIT=16'b0000000110101111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_6_LC_12_8_2  (
            .in0(N__45237),
            .in1(N__45064),
            .in2(N__44922),
            .in3(N__39562),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50220),
            .ce(),
            .sr(N__49624));
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_12_8_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_12_8_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_12_8_3 .LUT_INIT=16'b0011000011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_13_LC_12_8_3  (
            .in0(N__45060),
            .in1(N__45238),
            .in2(N__44918),
            .in3(N__39784),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50220),
            .ce(),
            .sr(N__49624));
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_12_8_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_12_8_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_12_8_4 .LUT_INIT=16'b0101000011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_14_LC_12_8_4  (
            .in0(N__45235),
            .in1(N__45062),
            .in2(N__44920),
            .in3(N__39769),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50220),
            .ce(),
            .sr(N__49624));
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_12_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_12_8_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_12_8_5 .LUT_INIT=16'b0011000011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_15_LC_12_8_5  (
            .in0(N__45061),
            .in1(N__45239),
            .in2(N__44919),
            .in3(N__39736),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50220),
            .ce(),
            .sr(N__49624));
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_12_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_12_8_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_12_8_6 .LUT_INIT=16'b0101000011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_16_LC_12_8_6  (
            .in0(N__45236),
            .in1(N__45063),
            .in2(N__44921),
            .in3(N__39706),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50220),
            .ce(),
            .sr(N__49624));
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_12_8_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_12_8_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_12_8_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_3_LC_12_8_7  (
            .in0(N__33421),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50220),
            .ce(),
            .sr(N__49624));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI758M_30_LC_12_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI758M_30_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI758M_30_LC_12_9_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI758M_30_LC_12_9_1  (
            .in0(N__41515),
            .in1(N__37099),
            .in2(N__32211),
            .in3(N__44119),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI637M_0_11_LC_12_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI637M_0_11_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI637M_0_11_LC_12_9_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI637M_0_11_LC_12_9_2  (
            .in0(N__41799),
            .in1(N__36907),
            .in2(N__41740),
            .in3(N__40259),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIKFFC1_21_LC_12_9_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIKFFC1_21_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIKFFC1_21_LC_12_9_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIKFFC1_21_LC_12_9_3  (
            .in0(N__39478),
            .in1(N__41454),
            .in2(N__28984),
            .in3(N__29002),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNID8UD2_28_LC_12_9_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID8UD2_28_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID8UD2_28_LC_12_9_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNID8UD2_28_LC_12_9_4  (
            .in0(N__44513),
            .in1(N__29062),
            .in2(N__28981),
            .in3(N__41663),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIC35V7_28_LC_12_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIC35V7_28_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIC35V7_28_LC_12_9_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIC35V7_28_LC_12_9_5  (
            .in0(N__32047),
            .in1(N__29146),
            .in2(N__29089),
            .in3(N__29086),
            .lcout(\current_shift_inst.PI_CTRL.N_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI203B_12_LC_12_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI203B_12_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI203B_12_LC_12_9_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI203B_12_LC_12_9_6  (
            .in0(_gnd_net_),
            .in1(N__41514),
            .in2(_gnd_net_),
            .in3(N__41662),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFD8M_29_LC_12_9_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFD8M_29_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFD8M_29_LC_12_9_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIFD8M_29_LC_12_9_7  (
            .in0(N__44454),
            .in1(N__37098),
            .in2(N__44126),
            .in3(N__39985),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIIIAM_24_LC_12_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIIIAM_24_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIIIAM_24_LC_12_10_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIIIAM_24_LC_12_10_0  (
            .in0(N__41340),
            .in1(N__44650),
            .in2(N__36819),
            .in3(N__44562),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_12_10_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_12_10_2 .LUT_INIT=16'b1111000011111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_12_10_2  (
            .in0(N__29170),
            .in1(N__29116),
            .in2(N__37936),
            .in3(N__29383),
            .lcout(\delay_measurement_inst.N_267 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7GAF_1_LC_12_10_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7GAF_1_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7GAF_1_LC_12_10_3 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7GAF_1_LC_12_10_3  (
            .in0(N__37369),
            .in1(N__37474),
            .in2(N__50304),
            .in3(N__37035),
            .lcout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDB3B_18_LC_12_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDB3B_18_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDB3B_18_LC_12_10_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIDB3B_18_LC_12_10_4  (
            .in0(_gnd_net_),
            .in1(N__40141),
            .in2(_gnd_net_),
            .in3(N__40195),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_12_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_12_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_12_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36911),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_12_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_12_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_12_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34135),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI99AM_29_LC_12_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI99AM_29_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI99AM_29_LC_12_10_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI99AM_29_LC_12_10_7  (
            .in0(N__44443),
            .in1(N__43789),
            .in2(N__44884),
            .in3(N__39989),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIDKK3_23_LC_12_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIDKK3_23_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIDKK3_23_LC_12_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIDKK3_23_LC_12_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36725),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_19_LC_12_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_19_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_19_LC_12_11_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICCAM_19_LC_12_11_3  (
            .in0(N__40142),
            .in1(N__44867),
            .in2(N__39493),
            .in3(N__44563),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_12_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_12_11_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_12_11_5 .LUT_INIT=16'b0011000011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_24_LC_12_11_5  (
            .in0(N__45065),
            .in1(N__45222),
            .in2(N__44914),
            .in3(N__39835),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50198),
            .ce(),
            .sr(N__49643));
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_12_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_12_11_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_12_11_7 .LUT_INIT=16'b0011001111110010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_27_LC_12_11_7  (
            .in0(N__45066),
            .in1(N__40054),
            .in2(N__44915),
            .in3(N__45223),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50198),
            .ce(),
            .sr(N__49643));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_12_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_12_12_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_12_12_1  (
            .in0(_gnd_net_),
            .in1(N__36972),
            .in2(_gnd_net_),
            .in3(N__36993),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_287_4 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_287_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRN391_2_LC_12_12_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRN391_2_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRN391_2_LC_12_12_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRN391_2_LC_12_12_2  (
            .in0(N__44303),
            .in1(N__29128),
            .in2(N__29119),
            .in3(N__37731),
            .lcout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_12_12_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_12_12_3 .LUT_INIT=16'b0001001100010001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_12_12_3  (
            .in0(N__37732),
            .in1(N__37695),
            .in2(N__37381),
            .in3(N__29097),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_290 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_esr_RNO_0_9_LC_12_12_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_RNO_0_9_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_RNO_0_9_LC_12_12_4 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_RNO_0_9_LC_12_12_4  (
            .in0(N__29098),
            .in1(N__37380),
            .in2(N__37699),
            .in3(N__29358),
            .lcout(\delay_measurement_inst.N_59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_12_12_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_12_12_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_12_12_5  (
            .in0(N__37278),
            .in1(N__37299),
            .in2(N__37257),
            .in3(N__37323),
            .lcout(\delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10 ),
            .ltout(\delay_measurement_inst.elapsed_time_ns_1_RNIUG5P1_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6_7_LC_12_12_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6_7_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6_7_LC_12_12_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6_7_LC_12_12_6  (
            .in0(N__37405),
            .in1(N__37431),
            .in2(N__29260),
            .in3(N__29357),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CKPA_31_LC_12_13_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CKPA_31_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CKPA_31_LC_12_13_0 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CKPA_31_LC_12_13_0  (
            .in0(N__29230),
            .in1(N__29176),
            .in2(N__37935),
            .in3(N__29224),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_2_LC_12_13_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_2_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_2_LC_12_13_1 .LUT_INIT=16'b0000101100001111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_2_LC_12_13_1  (
            .in0(N__29162),
            .in1(N__29257),
            .in2(N__29251),
            .in3(N__29209),
            .lcout(\delay_measurement_inst.un3_elapsed_time_tr_0_i ),
            .ltout(\delay_measurement_inst.un3_elapsed_time_tr_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_2_LC_12_13_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_2_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_2_LC_12_13_2 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_2_LC_12_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29233),
            .in3(N__49786),
            .lcout(\delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC841_9_LC_12_13_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC841_9_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC841_9_LC_12_13_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC841_9_LC_12_13_3  (
            .in0(N__37370),
            .in1(N__37736),
            .in2(N__37694),
            .in3(N__37480),
            .lcout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAPC7_15_LC_12_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAPC7_15_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAPC7_15_LC_12_13_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAPC7_15_LC_12_13_4  (
            .in0(_gnd_net_),
            .in1(N__37686),
            .in2(_gnd_net_),
            .in3(N__29223),
            .lcout(\delay_measurement_inst.N_299 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_12_13_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_12_13_6 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_12_13_6  (
            .in0(N__37571),
            .in1(N__37031),
            .in2(N__37532),
            .in3(N__44310),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIOKG82_16_LC_12_13_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIOKG82_16_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIOKG82_16_LC_12_13_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIOKG82_16_LC_12_13_7  (
            .in0(N__37610),
            .in1(N__37646),
            .in2(N__29185),
            .in3(N__29182),
            .lcout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_12_14_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_12_14_0 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_12_14_0  (
            .in0(N__37647),
            .in1(N__37533),
            .in2(N__37615),
            .in3(N__37572),
            .lcout(\delay_measurement_inst.N_265 ),
            .ltout(\delay_measurement_inst.N_265_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_12_14_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_12_14_1 .LUT_INIT=16'b1111111100001110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_12_14_1  (
            .in0(N__37692),
            .in1(N__37737),
            .in2(N__29500),
            .in3(N__29373),
            .lcout(\delay_measurement_inst.N_270 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVALS_28_LC_12_14_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVALS_28_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVALS_28_LC_12_14_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVALS_28_LC_12_14_7  (
            .in0(N__37768),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37780),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_12_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_12_15_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_12_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_12_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48856),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_fast_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50175),
            .ce(N__48264),
            .sr(N__49665));
    defparam \delay_measurement_inst.delay_tr_reg_esr_17_LC_12_16_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_17_LC_12_16_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_17_LC_12_16_1 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_17_LC_12_16_1  (
            .in0(N__37932),
            .in1(N__37614),
            .in2(_gnd_net_),
            .in3(N__29384),
            .lcout(measured_delay_tr_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50169),
            .ce(N__29296),
            .sr(N__49672));
    defparam \delay_measurement_inst.delay_tr_reg_esr_18_LC_12_16_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_18_LC_12_16_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_18_LC_12_16_2 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_18_LC_12_16_2  (
            .in0(N__29385),
            .in1(N__37933),
            .in2(_gnd_net_),
            .in3(N__37573),
            .lcout(measured_delay_tr_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50169),
            .ce(N__29296),
            .sr(N__49672));
    defparam \delay_measurement_inst.delay_tr_reg_esr_19_LC_12_16_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_19_LC_12_16_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_19_LC_12_16_3 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_19_LC_12_16_3  (
            .in0(N__37934),
            .in1(N__37534),
            .in2(_gnd_net_),
            .in3(N__29386),
            .lcout(measured_delay_tr_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50169),
            .ce(N__29296),
            .sr(N__49672));
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_12_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_12_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_12_16_7 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_inv_LC_12_16_7  (
            .in0(N__38288),
            .in1(N__29266),
            .in2(_gnd_net_),
            .in3(N__45364),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_12_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_12_17_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_12_17_0  (
            .in0(N__46528),
            .in1(N__47755),
            .in2(N__46019),
            .in3(N__42970),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_12_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_12_17_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_12_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_12_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48852),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50165),
            .ce(N__48261),
            .sr(N__49679));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_12_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_12_17_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_12_17_3  (
            .in0(N__46531),
            .in1(N__47517),
            .in2(N__46168),
            .in3(N__47145),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_12_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_12_17_4 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_12_17_4  (
            .in0(N__47146),
            .in1(N__45921),
            .in2(N__47521),
            .in3(N__46529),
            .lcout(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_12_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_12_17_5 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_12_17_5  (
            .in0(N__46530),
            .in1(N__29557),
            .in2(_gnd_net_),
            .in3(N__47314),
            .lcout(\current_shift_inst.un38_control_input_cry_0_s0_sf ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_12_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_12_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_12_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_12_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45397),
            .lcout(\current_shift_inst.un4_control_input1_1 ),
            .ltout(\current_shift_inst.un4_control_input1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_12_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_12_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_12_17_7 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_12_17_7  (
            .in0(_gnd_net_),
            .in1(N__46527),
            .in2(N__29551),
            .in3(N__47313),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_12_18_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_12_18_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_12_18_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_8_LC_12_18_1  (
            .in0(N__31479),
            .in1(N__32946),
            .in2(_gnd_net_),
            .in3(N__31755),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50160),
            .ce(N__30613),
            .sr(N__49686));
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_12_18_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_12_18_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_12_18_2 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_9_LC_12_18_2  (
            .in0(N__31756),
            .in1(N__31482),
            .in2(_gnd_net_),
            .in3(N__32001),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50160),
            .ce(N__30613),
            .sr(N__49686));
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_12_18_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_12_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_12_18_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_15_LC_12_18_4  (
            .in0(N__31754),
            .in1(N__31481),
            .in2(_gnd_net_),
            .in3(N__32892),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50160),
            .ce(N__30613),
            .sr(N__49686));
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_12_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_12_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_12_18_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_12_LC_12_18_6  (
            .in0(N__31753),
            .in1(N__31480),
            .in2(_gnd_net_),
            .in3(N__31281),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50160),
            .ce(N__30613),
            .sr(N__49686));
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_12_18_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_12_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_12_18_7 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_10_LC_12_18_7  (
            .in0(N__31478),
            .in1(N__31560),
            .in2(_gnd_net_),
            .in3(N__31752),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50160),
            .ce(N__30613),
            .sr(N__49686));
    defparam \phase_controller_inst2.stoper_hc.stoper_state_0_LC_12_19_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.stoper_state_0_LC_12_19_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.stoper_state_0_LC_12_19_0 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \phase_controller_inst2.stoper_hc.stoper_state_0_LC_12_19_0  (
            .in0(N__30032),
            .in1(N__30139),
            .in2(N__30331),
            .in3(N__30390),
            .lcout(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50156),
            .ce(N__36409),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.stoper_state_1_LC_12_19_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.stoper_state_1_LC_12_19_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.stoper_state_1_LC_12_19_1 .LUT_INIT=16'b0100000001001010;
    LogicCell40 \phase_controller_inst2.stoper_hc.stoper_state_1_LC_12_19_1  (
            .in0(N__30389),
            .in1(N__30327),
            .in2(N__30185),
            .in3(N__30033),
            .lcout(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50156),
            .ce(N__36409),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIUO2P_LC_12_19_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIUO2P_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIUO2P_LC_12_19_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIUO2P_LC_12_19_3  (
            .in0(_gnd_net_),
            .in1(N__30075),
            .in2(_gnd_net_),
            .in3(N__30031),
            .lcout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIUO2PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.stoper_state_0_LC_12_19_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.stoper_state_0_LC_12_19_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.stoper_state_0_LC_12_19_4 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.stoper_state_0_LC_12_19_4  (
            .in0(N__29611),
            .in1(N__29995),
            .in2(N__29733),
            .in3(N__29859),
            .lcout(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50156),
            .ce(N__36409),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.stoper_state_1_LC_12_19_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.stoper_state_1_LC_12_19_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.stoper_state_1_LC_12_19_5 .LUT_INIT=16'b0000101000110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.stoper_state_1_LC_12_19_5  (
            .in0(N__29994),
            .in1(N__29858),
            .in2(N__29734),
            .in3(N__29612),
            .lcout(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50156),
            .ce(N__36409),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_12_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_12_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_12_19_6  (
            .in0(N__37992),
            .in1(N__38287),
            .in2(_gnd_net_),
            .in3(N__37845),
            .lcout(\current_shift_inst.un38_control_input_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_12_20_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_12_20_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_12_20_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_4_LC_12_20_1  (
            .in0(N__31484),
            .in1(N__32835),
            .in2(_gnd_net_),
            .in3(N__31664),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50151),
            .ce(N__30611),
            .sr(N__49699));
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_12_20_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_12_20_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_12_20_4 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_17_LC_12_20_4  (
            .in0(N__31663),
            .in1(N__31485),
            .in2(_gnd_net_),
            .in3(N__31204),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50151),
            .ce(N__30611),
            .sr(N__49699));
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_12_20_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_12_20_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_12_20_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_11_LC_12_20_5  (
            .in0(N__31483),
            .in1(N__32037),
            .in2(_gnd_net_),
            .in3(N__31662),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50151),
            .ce(N__30611),
            .sr(N__49699));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto5_3_LC_12_21_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto5_3_LC_12_21_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto5_3_LC_12_21_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto5_3_LC_12_21_0  (
            .in0(N__32834),
            .in1(N__31318),
            .in2(N__31163),
            .in3(N__33068),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto5Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_12_21_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_12_21_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_12_21_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_12_21_1  (
            .in0(N__31240),
            .in1(N__31202),
            .in2(N__33139),
            .in3(N__33025),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_LC_12_21_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_LC_12_21_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_LC_12_21_2 .LUT_INIT=16'b0000101000101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto30_LC_12_21_2  (
            .in0(N__32701),
            .in1(N__31120),
            .in2(N__30562),
            .in3(N__32891),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlt31_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_12_21_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_12_21_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_12_21_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_12_21_4  (
            .in0(N__32890),
            .in1(N__31941),
            .in2(N__33028),
            .in3(N__31850),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_11_LC_12_21_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_11_LC_12_21_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_11_LC_12_21_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_11_LC_12_21_5  (
            .in0(N__31239),
            .in1(N__31203),
            .in2(N__30559),
            .in3(N__30682),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_LC_12_21_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_LC_12_21_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_LC_12_21_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_LC_12_21_6  (
            .in0(N__32717),
            .in1(N__30661),
            .in2(N__30556),
            .in3(N__38777),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlt31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_12_21_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_12_21_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_12_21_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_12_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30508),
            .lcout(\delay_measurement_inst.delay_hc_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto8_LC_12_22_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto8_LC_12_22_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto8_LC_12_22_0 .LUT_INIT=16'b1000110000001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto8_LC_12_22_0  (
            .in0(N__32742),
            .in1(N__30681),
            .in2(N__31901),
            .in3(N__30469),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un1_startlt9_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto14_LC_12_22_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto14_LC_12_22_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto14_LC_12_22_1 .LUT_INIT=16'b0000100010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto14_LC_12_22_1  (
            .in0(N__31952),
            .in1(N__32000),
            .in2(N__31123),
            .in3(N__31114),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlt15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto13_1_LC_12_22_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto13_1_LC_12_22_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto13_1_LC_12_22_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto13_1_LC_12_22_2  (
            .in0(N__31278),
            .in1(N__31558),
            .in2(N__31849),
            .in3(N__32034),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto13Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_12_22_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_12_22_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_12_22_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_12_22_3  (
            .in0(N__31026),
            .in1(N__30895),
            .in2(_gnd_net_),
            .in3(N__30769),
            .lcout(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_9_LC_12_22_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_9_LC_12_22_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_9_LC_12_22_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_9_LC_12_22_4  (
            .in0(N__31279),
            .in1(N__31559),
            .in2(N__32002),
            .in3(N__32035),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto8_0_LC_12_22_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto8_0_LC_12_22_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto8_0_LC_12_22_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto8_0_LC_12_22_5  (
            .in0(_gnd_net_),
            .in1(N__32939),
            .in2(_gnd_net_),
            .in3(N__32656),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto8Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_6_LC_12_22_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_6_LC_12_22_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_6_LC_12_22_6 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_6_LC_12_22_6  (
            .in0(N__32827),
            .in1(_gnd_net_),
            .in2(N__31902),
            .in3(N__31156),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_12_LC_12_22_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_12_LC_12_22_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_12_LC_12_22_7 .LUT_INIT=16'b1010000000100000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_12_LC_12_22_7  (
            .in0(N__30670),
            .in1(N__31326),
            .in2(N__30664),
            .in3(N__32743),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_12_23_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_12_23_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_12_23_1 .LUT_INIT=16'b0100010001010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_9_LC_12_23_1  (
            .in0(N__31391),
            .in1(N__31992),
            .in2(_gnd_net_),
            .in3(N__31734),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50138),
            .ce(N__31583),
            .sr(N__49715));
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_12_23_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_12_23_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_12_23_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_12_LC_12_23_2  (
            .in0(N__31732),
            .in1(N__31280),
            .in2(_gnd_net_),
            .in3(N__31392),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50138),
            .ce(N__31583),
            .sr(N__49715));
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_12_23_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_12_23_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_12_23_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_11_LC_12_23_5  (
            .in0(N__31389),
            .in1(N__32036),
            .in2(_gnd_net_),
            .in3(N__31731),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50138),
            .ce(N__31583),
            .sr(N__49715));
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_12_23_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_12_23_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_12_23_7 .LUT_INIT=16'b0100010001010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_17_LC_12_23_7  (
            .in0(N__31390),
            .in1(N__31197),
            .in2(_gnd_net_),
            .in3(N__31733),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50138),
            .ce(N__31583),
            .sr(N__49715));
    defparam \delay_measurement_inst.delay_hc_reg_10_LC_12_24_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_10_LC_12_24_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_10_LC_12_24_0 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_10_LC_12_24_0  (
            .in0(N__41199),
            .in1(N__35578),
            .in2(N__31561),
            .in3(N__41047),
            .lcout(measured_delay_hc_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50135),
            .ce(),
            .sr(N__49724));
    defparam \delay_measurement_inst.delay_hc_reg_31_LC_12_24_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_31_LC_12_24_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_31_LC_12_24_5 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_31_LC_12_24_5  (
            .in0(N__41048),
            .in1(N__31401),
            .in2(_gnd_net_),
            .in3(N__41203),
            .lcout(measured_delay_hc_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50135),
            .ce(),
            .sr(N__49724));
    defparam \delay_measurement_inst.delay_hc_reg_3_LC_12_24_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_3_LC_12_24_6 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_hc_reg_3_LC_12_24_6 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_3_LC_12_24_6  (
            .in0(N__35209),
            .in1(N__31317),
            .in2(N__41219),
            .in3(N__41049),
            .lcout(measured_delay_hc_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50135),
            .ce(),
            .sr(N__49724));
    defparam \delay_measurement_inst.delay_hc_reg_12_LC_12_25_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_12_LC_12_25_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_12_LC_12_25_0 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_12_LC_12_25_0  (
            .in0(N__41017),
            .in1(N__35467),
            .in2(N__31282),
            .in3(N__41156),
            .lcout(measured_delay_hc_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50133),
            .ce(),
            .sr(N__49730));
    defparam \delay_measurement_inst.delay_hc_reg_18_LC_12_25_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_18_LC_12_25_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_18_LC_12_25_1 .LUT_INIT=16'b1111111111011000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_18_LC_12_25_1  (
            .in0(N__41154),
            .in1(N__39052),
            .in2(N__31245),
            .in3(N__41019),
            .lcout(measured_delay_hc_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50133),
            .ce(),
            .sr(N__49730));
    defparam \delay_measurement_inst.delay_hc_reg_17_LC_12_25_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_17_LC_12_25_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_17_LC_12_25_2 .LUT_INIT=16'b1110111011111010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_17_LC_12_25_2  (
            .in0(N__41018),
            .in1(N__39022),
            .in2(N__31201),
            .in3(N__41157),
            .lcout(measured_delay_hc_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50133),
            .ce(),
            .sr(N__49730));
    defparam \delay_measurement_inst.delay_hc_reg_5_LC_12_25_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_5_LC_12_25_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_5_LC_12_25_4 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_5_LC_12_25_4  (
            .in0(N__41020),
            .in1(N__31152),
            .in2(N__41220),
            .in3(N__35143),
            .lcout(measured_delay_hc_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50133),
            .ce(),
            .sr(N__49730));
    defparam \delay_measurement_inst.delay_hc_reg_11_LC_12_25_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_11_LC_12_25_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_11_LC_12_25_5 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_11_LC_12_25_5  (
            .in0(N__41153),
            .in1(N__35521),
            .in2(N__32038),
            .in3(N__41016),
            .lcout(measured_delay_hc_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50133),
            .ce(),
            .sr(N__49730));
    defparam \delay_measurement_inst.delay_hc_reg_9_LC_12_25_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_9_LC_12_25_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_9_LC_12_25_7 .LUT_INIT=16'b1111111111011000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_9_LC_12_25_7  (
            .in0(N__41155),
            .in1(N__34924),
            .in2(N__31996),
            .in3(N__41021),
            .lcout(measured_delay_hc_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50133),
            .ce(),
            .sr(N__49730));
    defparam \delay_measurement_inst.delay_hc_reg_24_LC_12_26_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_24_LC_12_26_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_24_LC_12_26_2 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_24_LC_12_26_2  (
            .in0(N__40980),
            .in1(_gnd_net_),
            .in2(N__41207),
            .in3(N__31807),
            .lcout(measured_delay_hc_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50131),
            .ce(),
            .sr(N__49735));
    defparam \delay_measurement_inst.delay_hc_reg_14_LC_12_26_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_14_LC_12_26_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_14_LC_12_26_3 .LUT_INIT=16'b1111111110111000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_14_LC_12_26_3  (
            .in0(N__35356),
            .in1(N__41159),
            .in2(N__31951),
            .in3(N__40979),
            .lcout(measured_delay_hc_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50131),
            .ce(),
            .sr(N__49735));
    defparam \delay_measurement_inst.delay_hc_reg_6_LC_12_26_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_6_LC_12_26_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_6_LC_12_26_4 .LUT_INIT=16'b1111111010101110;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_6_LC_12_26_4  (
            .in0(N__40982),
            .in1(N__31879),
            .in2(N__41209),
            .in3(N__35095),
            .lcout(measured_delay_hc_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50131),
            .ce(),
            .sr(N__49735));
    defparam \delay_measurement_inst.delay_hc_reg_25_LC_12_26_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_25_LC_12_26_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_25_LC_12_26_6 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_25_LC_12_26_6  (
            .in0(N__40981),
            .in1(_gnd_net_),
            .in2(N__41208),
            .in3(N__31795),
            .lcout(measured_delay_hc_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50131),
            .ce(),
            .sr(N__49735));
    defparam \delay_measurement_inst.delay_hc_reg_13_LC_12_26_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_13_LC_12_26_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_13_LC_12_26_7 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_13_LC_12_26_7  (
            .in0(N__35413),
            .in1(N__41158),
            .in2(N__31848),
            .in3(N__40978),
            .lcout(measured_delay_hc_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50131),
            .ce(),
            .sr(N__49735));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_1_4_LC_12_27_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_1_4_LC_12_27_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_1_4_LC_12_27_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto30_1_4_LC_12_27_5  (
            .in0(N__31806),
            .in1(N__31794),
            .in2(N__31783),
            .in3(N__32166),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_12_27_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_12_27_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_12_27_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_12_27_6  (
            .in0(N__35466),
            .in1(N__35517),
            .in2(N__35412),
            .in3(N__35577),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_LC_12_28_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_LC_12_28_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.running_LC_12_28_1 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \current_shift_inst.timer_s1.running_LC_12_28_1  (
            .in0(N__33177),
            .in1(N__43662),
            .in2(_gnd_net_),
            .in3(N__33319),
            .lcout(\current_shift_inst.timer_s1.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50127),
            .ce(),
            .sr(N__49739));
    defparam \delay_measurement_inst.delay_hc_reg_23_LC_12_28_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_23_LC_12_28_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_23_LC_12_28_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_23_LC_12_28_2  (
            .in0(N__41212),
            .in1(N__32167),
            .in2(_gnd_net_),
            .in3(N__40983),
            .lcout(measured_delay_hc_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50127),
            .ce(),
            .sr(N__49739));
    defparam \current_shift_inst.start_timer_s1_LC_12_28_5 .C_ON=1'b0;
    defparam \current_shift_inst.start_timer_s1_LC_12_28_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.start_timer_s1_LC_12_28_5 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \current_shift_inst.start_timer_s1_LC_12_28_5  (
            .in0(N__32075),
            .in1(N__33176),
            .in2(_gnd_net_),
            .in3(N__32147),
            .lcout(\current_shift_inst.start_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50127),
            .ce(),
            .sr(N__49739));
    defparam \current_shift_inst.stop_timer_s1_LC_12_29_2 .C_ON=1'b0;
    defparam \current_shift_inst.stop_timer_s1_LC_12_29_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.stop_timer_s1_LC_12_29_2 .LUT_INIT=16'b1111101100001000;
    LogicCell40 \current_shift_inst.stop_timer_s1_LC_12_29_2  (
            .in0(N__33178),
            .in1(N__32154),
            .in2(N__32082),
            .in3(N__33318),
            .lcout(\current_shift_inst.stop_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50126),
            .ce(),
            .sr(N__49744));
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_13_6_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_13_6_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_13_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_0_LC_13_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33838),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50240),
            .ce(),
            .sr(N__49616));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI637M_11_LC_13_7_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI637M_11_LC_13_7_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI637M_11_LC_13_7_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI637M_11_LC_13_7_2  (
            .in0(N__36906),
            .in1(N__41789),
            .in2(N__40270),
            .in3(N__41729),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_13_7_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_13_7_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_13_7_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_13_7_6  (
            .in0(N__39402),
            .in1(N__36517),
            .in2(_gnd_net_),
            .in3(N__39432),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un1_enablelt3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_13_7_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_13_7_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_13_7_7 .LUT_INIT=16'b1111111101010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_13_7_7  (
            .in0(N__39353),
            .in1(N__40873),
            .in2(N__32050),
            .in3(N__43495),
            .lcout(\current_shift_inst.PI_CTRL.N_71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_13_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_13_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_13_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_13_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36677),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_13_8_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_13_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_13_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_13_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36233),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_13_8_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_13_8_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_13_8_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_13_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36269),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_13_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_13_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_13_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_13_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36197),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_13_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_13_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_13_8_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_13_8_6  (
            .in0(N__32201),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_13_8_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_13_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_13_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_13_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36560),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_13_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_13_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_13_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_13_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36161),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIFLJ3_16_LC_13_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIFLJ3_16_LC_13_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIFLJ3_16_LC_13_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIFLJ3_16_LC_13_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36764),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_13_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_13_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_13_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_13_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36479),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_13_9_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_13_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_13_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_13_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36602),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_13_9_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_13_9_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_13_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_13_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36638),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNICIJ3_13_LC_13_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNICIJ3_13_LC_13_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNICIJ3_13_LC_13_9_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNICIJ3_13_LC_13_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36311),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIEKJ3_15_LC_13_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIEKJ3_15_LC_13_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIEKJ3_15_LC_13_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIEKJ3_15_LC_13_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36854),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_14_LC_13_9_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_14_LC_13_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_14_LC_13_9_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_14_LC_13_9_7  (
            .in0(N__43859),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_13_10_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_13_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_13_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_13_10_0  (
            .in0(_gnd_net_),
            .in1(N__32248),
            .in2(_gnd_net_),
            .in3(N__33834),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ),
            .ltout(),
            .carryin(bfn_13_10_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_13_10_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_13_10_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_13_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_1_LC_13_10_1  (
            .in0(_gnd_net_),
            .in1(N__33628),
            .in2(_gnd_net_),
            .in3(N__32242),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .clk(N__50211),
            .ce(),
            .sr(N__49629));
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_13_10_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_13_10_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_13_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_LC_13_10_2  (
            .in0(_gnd_net_),
            .in1(N__33862),
            .in2(_gnd_net_),
            .in3(N__32239),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .clk(N__50211),
            .ce(),
            .sr(N__49629));
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_13_10_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_13_10_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_13_10_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_3_LC_13_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33727),
            .in3(N__32236),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .clk(N__50211),
            .ce(),
            .sr(N__49629));
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_13_10_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_13_10_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_13_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_4_LC_13_10_4  (
            .in0(_gnd_net_),
            .in1(N__32233),
            .in2(_gnd_net_),
            .in3(N__32221),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .clk(N__50211),
            .ce(),
            .sr(N__49629));
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_13_10_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_13_10_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_13_10_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_5_LC_13_10_5  (
            .in0(_gnd_net_),
            .in1(N__33706),
            .in2(_gnd_net_),
            .in3(N__32218),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .clk(N__50211),
            .ce(),
            .sr(N__49629));
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_13_10_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_13_10_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_13_10_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_6_LC_13_10_6  (
            .in0(_gnd_net_),
            .in1(N__32356),
            .in2(_gnd_net_),
            .in3(N__32215),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .clk(N__50211),
            .ce(),
            .sr(N__49629));
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_13_10_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_13_10_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_13_10_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_7_LC_13_10_7  (
            .in0(_gnd_net_),
            .in1(N__33592),
            .in2(_gnd_net_),
            .in3(N__32281),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .clk(N__50211),
            .ce(),
            .sr(N__49629));
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_13_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_13_11_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_13_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_8_LC_13_11_0  (
            .in0(_gnd_net_),
            .in1(N__33748),
            .in2(_gnd_net_),
            .in3(N__32278),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_8 ),
            .ltout(),
            .carryin(bfn_13_11_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .clk(N__50207),
            .ce(),
            .sr(N__49638));
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_13_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_13_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_13_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_9_LC_13_11_1  (
            .in0(_gnd_net_),
            .in1(N__32275),
            .in2(_gnd_net_),
            .in3(N__32269),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .clk(N__50207),
            .ce(),
            .sr(N__49638));
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_13_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_13_11_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_13_11_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_10_LC_13_11_2  (
            .in0(_gnd_net_),
            .in1(N__33742),
            .in2(_gnd_net_),
            .in3(N__32266),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .clk(N__50207),
            .ce(),
            .sr(N__49638));
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_13_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_13_11_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_13_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_11_LC_13_11_3  (
            .in0(_gnd_net_),
            .in1(N__33652),
            .in2(_gnd_net_),
            .in3(N__32263),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .clk(N__50207),
            .ce(),
            .sr(N__49638));
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_13_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_13_11_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_13_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_12_LC_13_11_4  (
            .in0(_gnd_net_),
            .in1(N__33697),
            .in2(_gnd_net_),
            .in3(N__32260),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ),
            .clk(N__50207),
            .ce(),
            .sr(N__49638));
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_13_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_13_11_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_13_11_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_13_LC_13_11_5  (
            .in0(_gnd_net_),
            .in1(N__33664),
            .in2(_gnd_net_),
            .in3(N__32257),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ),
            .clk(N__50207),
            .ce(),
            .sr(N__49638));
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_13_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_13_11_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_13_11_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_14_LC_13_11_6  (
            .in0(_gnd_net_),
            .in1(N__33715),
            .in2(_gnd_net_),
            .in3(N__32254),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_14 ),
            .clk(N__50207),
            .ce(),
            .sr(N__49638));
    defparam \current_shift_inst.PI_CTRL.error_control_15_LC_13_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_15_LC_13_11_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_15_LC_13_11_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_15_LC_13_11_7  (
            .in0(_gnd_net_),
            .in1(N__34060),
            .in2(_gnd_net_),
            .in3(N__32251),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_15 ),
            .clk(N__50207),
            .ce(),
            .sr(N__49638));
    defparam \current_shift_inst.PI_CTRL.error_control_16_LC_13_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_16_LC_13_12_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_16_LC_13_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_16_LC_13_12_0  (
            .in0(_gnd_net_),
            .in1(N__33658),
            .in2(_gnd_net_),
            .in3(N__32320),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_16 ),
            .ltout(),
            .carryin(bfn_13_12_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_16 ),
            .clk(N__50201),
            .ce(),
            .sr(N__49644));
    defparam \current_shift_inst.PI_CTRL.error_control_17_LC_13_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_17_LC_13_12_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_17_LC_13_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_17_LC_13_12_1  (
            .in0(_gnd_net_),
            .in1(N__33277),
            .in2(_gnd_net_),
            .in3(N__32317),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_17 ),
            .clk(N__50201),
            .ce(),
            .sr(N__49644));
    defparam \current_shift_inst.PI_CTRL.error_control_18_LC_13_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_18_LC_13_12_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_18_LC_13_12_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_18_LC_13_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33736),
            .in3(N__32314),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_18 ),
            .clk(N__50201),
            .ce(),
            .sr(N__49644));
    defparam \current_shift_inst.PI_CTRL.error_control_19_LC_13_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_19_LC_13_12_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_19_LC_13_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_19_LC_13_12_3  (
            .in0(_gnd_net_),
            .in1(N__33676),
            .in2(_gnd_net_),
            .in3(N__32311),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_19 ),
            .clk(N__50201),
            .ce(),
            .sr(N__49644));
    defparam \current_shift_inst.PI_CTRL.error_control_20_LC_13_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_20_LC_13_12_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_20_LC_13_12_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_20_LC_13_12_4  (
            .in0(_gnd_net_),
            .in1(N__33619),
            .in2(_gnd_net_),
            .in3(N__32308),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_20 ),
            .clk(N__50201),
            .ce(),
            .sr(N__49644));
    defparam \current_shift_inst.PI_CTRL.error_control_21_LC_13_12_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_21_LC_13_12_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_21_LC_13_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_21_LC_13_12_5  (
            .in0(_gnd_net_),
            .in1(N__32329),
            .in2(_gnd_net_),
            .in3(N__32305),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_21 ),
            .clk(N__50201),
            .ce(),
            .sr(N__49644));
    defparam \current_shift_inst.PI_CTRL.error_control_22_LC_13_12_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_22_LC_13_12_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_22_LC_13_12_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_22_LC_13_12_6  (
            .in0(_gnd_net_),
            .in1(N__32302),
            .in2(_gnd_net_),
            .in3(N__32290),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_22 ),
            .clk(N__50201),
            .ce(),
            .sr(N__49644));
    defparam \current_shift_inst.PI_CTRL.error_control_23_LC_13_12_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_23_LC_13_12_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_23_LC_13_12_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_23_LC_13_12_7  (
            .in0(_gnd_net_),
            .in1(N__33850),
            .in2(_gnd_net_),
            .in3(N__32287),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_23 ),
            .clk(N__50201),
            .ce(),
            .sr(N__49644));
    defparam \current_shift_inst.PI_CTRL.error_control_24_LC_13_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_24_LC_13_13_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_24_LC_13_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_24_LC_13_13_0  (
            .in0(_gnd_net_),
            .in1(N__32335),
            .in2(_gnd_net_),
            .in3(N__32284),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_24 ),
            .ltout(),
            .carryin(bfn_13_13_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_24 ),
            .clk(N__50193),
            .ce(),
            .sr(N__49649));
    defparam \current_shift_inst.PI_CTRL.error_control_25_LC_13_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_25_LC_13_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_25_LC_13_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_25_LC_13_13_1  (
            .in0(_gnd_net_),
            .in1(N__32341),
            .in2(_gnd_net_),
            .in3(N__32347),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_25 ),
            .clk(N__50193),
            .ce(),
            .sr(N__49649));
    defparam \current_shift_inst.PI_CTRL.error_control_26_LC_13_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_26_LC_13_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_26_LC_13_13_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_26_LC_13_13_2  (
            .in0(_gnd_net_),
            .in1(N__34387),
            .in2(_gnd_net_),
            .in3(N__32344),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50193),
            .ce(),
            .sr(N__49649));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_13_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_13_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_13_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_13_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34386),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_13_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_13_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_13_13_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_13_13_6  (
            .in0(N__34417),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_13_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_13_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_13_14_0 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_13_14_0  (
            .in0(N__38614),
            .in1(N__32554),
            .in2(_gnd_net_),
            .in3(N__46993),
            .lcout(\current_shift_inst.control_input_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_13_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_13_14_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_13_14_2  (
            .in0(N__34462),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_13_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_13_14_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_13_14_3  (
            .in0(N__46744),
            .in1(N__48190),
            .in2(N__46341),
            .in3(N__42819),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_13_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_13_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_13_14_4 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_13_14_4  (
            .in0(N__32488),
            .in1(N__38557),
            .in2(_gnd_net_),
            .in3(N__46994),
            .lcout(\current_shift_inst.control_input_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_13_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_13_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_13_14_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_13_14_5  (
            .in0(N__46743),
            .in1(N__47590),
            .in2(N__46340),
            .in3(N__42880),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_13_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_13_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_13_14_6 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_13_14_6  (
            .in0(N__46026),
            .in1(N__46745),
            .in2(N__48586),
            .in3(N__43060),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_13_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_13_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_13_14_7 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_13_14_7  (
            .in0(N__46995),
            .in1(N__38503),
            .in2(_gnd_net_),
            .in3(N__32635),
            .lcout(\current_shift_inst.control_input_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_13_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_13_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_13_15_0 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_13_15_0  (
            .in0(N__38485),
            .in1(N__32620),
            .in2(_gnd_net_),
            .in3(N__46973),
            .lcout(\current_shift_inst.control_input_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_13_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_13_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_13_15_1 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_13_15_1  (
            .in0(N__46974),
            .in1(N__38734),
            .in2(_gnd_net_),
            .in3(N__32608),
            .lcout(\current_shift_inst.control_input_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_13_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_13_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_13_15_2 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_13_15_2  (
            .in0(N__32371),
            .in1(N__38419),
            .in2(_gnd_net_),
            .in3(N__46969),
            .lcout(\current_shift_inst.control_input_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_13_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_13_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_13_15_3 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_13_15_3  (
            .in0(N__47905),
            .in1(N__42558),
            .in2(N__46228),
            .in3(N__46707),
            .lcout(\current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_13_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_13_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_13_15_4 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_13_15_4  (
            .in0(N__38593),
            .in1(N__32521),
            .in2(_gnd_net_),
            .in3(N__46970),
            .lcout(\current_shift_inst.control_input_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_13_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_13_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_13_15_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_13_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34180),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_13_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_13_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_13_15_6 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_13_15_6  (
            .in0(N__32473),
            .in1(N__38539),
            .in2(_gnd_net_),
            .in3(N__46971),
            .lcout(\current_shift_inst.control_input_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_13_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_13_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_13_15_7 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_13_15_7  (
            .in0(N__46972),
            .in1(N__38521),
            .in2(_gnd_net_),
            .in3(N__32458),
            .lcout(\current_shift_inst.control_input_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_13_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_13_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_13_16_0 .LUT_INIT=16'b1111010100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_13_16_0  (
            .in0(N__47800),
            .in1(N__46006),
            .in2(N__46742),
            .in3(N__42999),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_13_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_13_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_13_16_1 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_13_16_1  (
            .in0(N__32581),
            .in1(N__38701),
            .in2(_gnd_net_),
            .in3(N__46980),
            .lcout(\current_shift_inst.control_input_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_13_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_13_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_13_16_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_13_16_2  (
            .in0(N__46651),
            .in1(N__47713),
            .in2(N__46217),
            .in3(N__42936),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_13_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_13_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_13_16_3 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_13_16_3  (
            .in0(N__32500),
            .in1(N__38575),
            .in2(_gnd_net_),
            .in3(N__46979),
            .lcout(\current_shift_inst.control_input_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_13_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_13_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_13_16_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_13_16_4  (
            .in0(N__46647),
            .in1(N__47833),
            .in2(N__46218),
            .in3(N__47407),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_13_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_13_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_13_16_5 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_13_16_5  (
            .in0(N__38449),
            .in1(N__32410),
            .in2(_gnd_net_),
            .in3(N__46975),
            .lcout(\current_shift_inst.control_input_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_13_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_13_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_13_16_6 .LUT_INIT=16'b0000001111110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_13_16_6  (
            .in0(_gnd_net_),
            .in1(N__38434),
            .in2(N__46992),
            .in3(N__32392),
            .lcout(\current_shift_inst.control_input_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_13_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_13_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_13_16_7 .LUT_INIT=16'b1111001100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_13_16_7  (
            .in0(N__46007),
            .in1(N__48235),
            .in2(N__46797),
            .in3(N__42846),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_13_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_13_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_LC_13_17_0  (
            .in0(_gnd_net_),
            .in1(N__32362),
            .in2(N__37975),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_17_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_13_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_13_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_13_17_1  (
            .in0(_gnd_net_),
            .in1(N__40438),
            .in2(N__40417),
            .in3(N__37843),
            .lcout(\current_shift_inst.un38_control_input_5_1 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_13_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_13_17_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_13_17_2  (
            .in0(N__37844),
            .in1(N__32446),
            .in2(N__45925),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un38_control_input_5_2 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_LC_13_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_LC_13_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_LC_13_17_3  (
            .in0(_gnd_net_),
            .in1(N__40099),
            .in2(N__45928),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_LC_13_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_LC_13_17_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_LC_13_17_4  (
            .in0(_gnd_net_),
            .in1(N__45547),
            .in2(N__45926),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_LC_13_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_LC_13_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_LC_13_17_5  (
            .in0(_gnd_net_),
            .in1(N__32440),
            .in2(N__45929),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_13_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_13_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_13_17_6  (
            .in0(_gnd_net_),
            .in1(N__45532),
            .in2(N__45927),
            .in3(N__32431),
            .lcout(\current_shift_inst.un38_control_input_0_s0_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_13_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_13_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_13_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_13_17_7  (
            .in0(_gnd_net_),
            .in1(N__32428),
            .in2(N__45930),
            .in3(N__32422),
            .lcout(\current_shift_inst.un38_control_input_0_s0_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_13_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_13_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_13_18_0  (
            .in0(_gnd_net_),
            .in1(N__32419),
            .in2(N__45991),
            .in3(N__32401),
            .lcout(\current_shift_inst.un38_control_input_0_s0_8 ),
            .ltout(),
            .carryin(bfn_13_18_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_13_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_13_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_13_18_1  (
            .in0(_gnd_net_),
            .in1(N__32398),
            .in2(N__45995),
            .in3(N__32383),
            .lcout(\current_shift_inst.un38_control_input_0_s0_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_13_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_13_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_13_18_2  (
            .in0(_gnd_net_),
            .in1(N__32380),
            .in2(N__45992),
            .in3(N__32560),
            .lcout(\current_shift_inst.un38_control_input_0_s0_10 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_13_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_13_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_13_18_3  (
            .in0(_gnd_net_),
            .in1(N__47095),
            .in2(N__45996),
            .in3(N__32557),
            .lcout(\current_shift_inst.un38_control_input_0_s0_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_13_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_13_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_13_18_4  (
            .in0(_gnd_net_),
            .in1(N__34513),
            .in2(N__45993),
            .in3(N__32545),
            .lcout(\current_shift_inst.un38_control_input_0_s0_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_13_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_13_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_13_18_5  (
            .in0(_gnd_net_),
            .in1(N__32542),
            .in2(N__45997),
            .in3(N__32533),
            .lcout(\current_shift_inst.un38_control_input_0_s0_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_13_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_13_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_13_18_6  (
            .in0(_gnd_net_),
            .in1(N__32530),
            .in2(N__45994),
            .in3(N__32512),
            .lcout(\current_shift_inst.un38_control_input_0_s0_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_13_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_13_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_13_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_13_18_7  (
            .in0(_gnd_net_),
            .in1(N__32509),
            .in2(N__45998),
            .in3(N__32491),
            .lcout(\current_shift_inst.un38_control_input_0_s0_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_13_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_13_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_13_19_0  (
            .in0(_gnd_net_),
            .in1(N__45959),
            .in2(N__45487),
            .in3(N__32476),
            .lcout(\current_shift_inst.un38_control_input_0_s0_16 ),
            .ltout(),
            .carryin(bfn_13_19_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_13_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_13_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_13_19_1  (
            .in0(_gnd_net_),
            .in1(N__43351),
            .in2(N__46208),
            .in3(N__32461),
            .lcout(\current_shift_inst.un38_control_input_0_s0_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_13_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_13_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_13_19_2  (
            .in0(_gnd_net_),
            .in1(N__45963),
            .in2(N__34507),
            .in3(N__32449),
            .lcout(\current_shift_inst.un38_control_input_0_s0_18 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_13_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_13_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_13_19_3  (
            .in0(_gnd_net_),
            .in1(N__40591),
            .in2(N__46209),
            .in3(N__32623),
            .lcout(\current_shift_inst.un38_control_input_0_s0_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_13_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_13_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_13_19_4  (
            .in0(_gnd_net_),
            .in1(N__45967),
            .in2(N__40681),
            .in3(N__32611),
            .lcout(\current_shift_inst.un38_control_input_0_s0_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_13_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_13_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_13_19_5  (
            .in0(_gnd_net_),
            .in1(N__34483),
            .in2(N__46210),
            .in3(N__32599),
            .lcout(\current_shift_inst.un38_control_input_0_s0_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_13_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_13_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_13_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_13_19_6  (
            .in0(_gnd_net_),
            .in1(N__45971),
            .in2(N__32596),
            .in3(N__32584),
            .lcout(\current_shift_inst.un38_control_input_0_s0_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_13_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_13_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_13_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_13_19_7  (
            .in0(_gnd_net_),
            .in1(N__45999),
            .in2(N__43150),
            .in3(N__32572),
            .lcout(\current_shift_inst.un38_control_input_0_s0_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_13_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_13_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_13_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_13_20_0  (
            .in0(_gnd_net_),
            .in1(N__34600),
            .in2(N__46211),
            .in3(N__32569),
            .lcout(\current_shift_inst.un38_control_input_0_s0_24 ),
            .ltout(),
            .carryin(bfn_13_20_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_13_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_13_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_13_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_13_20_1  (
            .in0(_gnd_net_),
            .in1(N__43681),
            .in2(N__46215),
            .in3(N__32566),
            .lcout(\current_shift_inst.un38_control_input_0_s0_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_13_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_13_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_13_20_2  (
            .in0(_gnd_net_),
            .in1(N__34606),
            .in2(N__46212),
            .in3(N__32563),
            .lcout(\current_shift_inst.un38_control_input_0_s0_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_13_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_13_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_13_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_13_20_3  (
            .in0(_gnd_net_),
            .in1(N__43300),
            .in2(N__46216),
            .in3(N__32758),
            .lcout(\current_shift_inst.un38_control_input_0_s0_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_13_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_13_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_13_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_13_20_4  (
            .in0(_gnd_net_),
            .in1(N__34612),
            .in2(N__46213),
            .in3(N__32755),
            .lcout(\current_shift_inst.un38_control_input_0_s0_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_13_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_13_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_13_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_13_20_5  (
            .in0(_gnd_net_),
            .in1(N__45981),
            .in2(N__40711),
            .in3(N__32752),
            .lcout(\current_shift_inst.un38_control_input_0_s0_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNII18T_LC_13_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNII18T_LC_13_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNII18T_LC_13_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNII18T_LC_13_20_6  (
            .in0(_gnd_net_),
            .in1(N__40783),
            .in2(N__46214),
            .in3(N__32749),
            .lcout(\current_shift_inst.un38_control_input_0_s0_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_RNO_0_25_LC_13_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_RNO_0_25_LC_13_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_RNO_0_25_LC_13_20_7 .LUT_INIT=16'b1010001101010011;
    LogicCell40 \current_shift_inst.control_input_RNO_0_25_LC_13_20_7  (
            .in0(N__45457),
            .in1(N__39064),
            .in2(N__46996),
            .in3(N__32746),
            .lcout(\current_shift_inst.control_input_1_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto5_2_LC_13_21_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto5_2_LC_13_21_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto5_2_LC_13_21_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto5_2_LC_13_21_5  (
            .in0(_gnd_net_),
            .in1(N__32778),
            .in2(_gnd_net_),
            .in3(N__32974),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlt3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_1_LC_13_22_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_1_LC_13_22_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_1_LC_13_22_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_26_1_LC_13_22_2  (
            .in0(N__33042),
            .in1(N__32690),
            .in2(N__33135),
            .in3(N__32911),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_1_6_LC_13_22_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_1_6_LC_13_22_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_1_6_LC_13_22_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto30_1_6_LC_13_22_5  (
            .in0(N__32910),
            .in1(N__33041),
            .in2(N__32692),
            .in3(N__38776),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_22_LC_13_23_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_22_LC_13_23_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_22_LC_13_23_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_22_LC_13_23_0  (
            .in0(N__41185),
            .in1(N__32691),
            .in2(_gnd_net_),
            .in3(N__41038),
            .lcout(measured_delay_hc_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50144),
            .ce(),
            .sr(N__49708));
    defparam \delay_measurement_inst.delay_hc_reg_7_LC_13_23_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_7_LC_13_23_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_7_LC_13_23_1 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_7_LC_13_23_1  (
            .in0(N__41039),
            .in1(N__41186),
            .in2(N__32672),
            .in3(N__35044),
            .lcout(measured_delay_hc_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50144),
            .ce(),
            .sr(N__49708));
    defparam \delay_measurement_inst.delay_hc_reg_0_LC_13_23_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_0_LC_13_23_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_0_LC_13_23_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_0_LC_13_23_2  (
            .in0(N__41183),
            .in1(N__33067),
            .in2(_gnd_net_),
            .in3(N__41036),
            .lcout(measured_delay_hc_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50144),
            .ce(),
            .sr(N__49708));
    defparam \delay_measurement_inst.delay_hc_reg_20_LC_13_23_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_20_LC_13_23_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_20_LC_13_23_6 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_20_LC_13_23_6  (
            .in0(N__41184),
            .in1(N__33043),
            .in2(_gnd_net_),
            .in3(N__41037),
            .lcout(measured_delay_hc_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50144),
            .ce(),
            .sr(N__49708));
    defparam \delay_measurement_inst.delay_hc_reg_16_LC_13_24_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_16_LC_13_24_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_16_LC_13_24_0 .LUT_INIT=16'b1111111111011000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_16_LC_13_24_0  (
            .in0(N__41195),
            .in1(N__38992),
            .in2(N__33021),
            .in3(N__41032),
            .lcout(measured_delay_hc_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50139),
            .ce(),
            .sr(N__49716));
    defparam \delay_measurement_inst.delay_hc_reg_1_LC_13_24_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_1_LC_13_24_1 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_hc_reg_1_LC_13_24_1 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_1_LC_13_24_1  (
            .in0(N__41033),
            .in1(N__41197),
            .in2(N__32981),
            .in3(N__38881),
            .lcout(measured_delay_hc_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50139),
            .ce(),
            .sr(N__49716));
    defparam \delay_measurement_inst.delay_hc_reg_8_LC_13_24_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_8_LC_13_24_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_8_LC_13_24_2 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_8_LC_13_24_2  (
            .in0(N__41196),
            .in1(N__32938),
            .in2(N__34987),
            .in3(N__41035),
            .lcout(measured_delay_hc_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50139),
            .ce(),
            .sr(N__49716));
    defparam \delay_measurement_inst.delay_hc_reg_21_LC_13_24_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_21_LC_13_24_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_21_LC_13_24_5 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_21_LC_13_24_5  (
            .in0(N__41034),
            .in1(N__32909),
            .in2(_gnd_net_),
            .in3(N__41198),
            .lcout(measured_delay_hc_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50139),
            .ce(),
            .sr(N__49716));
    defparam \delay_measurement_inst.delay_hc_reg_15_LC_13_25_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_15_LC_13_25_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_15_LC_13_25_1 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_15_LC_13_25_1  (
            .in0(N__35299),
            .in1(N__41169),
            .in2(N__32889),
            .in3(N__41012),
            .lcout(measured_delay_hc_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50136),
            .ce(),
            .sr(N__49725));
    defparam \delay_measurement_inst.delay_hc_reg_4_LC_13_25_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_4_LC_13_25_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_4_LC_13_25_4 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_4_LC_13_25_4  (
            .in0(N__41015),
            .in1(N__35185),
            .in2(N__41211),
            .in3(N__32823),
            .lcout(measured_delay_hc_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50136),
            .ce(),
            .sr(N__49725));
    defparam \delay_measurement_inst.delay_hc_reg_2_LC_13_25_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_2_LC_13_25_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_2_LC_13_25_6 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_2_LC_13_25_6  (
            .in0(N__41014),
            .in1(N__32777),
            .in2(N__41210),
            .in3(N__38836),
            .lcout(measured_delay_hc_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50136),
            .ce(),
            .sr(N__49725));
    defparam \delay_measurement_inst.delay_hc_reg_19_LC_13_25_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_19_LC_13_25_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_19_LC_13_25_7 .LUT_INIT=16'b1111111110111000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_19_LC_13_25_7  (
            .in0(N__38960),
            .in1(N__41170),
            .in2(N__33134),
            .in3(N__41013),
            .lcout(measured_delay_hc_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50136),
            .ce(),
            .sr(N__49725));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI64F91_1_LC_13_26_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI64F91_1_LC_13_26_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI64F91_1_LC_13_26_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI64F91_1_LC_13_26_1  (
            .in0(N__35135),
            .in1(N__38832),
            .in2(_gnd_net_),
            .in3(N__38877),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto5_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHDUI2_3_LC_13_26_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHDUI2_3_LC_13_26_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHDUI2_3_LC_13_26_2 .LUT_INIT=16'b1110111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHDUI2_3_LC_13_26_2  (
            .in0(N__35183),
            .in1(N__35201),
            .in2(N__33103),
            .in3(N__35089),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI64AN1_6_LC_13_26_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI64AN1_6_LC_13_26_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI64AN1_6_LC_13_26_3 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI64AN1_6_LC_13_26_3  (
            .in0(N__35090),
            .in1(N__35038),
            .in2(N__34986),
            .in3(N__34912),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt13_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_13_LC_13_26_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_13_LC_13_26_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_13_LC_13_26_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_13_LC_13_26_4  (
            .in0(N__35402),
            .in1(N__38978),
            .in2(N__34920),
            .in3(N__35091),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_11_LC_13_26_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_11_LC_13_26_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_11_LC_13_26_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_11_LC_13_26_5  (
            .in0(N__33214),
            .in1(N__33094),
            .in2(N__33100),
            .in3(N__35215),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclt31_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOVQ9D_14_LC_13_26_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOVQ9D_14_LC_13_26_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOVQ9D_14_LC_13_26_6 .LUT_INIT=16'b0000110000000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOVQ9D_14_LC_13_26_6  (
            .in0(N__38935),
            .in1(N__33328),
            .in2(N__33097),
            .in3(N__33082),
            .lcout(\delay_measurement_inst.un1_elapsed_time_hc ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_17_LC_13_26_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_17_LC_13_26_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_17_LC_13_26_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_17_LC_13_26_7  (
            .in0(N__35136),
            .in1(N__39017),
            .in2(N__39047),
            .in3(N__35184),
            .lcout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINEU73_14_LC_13_27_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINEU73_14_LC_13_27_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINEU73_14_LC_13_27_3 .LUT_INIT=16'b0000000001110101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINEU73_14_LC_13_27_3  (
            .in0(N__35348),
            .in1(N__33088),
            .in2(N__33202),
            .in3(N__35293),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOJD01_11_LC_13_27_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOJD01_11_LC_13_27_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOJD01_11_LC_13_27_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOJD01_11_LC_13_27_4  (
            .in0(N__35347),
            .in1(N__35459),
            .in2(N__35298),
            .in3(N__35516),
            .lcout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI72ES3_7_LC_13_27_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI72ES3_7_LC_13_27_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI72ES3_7_LC_13_27_5 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI72ES3_7_LC_13_27_5  (
            .in0(N__34916),
            .in1(N__35039),
            .in2(N__34982),
            .in3(N__33208),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOC2D5_14_LC_13_27_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOC2D5_14_LC_13_27_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOC2D5_14_LC_13_27_6 .LUT_INIT=16'b0000001000110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOC2D5_14_LC_13_27_6  (
            .in0(N__33198),
            .in1(N__35294),
            .in2(N__33184),
            .in3(N__35349),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt19_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_13_27_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_13_27_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_13_27_7 .LUT_INIT=16'b0000001000110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_13_27_7  (
            .in0(N__38934),
            .in1(N__35914),
            .in2(N__33181),
            .in3(N__33151),
            .lcout(\delay_measurement_inst.delay_hc_reg3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILLI01_20_LC_13_28_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILLI01_20_LC_13_28_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILLI01_20_LC_13_28_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILLI01_20_LC_13_28_0  (
            .in0(N__35910),
            .in1(N__35718),
            .in2(N__35797),
            .in3(N__35755),
            .lcout(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_28_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_28_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_28_3 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_28_3  (
            .in0(N__43661),
            .in1(N__33175),
            .in2(_gnd_net_),
            .in3(N__33317),
            .lcout(\current_shift_inst.timer_s1.N_181_i_g ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_13_28_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_13_28_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_13_28_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_13_28_4  (
            .in0(_gnd_net_),
            .in1(N__35754),
            .in2(_gnd_net_),
            .in3(N__35719),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JIP2_20_LC_13_28_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JIP2_20_LC_13_28_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JIP2_20_LC_13_28_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JIP2_20_LC_13_28_5  (
            .in0(N__35796),
            .in1(N__33285),
            .in2(N__33154),
            .in3(N__33145),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_13_28_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_13_28_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_13_28_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_13_28_6  (
            .in0(N__35617),
            .in1(N__35647),
            .in2(N__36112),
            .in3(N__35680),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02O13_20_LC_13_28_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02O13_20_LC_13_28_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02O13_20_LC_13_28_7 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02O13_20_LC_13_28_7  (
            .in0(_gnd_net_),
            .in1(N__33337),
            .in2(N__33331),
            .in3(N__33286),
            .lcout(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_29_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_29_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_29_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.timer_s1.running_RNII51H_LC_13_29_1  (
            .in0(_gnd_net_),
            .in1(N__43657),
            .in2(_gnd_net_),
            .in3(N__33316),
            .lcout(\current_shift_inst.timer_s1.N_180_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_13_29_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_13_29_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_13_29_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_13_29_2  (
            .in0(N__35980),
            .in1(N__36034),
            .in2(N__35929),
            .in3(N__36073),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_14_6_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_14_6_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_14_6_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_14_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41779),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_14_6_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_14_6_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_14_6_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_14_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34249),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_14_6_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_14_6_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_14_6_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_14_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39465),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_14_6_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_14_6_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_14_6_7 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_14_6_7  (
            .in0(_gnd_net_),
            .in1(N__43469),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_14_7_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_14_7_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_14_7_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_14_7_0  (
            .in0(N__33258),
            .in1(N__33247),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_0 ),
            .ltout(),
            .carryin(bfn_14_7_0_),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_14_7_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_14_7_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_14_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_14_7_1  (
            .in0(_gnd_net_),
            .in1(N__33220),
            .in2(_gnd_net_),
            .in3(N__33237),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_14_7_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_14_7_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_14_7_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_14_7_2  (
            .in0(_gnd_net_),
            .in1(N__33427),
            .in2(_gnd_net_),
            .in3(N__33450),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_14_7_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_14_7_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_14_7_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_14_7_3  (
            .in0(_gnd_net_),
            .in1(N__33403),
            .in2(_gnd_net_),
            .in3(N__33420),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_14_7_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_14_7_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_14_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_14_7_4  (
            .in0(_gnd_net_),
            .in1(N__33397),
            .in2(_gnd_net_),
            .in3(N__33391),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_14_7_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_14_7_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_14_7_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_14_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33388),
            .in3(N__33379),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_14_7_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_14_7_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_14_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_14_7_6  (
            .in0(_gnd_net_),
            .in1(N__33376),
            .in2(_gnd_net_),
            .in3(N__33370),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_14_7_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_14_7_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_14_7_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_14_7_7  (
            .in0(_gnd_net_),
            .in1(N__33367),
            .in2(_gnd_net_),
            .in3(N__33358),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_14_8_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_14_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_14_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_14_8_0  (
            .in0(_gnd_net_),
            .in1(N__33355),
            .in2(_gnd_net_),
            .in3(N__33349),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_8 ),
            .ltout(),
            .carryin(bfn_14_8_0_),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_14_8_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_14_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_14_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_14_8_1  (
            .in0(_gnd_net_),
            .in1(N__33346),
            .in2(_gnd_net_),
            .in3(N__33340),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_14_8_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_14_8_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_14_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_14_8_2  (
            .in0(_gnd_net_),
            .in1(N__33520),
            .in2(_gnd_net_),
            .in3(N__33514),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_14_8_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_14_8_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_14_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_14_8_3  (
            .in0(_gnd_net_),
            .in1(N__33511),
            .in2(_gnd_net_),
            .in3(N__33505),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNI9BCC_LC_14_8_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNI9BCC_LC_14_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNI9BCC_LC_14_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNI9BCC_LC_14_8_4  (
            .in0(_gnd_net_),
            .in1(N__33502),
            .in2(_gnd_net_),
            .in3(N__33496),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNIBEDC_LC_14_8_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNIBEDC_LC_14_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNIBEDC_LC_14_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNIBEDC_LC_14_8_5  (
            .in0(_gnd_net_),
            .in1(N__33493),
            .in2(_gnd_net_),
            .in3(N__33487),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIDHEC_LC_14_8_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIDHEC_LC_14_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIDHEC_LC_14_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIDHEC_LC_14_8_6  (
            .in0(_gnd_net_),
            .in1(N__33484),
            .in2(_gnd_net_),
            .in3(N__33478),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIFKFC_LC_14_8_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIFKFC_LC_14_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIFKFC_LC_14_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNIFKFC_LC_14_8_7  (
            .in0(_gnd_net_),
            .in1(N__33475),
            .in2(_gnd_net_),
            .in3(N__33469),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIHNGC_LC_14_9_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIHNGC_LC_14_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIHNGC_LC_14_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIHNGC_LC_14_9_0  (
            .in0(_gnd_net_),
            .in1(N__33466),
            .in2(_gnd_net_),
            .in3(N__33460),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_16 ),
            .ltout(),
            .carryin(bfn_14_9_0_),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIJQHC_LC_14_9_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIJQHC_LC_14_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIJQHC_LC_14_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIJQHC_LC_14_9_1  (
            .in0(_gnd_net_),
            .in1(N__33586),
            .in2(_gnd_net_),
            .in3(N__33457),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNILTIC_LC_14_9_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNILTIC_LC_14_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNILTIC_LC_14_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNILTIC_LC_14_9_2  (
            .in0(_gnd_net_),
            .in1(N__33601),
            .in2(_gnd_net_),
            .in3(N__33454),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIN0KC_LC_14_9_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIN0KC_LC_14_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIN0KC_LC_14_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNIN0KC_LC_14_9_3  (
            .in0(_gnd_net_),
            .in1(N__33568),
            .in2(_gnd_net_),
            .in3(N__33559),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNIGRLC_LC_14_9_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNIGRLC_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNIGRLC_LC_14_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNIGRLC_LC_14_9_4  (
            .in0(_gnd_net_),
            .in1(N__33637),
            .in2(_gnd_net_),
            .in3(N__33556),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNI9DFD_LC_14_9_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNI9DFD_LC_14_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNI9DFD_LC_14_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNI9DFD_LC_14_9_5  (
            .in0(_gnd_net_),
            .in1(N__33646),
            .in2(_gnd_net_),
            .in3(N__33553),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIBGGD_LC_14_9_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIBGGD_LC_14_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIBGGD_LC_14_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNIBGGD_LC_14_9_6  (
            .in0(_gnd_net_),
            .in1(N__33577),
            .in2(_gnd_net_),
            .in3(N__33550),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIDJHD_LC_14_9_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIDJHD_LC_14_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIDJHD_LC_14_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIDJHD_LC_14_9_7  (
            .in0(_gnd_net_),
            .in1(N__33547),
            .in2(_gnd_net_),
            .in3(N__33535),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIFMID_LC_14_10_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIFMID_LC_14_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIFMID_LC_14_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNIFMID_LC_14_10_0  (
            .in0(_gnd_net_),
            .in1(N__33670),
            .in2(_gnd_net_),
            .in3(N__33532),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_24 ),
            .ltout(),
            .carryin(bfn_14_10_0_),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIHPJD_LC_14_10_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIHPJD_LC_14_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIHPJD_LC_14_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIHPJD_LC_14_10_1  (
            .in0(_gnd_net_),
            .in1(N__41365),
            .in2(_gnd_net_),
            .in3(N__33529),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_14_10_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_14_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_14_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_14_10_2  (
            .in0(_gnd_net_),
            .in1(N__37200),
            .in2(_gnd_net_),
            .in3(N__33526),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_14_10_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_14_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_14_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_14_10_3  (
            .in0(_gnd_net_),
            .in1(N__36702),
            .in2(_gnd_net_),
            .in3(N__33523),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_14_10_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_14_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_14_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_14_10_4  (
            .in0(_gnd_net_),
            .in1(N__37065),
            .in2(_gnd_net_),
            .in3(N__33613),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_14_10_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_14_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_14_10_5  (
            .in0(_gnd_net_),
            .in1(N__37172),
            .in2(_gnd_net_),
            .in3(N__33610),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_14_10_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_14_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_14_10_6  (
            .in0(_gnd_net_),
            .in1(N__37233),
            .in2(_gnd_net_),
            .in3(N__33607),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator1_31 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNILB5K_LC_14_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNILB5K_LC_14_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNILB5K_LC_14_10_7 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNILB5K_LC_14_10_7  (
            .in0(N__44017),
            .in1(N__36831),
            .in2(_gnd_net_),
            .in3(N__33604),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNILB5KZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIHNJ3_18_LC_14_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIHNJ3_18_LC_14_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIHNJ3_18_LC_14_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIHNJ3_18_LC_14_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41558),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_14_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_14_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_14_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_14_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34171),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_14_11_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_14_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_14_11_2  (
            .in0(N__37232),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43981),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIGMJ3_17_LC_14_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIGMJ3_17_LC_14_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIGMJ3_17_LC_14_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIGMJ3_17_LC_14_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44252),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNICJK3_22_LC_14_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNICJK3_22_LC_14_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNICJK3_22_LC_14_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNICJK3_22_LC_14_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36437),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIELK3_24_LC_14_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIELK3_24_LC_14_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIELK3_24_LC_14_11_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIELK3_24_LC_14_11_5  (
            .in0(N__40325),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_14_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_14_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_14_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_14_11_6  (
            .in0(N__37174),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43980),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_14_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_14_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_14_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_14_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34315),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_14_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_14_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_14_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_14_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34267),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_14_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_14_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_14_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34090),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBIK3_21_LC_14_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBIK3_21_LC_14_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBIK3_21_LC_14_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIBIK3_21_LC_14_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41828),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIAHK3_20_LC_14_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIAHK3_20_LC_14_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIAHK3_20_LC_14_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIAHK3_20_LC_14_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37133),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_14_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_14_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_14_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_14_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33817),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_14_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_14_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_14_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_14_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34210),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_14_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_14_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_14_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_14_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34153),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_14_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_14_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_14_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_14_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34108),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_14_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_14_13_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_14_13_0  (
            .in0(N__34234),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_14_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_14_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_14_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_14_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33784),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_14_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_14_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_14_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_14_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34297),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_14_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_14_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_14_13_3 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_14_13_3  (
            .in0(_gnd_net_),
            .in1(N__34198),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_14_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_14_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_14_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_14_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34072),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9AP1_24_LC_14_13_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9AP1_24_LC_14_13_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9AP1_24_LC_14_13_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9AP1_24_LC_14_13_5  (
            .in0(N__37801),
            .in1(N__37810),
            .in2(N__37792),
            .in3(N__37819),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_14_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_14_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_14_13_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_14_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34222),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_14_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_14_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_14_13_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_14_13_7  (
            .in0(N__34279),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_14_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_14_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_14_14_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_15_LC_14_14_0  (
            .in0(_gnd_net_),
            .in1(N__34042),
            .in2(_gnd_net_),
            .in3(N__33985),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50194),
            .ce(N__33927),
            .sr(N__49650));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_14_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_14_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_14_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_14_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33799),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_14_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_14_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_14_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_14_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34429),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_0_LC_14_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_0_LC_14_15_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_0_LC_14_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_0_LC_14_15_0  (
            .in0(_gnd_net_),
            .in1(N__34333),
            .in2(N__34357),
            .in3(N__34356),
            .lcout(\current_shift_inst.control_inputZ0Z_0 ),
            .ltout(),
            .carryin(bfn_14_15_0_),
            .carryout(\current_shift_inst.control_input_1_cry_0 ),
            .clk(N__50187),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_1_LC_14_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_1_LC_14_15_1 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_1_LC_14_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_1_LC_14_15_1  (
            .in0(_gnd_net_),
            .in1(N__34540),
            .in2(_gnd_net_),
            .in3(N__33808),
            .lcout(\current_shift_inst.control_inputZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_0 ),
            .carryout(\current_shift_inst.control_input_1_cry_1 ),
            .clk(N__50187),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_2_LC_14_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_2_LC_14_15_2 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_2_LC_14_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_2_LC_14_15_2  (
            .in0(_gnd_net_),
            .in1(N__33805),
            .in2(_gnd_net_),
            .in3(N__33793),
            .lcout(\current_shift_inst.control_inputZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_1 ),
            .carryout(\current_shift_inst.control_input_1_cry_2 ),
            .clk(N__50187),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_3_LC_14_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_3_LC_14_15_3 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_3_LC_14_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_3_LC_14_15_3  (
            .in0(_gnd_net_),
            .in1(N__33790),
            .in2(_gnd_net_),
            .in3(N__33775),
            .lcout(\current_shift_inst.control_inputZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_2 ),
            .carryout(\current_shift_inst.control_input_1_cry_3 ),
            .clk(N__50187),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_4_LC_14_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_4_LC_14_15_4 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_4_LC_14_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_4_LC_14_15_4  (
            .in0(_gnd_net_),
            .in1(N__33772),
            .in2(_gnd_net_),
            .in3(N__33751),
            .lcout(\current_shift_inst.control_inputZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_3 ),
            .carryout(\current_shift_inst.control_input_1_cry_4 ),
            .clk(N__50187),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_5_LC_14_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_5_LC_14_15_5 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_5_LC_14_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_5_LC_14_15_5  (
            .in0(_gnd_net_),
            .in1(N__47020),
            .in2(_gnd_net_),
            .in3(N__34189),
            .lcout(\current_shift_inst.control_inputZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_4 ),
            .carryout(\current_shift_inst.control_input_1_cry_5 ),
            .clk(N__50187),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_6_LC_14_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_6_LC_14_15_6 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_6_LC_14_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_6_LC_14_15_6  (
            .in0(_gnd_net_),
            .in1(N__34186),
            .in2(_gnd_net_),
            .in3(N__34174),
            .lcout(\current_shift_inst.control_inputZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_5 ),
            .carryout(\current_shift_inst.control_input_1_cry_6 ),
            .clk(N__50187),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_7_LC_14_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_7_LC_14_15_7 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_7_LC_14_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_7_LC_14_15_7  (
            .in0(_gnd_net_),
            .in1(N__46834),
            .in2(_gnd_net_),
            .in3(N__34162),
            .lcout(\current_shift_inst.control_inputZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_6 ),
            .carryout(\current_shift_inst.control_input_1_cry_7 ),
            .clk(N__50187),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_8_LC_14_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_8_LC_14_16_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_8_LC_14_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_8_LC_14_16_0  (
            .in0(_gnd_net_),
            .in1(N__34159),
            .in2(_gnd_net_),
            .in3(N__34144),
            .lcout(\current_shift_inst.control_inputZ0Z_8 ),
            .ltout(),
            .carryin(bfn_14_16_0_),
            .carryout(\current_shift_inst.control_input_1_cry_8 ),
            .clk(N__50181),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_9_LC_14_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_9_LC_14_16_1 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_9_LC_14_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_9_LC_14_16_1  (
            .in0(_gnd_net_),
            .in1(N__34141),
            .in2(_gnd_net_),
            .in3(N__34120),
            .lcout(\current_shift_inst.control_inputZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_8 ),
            .carryout(\current_shift_inst.control_input_1_cry_9 ),
            .clk(N__50181),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_10_LC_14_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_10_LC_14_16_2 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_10_LC_14_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_10_LC_14_16_2  (
            .in0(_gnd_net_),
            .in1(N__34117),
            .in2(_gnd_net_),
            .in3(N__34099),
            .lcout(\current_shift_inst.control_inputZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_9 ),
            .carryout(\current_shift_inst.control_input_1_cry_10 ),
            .clk(N__50181),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_11_LC_14_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_11_LC_14_16_3 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_11_LC_14_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_11_LC_14_16_3  (
            .in0(_gnd_net_),
            .in1(N__34096),
            .in2(_gnd_net_),
            .in3(N__34081),
            .lcout(\current_shift_inst.control_inputZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_10 ),
            .carryout(\current_shift_inst.control_input_1_cry_11 ),
            .clk(N__50181),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_12_LC_14_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_12_LC_14_16_4 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_12_LC_14_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_12_LC_14_16_4  (
            .in0(_gnd_net_),
            .in1(N__34078),
            .in2(_gnd_net_),
            .in3(N__34063),
            .lcout(\current_shift_inst.control_inputZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_11 ),
            .carryout(\current_shift_inst.control_input_1_cry_12 ),
            .clk(N__50181),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_13_LC_14_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_13_LC_14_16_5 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_13_LC_14_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_13_LC_14_16_5  (
            .in0(_gnd_net_),
            .in1(N__34324),
            .in2(_gnd_net_),
            .in3(N__34306),
            .lcout(\current_shift_inst.control_inputZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_12 ),
            .carryout(\current_shift_inst.control_input_1_cry_13 ),
            .clk(N__50181),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_14_LC_14_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_14_LC_14_16_6 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_14_LC_14_16_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_14_LC_14_16_6  (
            .in0(_gnd_net_),
            .in1(N__34303),
            .in2(_gnd_net_),
            .in3(N__34288),
            .lcout(\current_shift_inst.control_inputZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_13 ),
            .carryout(\current_shift_inst.control_input_1_cry_14 ),
            .clk(N__50181),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_15_LC_14_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_15_LC_14_16_7 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_15_LC_14_16_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_15_LC_14_16_7  (
            .in0(_gnd_net_),
            .in1(N__34285),
            .in2(_gnd_net_),
            .in3(N__34270),
            .lcout(\current_shift_inst.control_inputZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_14 ),
            .carryout(\current_shift_inst.control_input_1_cry_15 ),
            .clk(N__50181),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_16_LC_14_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_16_LC_14_17_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_16_LC_14_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_16_LC_14_17_0  (
            .in0(_gnd_net_),
            .in1(N__34573),
            .in2(_gnd_net_),
            .in3(N__34258),
            .lcout(\current_shift_inst.control_inputZ0Z_16 ),
            .ltout(),
            .carryin(bfn_14_17_0_),
            .carryout(\current_shift_inst.control_input_1_cry_16 ),
            .clk(N__50176),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_17_LC_14_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_17_LC_14_17_1 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_17_LC_14_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_17_LC_14_17_1  (
            .in0(_gnd_net_),
            .in1(N__34255),
            .in2(_gnd_net_),
            .in3(N__34237),
            .lcout(\current_shift_inst.control_inputZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_16 ),
            .carryout(\current_shift_inst.control_input_1_cry_17 ),
            .clk(N__50176),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_18_LC_14_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_18_LC_14_17_2 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_18_LC_14_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_18_LC_14_17_2  (
            .in0(_gnd_net_),
            .in1(N__34492),
            .in2(_gnd_net_),
            .in3(N__34225),
            .lcout(\current_shift_inst.control_inputZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_17 ),
            .carryout(\current_shift_inst.control_input_1_cry_18 ),
            .clk(N__50176),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_19_LC_14_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_19_LC_14_17_3 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_19_LC_14_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_19_LC_14_17_3  (
            .in0(_gnd_net_),
            .in1(N__34633),
            .in2(_gnd_net_),
            .in3(N__34213),
            .lcout(\current_shift_inst.control_inputZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_18 ),
            .carryout(\current_shift_inst.control_input_1_cry_19 ),
            .clk(N__50176),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_20_LC_14_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_20_LC_14_17_4 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_20_LC_14_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_20_LC_14_17_4  (
            .in0(_gnd_net_),
            .in1(N__34471),
            .in2(_gnd_net_),
            .in3(N__34201),
            .lcout(\current_shift_inst.control_inputZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_19 ),
            .carryout(\current_shift_inst.control_input_1_cry_20 ),
            .clk(N__50176),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_21_LC_14_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_21_LC_14_17_5 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_21_LC_14_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_21_LC_14_17_5  (
            .in0(_gnd_net_),
            .in1(N__34522),
            .in2(_gnd_net_),
            .in3(N__34447),
            .lcout(\current_shift_inst.control_inputZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_20 ),
            .carryout(\current_shift_inst.control_input_1_cry_21 ),
            .clk(N__50176),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_22_LC_14_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_22_LC_14_17_6 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_22_LC_14_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_22_LC_14_17_6  (
            .in0(_gnd_net_),
            .in1(N__34363),
            .in2(_gnd_net_),
            .in3(N__34432),
            .lcout(\current_shift_inst.control_inputZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_21 ),
            .carryout(\current_shift_inst.control_input_1_cry_22 ),
            .clk(N__50176),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_23_LC_14_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_23_LC_14_17_7 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_23_LC_14_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_23_LC_14_17_7  (
            .in0(_gnd_net_),
            .in1(N__34555),
            .in2(_gnd_net_),
            .in3(N__34420),
            .lcout(\current_shift_inst.control_inputZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_22 ),
            .carryout(\current_shift_inst.control_input_1_cry_23 ),
            .clk(N__50176),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_24_LC_14_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_24_LC_14_18_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_24_LC_14_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_24_LC_14_18_0  (
            .in0(_gnd_net_),
            .in1(N__34618),
            .in2(_gnd_net_),
            .in3(N__34405),
            .lcout(\current_shift_inst.control_inputZ0Z_24 ),
            .ltout(),
            .carryin(bfn_14_18_0_),
            .carryout(\current_shift_inst.control_input_1_cry_24 ),
            .clk(N__50171),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_25_LC_14_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_25_LC_14_18_1 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_25_LC_14_18_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.control_input_25_LC_14_18_1  (
            .in0(_gnd_net_),
            .in1(N__34402),
            .in2(_gnd_net_),
            .in3(N__34390),
            .lcout(\current_shift_inst.control_inputZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50171),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_14_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_14_18_2 .LUT_INIT=16'b0011010100110101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_14_18_2  (
            .in0(N__38629),
            .in1(N__34372),
            .in2(N__46930),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.control_input_1_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_14_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_14_18_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_14_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46901),
            .lcout(\current_shift_inst.N_1355_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_14_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_14_18_4 .LUT_INIT=16'b0101001101010011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_14_18_4  (
            .in0(N__34339),
            .in1(N__38470),
            .in2(N__46929),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.control_input_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_14_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_14_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_14_18_5 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_14_18_5  (
            .in0(N__34582),
            .in1(N__38716),
            .in2(_gnd_net_),
            .in3(N__46902),
            .lcout(\current_shift_inst.control_input_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_14_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_14_18_6 .LUT_INIT=16'b0011000000111111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_14_18_6  (
            .in0(_gnd_net_),
            .in1(N__34567),
            .in2(N__46931),
            .in3(N__39097),
            .lcout(\current_shift_inst.control_input_1_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_14_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_14_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_14_18_7 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_14_18_7  (
            .in0(N__38461),
            .in1(N__34549),
            .in2(_gnd_net_),
            .in3(N__46897),
            .lcout(\current_shift_inst.control_input_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_14_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_14_19_0 .LUT_INIT=16'b0000010110101111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_14_19_0  (
            .in0(N__46927),
            .in1(_gnd_net_),
            .in2(N__38644),
            .in3(N__34531),
            .lcout(\current_shift_inst.control_input_1_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_14_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_14_19_1 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_14_19_1  (
            .in0(N__46771),
            .in1(N__46232),
            .in2(N__47635),
            .in3(N__42907),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_14_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_14_19_2 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_14_19_2  (
            .in0(N__46231),
            .in1(N__46772),
            .in2(N__48064),
            .in3(N__45442),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI25021_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_14_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_14_19_3 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_14_19_3  (
            .in0(N__38683),
            .in1(N__34498),
            .in2(_gnd_net_),
            .in3(N__46924),
            .lcout(\current_shift_inst.control_input_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_14_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_14_19_4 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_14_19_4  (
            .in0(N__46233),
            .in1(N__46773),
            .in2(N__47953),
            .in3(N__43089),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_14_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_14_19_5 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_14_19_5  (
            .in0(N__34477),
            .in1(N__38656),
            .in2(_gnd_net_),
            .in3(N__46926),
            .lcout(\current_shift_inst.control_input_1_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_14_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_14_19_6 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_14_19_6  (
            .in0(N__46925),
            .in1(N__34639),
            .in2(_gnd_net_),
            .in3(N__38668),
            .lcout(\current_shift_inst.control_input_1_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNI9GMC2_LC_14_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNI9GMC2_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNI9GMC2_LC_14_19_7 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNI9GMC2_LC_14_19_7  (
            .in0(N__34624),
            .in1(N__39082),
            .in2(_gnd_net_),
            .in3(N__46928),
            .lcout(\current_shift_inst.control_input_1_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_14_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_14_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_14_20_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_14_20_0  (
            .in0(N__46740),
            .in1(N__48343),
            .in2(N__46342),
            .in3(N__43252),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_14_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_14_20_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_14_20_3  (
            .in0(N__46741),
            .in1(N__48427),
            .in2(N__46344),
            .in3(N__43288),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_14_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_14_20_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_14_20_4  (
            .in0(N__46739),
            .in1(N__48497),
            .in2(N__46343),
            .in3(N__43024),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_14_21_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_14_21_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_14_21_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_0_LC_14_21_0  (
            .in0(N__34823),
            .in1(N__38897),
            .in2(_gnd_net_),
            .in3(N__34594),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_14_21_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .clk(N__50158),
            .ce(N__34726),
            .sr(N__49691));
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_14_21_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_14_21_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_14_21_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_1_LC_14_21_1  (
            .in0(N__34818),
            .in1(N__38852),
            .in2(_gnd_net_),
            .in3(N__34591),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .clk(N__50158),
            .ce(N__34726),
            .sr(N__49691));
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_14_21_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_14_21_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_14_21_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_2_LC_14_21_2  (
            .in0(N__34824),
            .in1(N__35162),
            .in2(_gnd_net_),
            .in3(N__34588),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .clk(N__50158),
            .ce(N__34726),
            .sr(N__49691));
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_14_21_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_14_21_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_14_21_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_3_LC_14_21_3  (
            .in0(N__34819),
            .in1(N__35114),
            .in2(_gnd_net_),
            .in3(N__34585),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .clk(N__50158),
            .ce(N__34726),
            .sr(N__49691));
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_14_21_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_14_21_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_14_21_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_4_LC_14_21_4  (
            .in0(N__34825),
            .in1(N__35058),
            .in2(_gnd_net_),
            .in3(N__34666),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .clk(N__50158),
            .ce(N__34726),
            .sr(N__49691));
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_14_21_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_14_21_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_14_21_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_5_LC_14_21_5  (
            .in0(N__34820),
            .in1(N__35003),
            .in2(_gnd_net_),
            .in3(N__34663),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .clk(N__50158),
            .ce(N__34726),
            .sr(N__49691));
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_14_21_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_14_21_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_14_21_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_6_LC_14_21_6  (
            .in0(N__34822),
            .in1(N__34938),
            .in2(_gnd_net_),
            .in3(N__34660),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .clk(N__50158),
            .ce(N__34726),
            .sr(N__49691));
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_14_21_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_14_21_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_14_21_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_7_LC_14_21_7  (
            .in0(N__34821),
            .in1(N__35592),
            .in2(_gnd_net_),
            .in3(N__34657),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .clk(N__50158),
            .ce(N__34726),
            .sr(N__49691));
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_14_22_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_14_22_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_14_22_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_8_LC_14_22_0  (
            .in0(N__34852),
            .in1(N__35540),
            .in2(_gnd_net_),
            .in3(N__34654),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_14_22_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .clk(N__50154),
            .ce(N__34739),
            .sr(N__49700));
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_14_22_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_14_22_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_14_22_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_9_LC_14_22_1  (
            .in0(N__34870),
            .in1(N__35483),
            .in2(_gnd_net_),
            .in3(N__34651),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .clk(N__50154),
            .ce(N__34739),
            .sr(N__49700));
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_14_22_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_14_22_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_14_22_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_10_LC_14_22_2  (
            .in0(N__34849),
            .in1(N__35432),
            .in2(_gnd_net_),
            .in3(N__34648),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .clk(N__50154),
            .ce(N__34739),
            .sr(N__49700));
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_14_22_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_14_22_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_14_22_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_11_LC_14_22_3  (
            .in0(N__34867),
            .in1(N__35375),
            .in2(_gnd_net_),
            .in3(N__34645),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .clk(N__50154),
            .ce(N__34739),
            .sr(N__49700));
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_14_22_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_14_22_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_14_22_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_12_LC_14_22_4  (
            .in0(N__34850),
            .in1(N__35313),
            .in2(_gnd_net_),
            .in3(N__34642),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .clk(N__50154),
            .ce(N__34739),
            .sr(N__49700));
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_14_22_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_14_22_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_14_22_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_13_LC_14_22_5  (
            .in0(N__34868),
            .in1(N__35261),
            .in2(_gnd_net_),
            .in3(N__34693),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .clk(N__50154),
            .ce(N__34739),
            .sr(N__49700));
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_14_22_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_14_22_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_14_22_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_14_LC_14_22_6  (
            .in0(N__34851),
            .in1(N__35235),
            .in2(_gnd_net_),
            .in3(N__34690),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .clk(N__50154),
            .ce(N__34739),
            .sr(N__49700));
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_14_22_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_14_22_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_14_22_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_15_LC_14_22_7  (
            .in0(N__34869),
            .in1(N__35877),
            .in2(_gnd_net_),
            .in3(N__34687),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .clk(N__50154),
            .ce(N__34739),
            .sr(N__49700));
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_14_23_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_14_23_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_14_23_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_16_LC_14_23_0  (
            .in0(N__34863),
            .in1(N__35846),
            .in2(_gnd_net_),
            .in3(N__34684),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_14_23_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .clk(N__50150),
            .ce(N__34741),
            .sr(N__49704));
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_14_23_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_14_23_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_14_23_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_17_LC_14_23_1  (
            .in0(N__34853),
            .in1(N__35813),
            .in2(_gnd_net_),
            .in3(N__34681),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .clk(N__50150),
            .ce(N__34741),
            .sr(N__49704));
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_14_23_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_14_23_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_14_23_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_18_LC_14_23_2  (
            .in0(N__34864),
            .in1(N__35774),
            .in2(_gnd_net_),
            .in3(N__34678),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .clk(N__50150),
            .ce(N__34741),
            .sr(N__49704));
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_14_23_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_14_23_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_14_23_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_19_LC_14_23_3  (
            .in0(N__34854),
            .in1(N__35738),
            .in2(_gnd_net_),
            .in3(N__34675),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .clk(N__50150),
            .ce(N__34741),
            .sr(N__49704));
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_14_23_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_14_23_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_14_23_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_20_LC_14_23_4  (
            .in0(N__34865),
            .in1(N__35694),
            .in2(_gnd_net_),
            .in3(N__34672),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .clk(N__50150),
            .ce(N__34741),
            .sr(N__49704));
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_14_23_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_14_23_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_14_23_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_21_LC_14_23_5  (
            .in0(N__34855),
            .in1(N__35663),
            .in2(_gnd_net_),
            .in3(N__34669),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .clk(N__50150),
            .ce(N__34741),
            .sr(N__49704));
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_14_23_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_14_23_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_14_23_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_22_LC_14_23_6  (
            .in0(N__34866),
            .in1(N__35631),
            .in2(_gnd_net_),
            .in3(N__34891),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .clk(N__50150),
            .ce(N__34741),
            .sr(N__49704));
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_14_23_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_14_23_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_14_23_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_23_LC_14_23_7  (
            .in0(N__34856),
            .in1(N__36126),
            .in2(_gnd_net_),
            .in3(N__34888),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .clk(N__50150),
            .ce(N__34741),
            .sr(N__49704));
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_14_24_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_14_24_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_14_24_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_24_LC_14_24_0  (
            .in0(N__34857),
            .in1(N__36089),
            .in2(_gnd_net_),
            .in3(N__34885),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_14_24_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .clk(N__50145),
            .ce(N__34740),
            .sr(N__49709));
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_14_24_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_14_24_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_14_24_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_25_LC_14_24_1  (
            .in0(N__34861),
            .in1(N__36050),
            .in2(_gnd_net_),
            .in3(N__34882),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .clk(N__50145),
            .ce(N__34740),
            .sr(N__49709));
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_14_24_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_14_24_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_14_24_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_26_LC_14_24_2  (
            .in0(N__34858),
            .in1(N__36020),
            .in2(_gnd_net_),
            .in3(N__34879),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .clk(N__50145),
            .ce(N__34740),
            .sr(N__49709));
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_14_24_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_14_24_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_14_24_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_27_LC_14_24_3  (
            .in0(N__34862),
            .in1(N__35966),
            .in2(_gnd_net_),
            .in3(N__34876),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .clk(N__50145),
            .ce(N__34740),
            .sr(N__49709));
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_14_24_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_14_24_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_14_24_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_28_LC_14_24_4  (
            .in0(N__34859),
            .in1(N__35994),
            .in2(_gnd_net_),
            .in3(N__34873),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ),
            .clk(N__50145),
            .ce(N__34740),
            .sr(N__49709));
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_14_24_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_14_24_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_14_24_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_29_LC_14_24_5  (
            .in0(N__35943),
            .in1(N__34860),
            .in2(_gnd_net_),
            .in3(N__34744),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50145),
            .ce(N__34740),
            .sr(N__49709));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOKRB1_10_LC_14_25_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOKRB1_10_LC_14_25_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOKRB1_10_LC_14_25_4 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOKRB1_10_LC_14_25_4  (
            .in0(N__35564),
            .in1(N__35202),
            .in2(N__38962),
            .in3(N__38831),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRMG72_7_LC_14_25_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRMG72_7_LC_14_25_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRMG72_7_LC_14_25_5 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRMG72_7_LC_14_25_5  (
            .in0(_gnd_net_),
            .in1(N__34972),
            .in2(N__35218),
            .in3(N__35040),
            .lcout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_14_26_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_14_26_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_14_26_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_14_26_0  (
            .in0(_gnd_net_),
            .in1(N__38904),
            .in2(N__35167),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.elapsed_time_hc_3 ),
            .ltout(),
            .carryin(bfn_14_26_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__50137),
            .ce(N__38811),
            .sr(N__49726));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_14_26_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_14_26_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_14_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_14_26_1  (
            .in0(_gnd_net_),
            .in1(N__38859),
            .in2(N__35119),
            .in3(N__35170),
            .lcout(\delay_measurement_inst.elapsed_time_hc_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__50137),
            .ce(N__38811),
            .sr(N__49726));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_14_26_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_14_26_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_14_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_14_26_2  (
            .in0(_gnd_net_),
            .in1(N__35166),
            .in2(N__35070),
            .in3(N__35122),
            .lcout(\delay_measurement_inst.elapsed_time_hc_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__50137),
            .ce(N__38811),
            .sr(N__49726));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_14_26_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_14_26_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_14_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_14_26_3  (
            .in0(_gnd_net_),
            .in1(N__35118),
            .in2(N__35014),
            .in3(N__35074),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__50137),
            .ce(N__38811),
            .sr(N__49726));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_14_26_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_14_26_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_14_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_14_26_4  (
            .in0(_gnd_net_),
            .in1(N__34944),
            .in2(N__35071),
            .in3(N__35017),
            .lcout(\delay_measurement_inst.elapsed_time_hc_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__50137),
            .ce(N__38811),
            .sr(N__49726));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_14_26_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_14_26_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_14_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_14_26_5  (
            .in0(_gnd_net_),
            .in1(N__35013),
            .in2(N__35604),
            .in3(N__34948),
            .lcout(\delay_measurement_inst.elapsed_time_hc_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__50137),
            .ce(N__38811),
            .sr(N__49726));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_14_26_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_14_26_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_14_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_14_26_6  (
            .in0(_gnd_net_),
            .in1(N__34945),
            .in2(N__35545),
            .in3(N__34894),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__50137),
            .ce(N__38811),
            .sr(N__49726));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_14_26_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_14_26_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_14_26_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_14_26_7  (
            .in0(_gnd_net_),
            .in1(N__35490),
            .in2(N__35605),
            .in3(N__35548),
            .lcout(\delay_measurement_inst.elapsed_time_hc_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__50137),
            .ce(N__38811),
            .sr(N__49726));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_14_27_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_14_27_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_14_27_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_14_27_0  (
            .in0(_gnd_net_),
            .in1(N__35544),
            .in2(N__35437),
            .in3(N__35497),
            .lcout(\delay_measurement_inst.elapsed_time_hc_11 ),
            .ltout(),
            .carryin(bfn_14_27_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__50134),
            .ce(N__38810),
            .sr(N__49731));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_14_27_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_14_27_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_14_27_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_14_27_1  (
            .in0(_gnd_net_),
            .in1(N__35494),
            .in2(N__35380),
            .in3(N__35440),
            .lcout(\delay_measurement_inst.elapsed_time_hc_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__50134),
            .ce(N__38810),
            .sr(N__49731));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_14_27_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_14_27_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_14_27_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_14_27_2  (
            .in0(_gnd_net_),
            .in1(N__35436),
            .in2(N__35325),
            .in3(N__35383),
            .lcout(\delay_measurement_inst.elapsed_time_hc_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__50134),
            .ce(N__38810),
            .sr(N__49731));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_14_27_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_14_27_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_14_27_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_14_27_3  (
            .in0(_gnd_net_),
            .in1(N__35379),
            .in2(N__35268),
            .in3(N__35329),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__50134),
            .ce(N__38810),
            .sr(N__49731));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_14_27_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_14_27_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_14_27_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_14_27_4  (
            .in0(_gnd_net_),
            .in1(N__35241),
            .in2(N__35326),
            .in3(N__35272),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__50134),
            .ce(N__38810),
            .sr(N__49731));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_14_27_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_14_27_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_14_27_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_14_27_5  (
            .in0(_gnd_net_),
            .in1(N__35883),
            .in2(N__35269),
            .in3(N__35245),
            .lcout(\delay_measurement_inst.elapsed_time_hc_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__50134),
            .ce(N__38810),
            .sr(N__49731));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_14_27_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_14_27_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_14_27_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_14_27_6  (
            .in0(_gnd_net_),
            .in1(N__35242),
            .in2(N__35859),
            .in3(N__35221),
            .lcout(\delay_measurement_inst.elapsed_time_hc_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__50134),
            .ce(N__38810),
            .sr(N__49731));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_14_27_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_14_27_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_14_27_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_14_27_7  (
            .in0(_gnd_net_),
            .in1(N__35884),
            .in2(N__35826),
            .in3(N__35863),
            .lcout(\delay_measurement_inst.elapsed_time_hc_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__50134),
            .ce(N__38810),
            .sr(N__49731));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_14_28_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_14_28_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_14_28_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_14_28_0  (
            .in0(_gnd_net_),
            .in1(N__35860),
            .in2(N__35779),
            .in3(N__35830),
            .lcout(\delay_measurement_inst.elapsed_time_hc_19 ),
            .ltout(),
            .carryin(bfn_14_28_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__50132),
            .ce(N__38809),
            .sr(N__49736));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_14_28_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_14_28_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_14_28_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_14_28_1  (
            .in0(_gnd_net_),
            .in1(N__35827),
            .in2(N__35743),
            .in3(N__35782),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__50132),
            .ce(N__38809),
            .sr(N__49736));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_14_28_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_14_28_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_14_28_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_14_28_2  (
            .in0(_gnd_net_),
            .in1(N__35778),
            .in2(N__35706),
            .in3(N__35746),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__50132),
            .ce(N__38809),
            .sr(N__49736));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_14_28_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_14_28_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_14_28_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_14_28_3  (
            .in0(_gnd_net_),
            .in1(N__35742),
            .in2(N__35670),
            .in3(N__35710),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__50132),
            .ce(N__38809),
            .sr(N__49736));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_14_28_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_14_28_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_14_28_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_14_28_4  (
            .in0(_gnd_net_),
            .in1(N__35637),
            .in2(N__35707),
            .in3(N__35674),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__50132),
            .ce(N__38809),
            .sr(N__49736));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_14_28_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_14_28_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_14_28_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_14_28_5  (
            .in0(_gnd_net_),
            .in1(N__36132),
            .in2(N__35671),
            .in3(N__35641),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__50132),
            .ce(N__38809),
            .sr(N__49736));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_14_28_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_14_28_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_14_28_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_14_28_6  (
            .in0(_gnd_net_),
            .in1(N__35638),
            .in2(N__36100),
            .in3(N__35608),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__50132),
            .ce(N__38809),
            .sr(N__49736));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_14_28_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_14_28_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_14_28_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_14_28_7  (
            .in0(_gnd_net_),
            .in1(N__36133),
            .in2(N__36063),
            .in3(N__36103),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__50132),
            .ce(N__38809),
            .sr(N__49736));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_14_29_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_14_29_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_14_29_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_14_29_0  (
            .in0(_gnd_net_),
            .in1(N__36099),
            .in2(N__36025),
            .in3(N__36067),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ),
            .ltout(),
            .carryin(bfn_14_29_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__50130),
            .ce(N__38808),
            .sr(N__49738));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_14_29_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_14_29_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_14_29_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_14_29_1  (
            .in0(_gnd_net_),
            .in1(N__36064),
            .in2(N__35971),
            .in3(N__36028),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__50130),
            .ce(N__38808),
            .sr(N__49738));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_14_29_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_14_29_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_14_29_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_14_29_2  (
            .in0(_gnd_net_),
            .in1(N__36024),
            .in2(N__36001),
            .in3(N__35974),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__50130),
            .ce(N__38808),
            .sr(N__49738));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_14_29_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_14_29_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_14_29_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_14_29_3  (
            .in0(_gnd_net_),
            .in1(N__35970),
            .in2(N__35947),
            .in3(N__35920),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__50130),
            .ce(N__38808),
            .sr(N__49738));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_14_29_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_14_29_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_14_29_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_14_29_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35917),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50130),
            .ce(N__38808),
            .sr(N__49738));
    defparam SB_DFF_inst_DELAY_TR1_LC_15_2_1.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_TR1_LC_15_2_1.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_TR1_LC_15_2_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_DELAY_TR1_LC_15_2_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35899),
            .lcout(delay_tr_d1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50271),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_DELAY_TR2_LC_15_2_2.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_TR2_LC_15_2_2.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_TR2_LC_15_2_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_DELAY_TR2_LC_15_2_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35890),
            .lcout(delay_tr_d2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50271),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.stop_timer_tr_LC_15_2_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_tr_LC_15_2_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.stop_timer_tr_LC_15_2_6 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \delay_measurement_inst.stop_timer_tr_LC_15_2_6  (
            .in0(N__39187),
            .in1(N__39208),
            .in2(N__49791),
            .in3(N__39169),
            .lcout(\delay_measurement_inst.stop_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50271),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.tr_state_0_LC_15_3_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.tr_state_0_LC_15_3_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.tr_state_0_LC_15_3_0 .LUT_INIT=16'b1100110001100110;
    LogicCell40 \delay_measurement_inst.tr_state_0_LC_15_3_0  (
            .in0(N__39188),
            .in1(N__39206),
            .in2(_gnd_net_),
            .in3(N__39168),
            .lcout(\delay_measurement_inst.tr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50267),
            .ce(N__36415),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNITAU01_13_LC_15_6_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNITAU01_13_LC_15_6_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNITAU01_13_LC_15_6_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNITAU01_13_LC_15_6_0  (
            .in0(N__44079),
            .in1(N__36322),
            .in2(N__43588),
            .in3(N__36286),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNITAU01Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_15_6_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_15_6_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_15_6_2 .LUT_INIT=16'b0101010100000111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_9_LC_15_6_2  (
            .in0(N__39505),
            .in1(N__45124),
            .in2(N__44933),
            .in3(N__45338),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50252),
            .ce(),
            .sr(N__49612));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIC46U_6_LC_15_7_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIC46U_6_LC_15_7_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIC46U_6_LC_15_7_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIC46U_6_LC_15_7_1  (
            .in0(N__44051),
            .in1(N__36276),
            .in2(N__39392),
            .in3(N__36247),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIC46UZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI8V4U_5_LC_15_7_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI8V4U_5_LC_15_7_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI8V4U_5_LC_15_7_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI8V4U_5_LC_15_7_2  (
            .in0(N__44050),
            .in1(N__36240),
            .in2(N__36532),
            .in3(N__36211),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNI8V4UZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI4Q3U_4_LC_15_7_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI4Q3U_4_LC_15_7_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI4Q3U_4_LC_15_7_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI4Q3U_4_LC_15_7_4  (
            .in0(N__44049),
            .in1(N__36204),
            .in2(N__39286),
            .in3(N__36175),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNI4Q3UZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_15_7_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_15_7_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_15_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_15_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43569),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIKE8U_8_LC_15_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIKE8U_8_LC_15_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIKE8U_8_LC_15_8_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIKE8U_8_LC_15_8_0  (
            .in0(N__44053),
            .in1(N__36168),
            .in2(N__39361),
            .in3(N__36139),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIKE8UZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_15_8_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_15_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_15_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_15_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43528),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIG97U_7_LC_15_8_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIG97U_7_LC_15_8_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIG97U_7_LC_15_8_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIG97U_7_LC_15_8_2  (
            .in0(N__44052),
            .in1(N__36682),
            .in2(N__40881),
            .in3(N__36655),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIG97UZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIOJ9U_9_LC_15_8_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIOJ9U_9_LC_15_8_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIOJ9U_9_LC_15_8_3 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIOJ9U_9_LC_15_8_3  (
            .in0(N__43468),
            .in1(N__44054),
            .in2(N__36649),
            .in3(N__36616),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIOJ9UZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIA1B41_10_LC_15_8_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIA1B41_10_LC_15_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIA1B41_10_LC_15_8_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIA1B41_10_LC_15_8_4  (
            .in0(N__44055),
            .in1(N__36609),
            .in2(N__43536),
            .in3(N__36580),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIA1B41Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIP5T01_12_LC_15_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIP5T01_12_LC_15_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIP5T01_12_LC_15_8_5 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIP5T01_12_LC_15_8_5  (
            .in0(N__43625),
            .in1(N__44056),
            .in2(N__36574),
            .in3(N__36538),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIP5T01Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_15_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_15_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_15_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_15_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41718),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_15_8_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_15_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_15_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_15_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36531),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIL0S01_11_LC_15_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIL0S01_11_LC_15_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIL0S01_11_LC_15_9_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIL0S01_11_LC_15_9_0  (
            .in0(N__36486),
            .in1(N__43983),
            .in2(N__44203),
            .in3(N__36457),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIL0S01Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIDGBQ_22_LC_15_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIDGBQ_22_LC_15_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIDGBQ_22_LC_15_9_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIDGBQ_22_LC_15_9_1  (
            .in0(N__43987),
            .in1(N__36450),
            .in2(N__40207),
            .in3(N__36421),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIDGBQZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIGNK3_0_26_LC_15_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIGNK3_0_26_LC_15_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIGNK3_0_26_LC_15_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIGNK3_0_26_LC_15_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43982),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_i_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIS2EP_19_LC_15_9_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIS2EP_19_LC_15_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIS2EP_19_LC_15_9_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIS2EP_19_LC_15_9_3  (
            .in0(N__43986),
            .in1(N__36952),
            .in2(N__36928),
            .in3(N__36877),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIS2EPZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNICE9P_15_LC_15_9_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNICE9P_15_LC_15_9_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNICE9P_15_LC_15_9_4 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNICE9P_15_LC_15_9_4  (
            .in0(N__41728),
            .in1(N__43984),
            .in2(N__36871),
            .in3(N__36861),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNICE9PZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_15_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_15_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_15_9_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_15_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36827),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_15_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_15_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_15_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_15_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37115),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIGJAP_16_LC_15_9_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIGJAP_16_LC_15_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIGJAP_16_LC_15_9_7 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIGJAP_16_LC_15_9_7  (
            .in0(N__43985),
            .in1(N__36778),
            .in2(N__41674),
            .in3(N__36771),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIGJAPZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIHLCQ_23_LC_15_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIHLCQ_23_LC_15_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIHLCQ_23_LC_15_10_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIHLCQ_23_LC_15_10_0  (
            .in0(N__44068),
            .in1(N__36738),
            .in2(N__40150),
            .in3(N__36709),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIHLCQZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_15_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_15_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_15_10_1  (
            .in0(N__36703),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44066),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ),
            .ltout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_27_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIMG8J_LC_15_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIMG8J_LC_15_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIMG8J_LC_15_10_2 .LUT_INIT=16'b0101111111110101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIMG8J_LC_15_10_2  (
            .in0(N__44070),
            .in1(N__44453),
            .in2(N__36691),
            .in3(N__36688),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIMG8JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNISPBJ_LC_15_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNISPBJ_LC_15_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNISPBJ_LC_15_10_3 .LUT_INIT=16'b0111011110111011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNISPBJ_LC_15_10_3  (
            .in0(N__37234),
            .in1(N__44073),
            .in2(N__44651),
            .in3(N__37210),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNISPBJZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIKD7J_LC_15_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIKD7J_LC_15_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIKD7J_LC_15_10_4 .LUT_INIT=16'b0111011111011101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIKD7J_LC_15_10_4  (
            .in0(N__44069),
            .in1(N__37204),
            .in2(N__39492),
            .in3(N__37180),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIKD7JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNIQMAJ_LC_15_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNIQMAJ_LC_15_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNIQMAJ_LC_15_10_5 .LUT_INIT=16'b0111101101111011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNIQMAJ_LC_15_10_5  (
            .in0(N__37173),
            .in1(N__44072),
            .in2(N__37156),
            .in3(N__41338),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNIQMAJZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIENGP_20_LC_15_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIENGP_20_LC_15_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIENGP_20_LC_15_10_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIENGP_20_LC_15_10_6  (
            .in0(N__44067),
            .in1(N__37146),
            .in2(N__37120),
            .in3(N__37075),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIENGPZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIOJ9J_LC_15_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIOJ9J_LC_15_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIOJ9J_LC_15_10_7 .LUT_INIT=16'b0111011110111011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIOJ9J_LC_15_10_7  (
            .in0(N__37069),
            .in1(N__44071),
            .in2(N__44581),
            .in3(N__37045),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNIOJ9JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_15_11_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_15_11_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_15_11_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_15_11_0  (
            .in0(_gnd_net_),
            .in1(N__50328),
            .in2(N__41610),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.elapsed_time_tr_3 ),
            .ltout(),
            .carryin(bfn_15_11_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__50222),
            .ce(N__49811),
            .sr(N__49625));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_15_11_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_15_11_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_15_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_15_11_1  (
            .in0(_gnd_net_),
            .in1(N__44332),
            .in2(N__42090),
            .in3(N__36976),
            .lcout(\delay_measurement_inst.elapsed_time_tr_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__50222),
            .ce(N__49811),
            .sr(N__49625));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_15_11_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_15_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_15_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_15_11_2  (
            .in0(_gnd_net_),
            .in1(N__42063),
            .in2(N__41611),
            .in3(N__36955),
            .lcout(\delay_measurement_inst.elapsed_time_tr_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__50222),
            .ce(N__49811),
            .sr(N__49625));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_15_11_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_15_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_15_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_15_11_3  (
            .in0(_gnd_net_),
            .in1(N__42042),
            .in2(N__42091),
            .in3(N__37435),
            .lcout(\delay_measurement_inst.delay_tr_reg3lto6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__50222),
            .ce(N__49811),
            .sr(N__49625));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_15_11_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_15_11_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_15_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_15_11_4  (
            .in0(_gnd_net_),
            .in1(N__42064),
            .in2(N__42018),
            .in3(N__37408),
            .lcout(\delay_measurement_inst.elapsed_time_tr_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__50222),
            .ce(N__49811),
            .sr(N__49625));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_15_11_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_15_11_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_15_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_15_11_5  (
            .in0(_gnd_net_),
            .in1(N__42043),
            .in2(N__41991),
            .in3(N__37384),
            .lcout(\delay_measurement_inst.elapsed_time_tr_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__50222),
            .ce(N__49811),
            .sr(N__49625));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_15_11_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_15_11_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_15_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_15_11_6  (
            .in0(_gnd_net_),
            .in1(N__41965),
            .in2(N__42019),
            .in3(N__37330),
            .lcout(\delay_measurement_inst.delay_tr_reg3lto9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__50222),
            .ce(N__49811),
            .sr(N__49625));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_15_11_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_15_11_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_15_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_15_11_7  (
            .in0(_gnd_net_),
            .in1(N__41938),
            .in2(N__41992),
            .in3(N__37306),
            .lcout(\delay_measurement_inst.elapsed_time_tr_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__50222),
            .ce(N__49811),
            .sr(N__49625));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_15_12_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_15_12_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_15_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_15_12_0  (
            .in0(_gnd_net_),
            .in1(N__41964),
            .in2(N__41907),
            .in3(N__37285),
            .lcout(\delay_measurement_inst.elapsed_time_tr_11 ),
            .ltout(),
            .carryin(bfn_15_12_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__50212),
            .ce(N__49812),
            .sr(N__49630));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_15_12_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_15_12_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_15_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_15_12_1  (
            .in0(_gnd_net_),
            .in1(N__41937),
            .in2(N__41880),
            .in3(N__37261),
            .lcout(\delay_measurement_inst.elapsed_time_tr_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__50212),
            .ce(N__49812),
            .sr(N__49630));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_15_12_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_15_12_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_15_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_15_12_2  (
            .in0(_gnd_net_),
            .in1(N__42300),
            .in2(N__41908),
            .in3(N__37237),
            .lcout(\delay_measurement_inst.elapsed_time_tr_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__50212),
            .ce(N__49812),
            .sr(N__49630));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_15_12_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_15_12_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_15_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_15_12_3  (
            .in0(_gnd_net_),
            .in1(N__42276),
            .in2(N__41881),
            .in3(N__37702),
            .lcout(\delay_measurement_inst.delay_tr_reg3lto14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__50212),
            .ce(N__49812),
            .sr(N__49630));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_15_12_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_15_12_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_15_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_15_12_4  (
            .in0(_gnd_net_),
            .in1(N__42301),
            .in2(N__42255),
            .in3(N__37654),
            .lcout(\delay_measurement_inst.delay_tr_reg3lto15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__50212),
            .ce(N__49812),
            .sr(N__49630));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_15_12_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_15_12_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_15_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_15_12_5  (
            .in0(_gnd_net_),
            .in1(N__42277),
            .in2(N__42228),
            .in3(N__37618),
            .lcout(\delay_measurement_inst.elapsed_time_tr_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__50212),
            .ce(N__49812),
            .sr(N__49630));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_15_12_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_15_12_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_15_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_15_12_6  (
            .in0(_gnd_net_),
            .in1(N__42202),
            .in2(N__42256),
            .in3(N__37576),
            .lcout(\delay_measurement_inst.elapsed_time_tr_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__50212),
            .ce(N__49812),
            .sr(N__49630));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_15_12_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_15_12_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_15_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_15_12_7  (
            .in0(_gnd_net_),
            .in1(N__42172),
            .in2(N__42229),
            .in3(N__37537),
            .lcout(\delay_measurement_inst.elapsed_time_tr_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__50212),
            .ce(N__49812),
            .sr(N__49630));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_15_13_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_15_13_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_15_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_15_13_0  (
            .in0(_gnd_net_),
            .in1(N__42201),
            .in2(N__42144),
            .in3(N__37498),
            .lcout(\delay_measurement_inst.elapsed_time_tr_19 ),
            .ltout(),
            .carryin(bfn_15_13_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__50208),
            .ce(N__49813),
            .sr(N__49639));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_15_13_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_15_13_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_15_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_15_13_1  (
            .in0(_gnd_net_),
            .in1(N__42171),
            .in2(N__42117),
            .in3(N__37495),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__50208),
            .ce(N__49813),
            .sr(N__49639));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_15_13_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_15_13_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_15_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_15_13_2  (
            .in0(_gnd_net_),
            .in1(N__42525),
            .in2(N__42145),
            .in3(N__37492),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__50208),
            .ce(N__49813),
            .sr(N__49639));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_15_13_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_15_13_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_15_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_15_13_3  (
            .in0(_gnd_net_),
            .in1(N__42504),
            .in2(N__42118),
            .in3(N__37489),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__50208),
            .ce(N__49813),
            .sr(N__49639));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_15_13_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_15_13_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_15_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_15_13_4  (
            .in0(_gnd_net_),
            .in1(N__42526),
            .in2(N__42483),
            .in3(N__37822),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__50208),
            .ce(N__49813),
            .sr(N__49639));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_15_13_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_15_13_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_15_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_15_13_5  (
            .in0(_gnd_net_),
            .in1(N__42505),
            .in2(N__42456),
            .in3(N__37813),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__50208),
            .ce(N__49813),
            .sr(N__49639));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_15_13_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_15_13_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_15_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_15_13_6  (
            .in0(_gnd_net_),
            .in1(N__42430),
            .in2(N__42484),
            .in3(N__37804),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__50208),
            .ce(N__49813),
            .sr(N__49639));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_15_13_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_15_13_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_15_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_15_13_7  (
            .in0(_gnd_net_),
            .in1(N__42403),
            .in2(N__42457),
            .in3(N__37795),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__50208),
            .ce(N__49813),
            .sr(N__49639));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_15_14_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_15_14_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_15_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_15_14_0  (
            .in0(_gnd_net_),
            .in1(N__42429),
            .in2(N__42372),
            .in3(N__37783),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ),
            .ltout(),
            .carryin(bfn_15_14_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__50202),
            .ce(N__49814),
            .sr(N__49645));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_15_14_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_15_14_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_15_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_15_14_1  (
            .in0(_gnd_net_),
            .in1(N__42402),
            .in2(N__42345),
            .in3(N__37771),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__50202),
            .ce(N__49814),
            .sr(N__49645));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_15_14_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_15_14_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_15_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_15_14_2  (
            .in0(_gnd_net_),
            .in1(N__42319),
            .in2(N__42373),
            .in3(N__37759),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__50202),
            .ce(N__49814),
            .sr(N__49645));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_15_14_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_15_14_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_15_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_15_14_3  (
            .in0(_gnd_net_),
            .in1(N__42655),
            .in2(N__42346),
            .in3(N__37741),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__50202),
            .ce(N__49814),
            .sr(N__49645));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_15_14_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_15_14_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_15_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_15_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37939),
            .lcout(\delay_measurement_inst.elapsed_time_tr_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50202),
            .ce(N__49814),
            .sr(N__49645));
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_15_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_15_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_LC_15_15_0  (
            .in0(_gnd_net_),
            .in1(N__45360),
            .in2(N__37852),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_15_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_15_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_15_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_15_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_LC_15_15_1  (
            .in0(_gnd_net_),
            .in1(N__40357),
            .in2(N__38380),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_0 ),
            .carryout(\current_shift_inst.un10_control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_15_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_15_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_15_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_LC_15_15_2  (
            .in0(_gnd_net_),
            .in1(N__47125),
            .in2(N__38384),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_1 ),
            .carryout(\current_shift_inst.un10_control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_15_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_15_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_15_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_LC_15_15_3  (
            .in0(_gnd_net_),
            .in1(N__40465),
            .in2(N__38381),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_2 ),
            .carryout(\current_shift_inst.un10_control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_15_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_15_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_15_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_LC_15_15_4  (
            .in0(_gnd_net_),
            .in1(N__38326),
            .in2(N__40447),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_3 ),
            .carryout(\current_shift_inst.un10_control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_15_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_15_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_15_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_LC_15_15_5  (
            .in0(_gnd_net_),
            .in1(N__40453),
            .in2(N__38382),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_4 ),
            .carryout(\current_shift_inst.un10_control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_15_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_15_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_15_15_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_LC_15_15_6  (
            .in0(_gnd_net_),
            .in1(N__45469),
            .in2(N__38385),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_5 ),
            .carryout(\current_shift_inst.un10_control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_15_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_15_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_15_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_LC_15_15_7  (
            .in0(_gnd_net_),
            .in1(N__40459),
            .in2(N__38383),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_6 ),
            .carryout(\current_shift_inst.un10_control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_15_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_15_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_15_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_LC_15_16_0  (
            .in0(_gnd_net_),
            .in1(N__40525),
            .in2(N__38375),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_16_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_15_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_15_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_15_16_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_LC_15_16_1  (
            .in0(_gnd_net_),
            .in1(N__40489),
            .in2(N__38379),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_8 ),
            .carryout(\current_shift_inst.un10_control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_15_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_15_16_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_LC_15_16_2  (
            .in0(_gnd_net_),
            .in1(N__40495),
            .in2(N__38372),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_9 ),
            .carryout(\current_shift_inst.un10_control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_15_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_15_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_15_16_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_LC_15_16_3  (
            .in0(_gnd_net_),
            .in1(N__40507),
            .in2(N__38376),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_10 ),
            .carryout(\current_shift_inst.un10_control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_15_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_15_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_15_16_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_LC_15_16_4  (
            .in0(_gnd_net_),
            .in1(N__40519),
            .in2(N__38373),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_11 ),
            .carryout(\current_shift_inst.un10_control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_15_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_15_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_15_16_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_LC_15_16_5  (
            .in0(_gnd_net_),
            .in1(N__40531),
            .in2(N__38377),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_12 ),
            .carryout(\current_shift_inst.un10_control_input_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_15_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_15_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_15_16_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_LC_15_16_6  (
            .in0(_gnd_net_),
            .in1(N__40501),
            .in2(N__38374),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_13 ),
            .carryout(\current_shift_inst.un10_control_input_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_15_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_15_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_15_16_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_LC_15_16_7  (
            .in0(_gnd_net_),
            .in1(N__40513),
            .in2(N__38378),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_14 ),
            .carryout(\current_shift_inst.un10_control_input_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_15_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_15_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_LC_15_17_0  (
            .in0(_gnd_net_),
            .in1(N__40609),
            .in2(N__38289),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_17_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_15_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_15_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_LC_15_17_1  (
            .in0(_gnd_net_),
            .in1(N__40603),
            .in2(N__38293),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_16 ),
            .carryout(\current_shift_inst.un10_control_input_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_15_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_15_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_LC_15_17_2  (
            .in0(_gnd_net_),
            .in1(N__45409),
            .in2(N__38290),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_17 ),
            .carryout(\current_shift_inst.un10_control_input_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_15_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_15_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_LC_15_17_3  (
            .in0(_gnd_net_),
            .in1(N__40483),
            .in2(N__38294),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_18 ),
            .carryout(\current_shift_inst.un10_control_input_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_15_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_15_17_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_LC_15_17_4  (
            .in0(_gnd_net_),
            .in1(N__40654),
            .in2(N__38291),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_19 ),
            .carryout(\current_shift_inst.un10_control_input_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_15_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_15_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_LC_15_17_5  (
            .in0(_gnd_net_),
            .in1(N__38200),
            .in2(N__40648),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_20 ),
            .carryout(\current_shift_inst.un10_control_input_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_15_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_15_17_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_LC_15_17_6  (
            .in0(_gnd_net_),
            .in1(N__40597),
            .in2(N__38292),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_21 ),
            .carryout(\current_shift_inst.un10_control_input_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_15_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_15_17_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_LC_15_17_7  (
            .in0(_gnd_net_),
            .in1(N__40567),
            .in2(N__38295),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_22 ),
            .carryout(\current_shift_inst.un10_control_input_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_15_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_15_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_LC_15_18_0  (
            .in0(_gnd_net_),
            .in1(N__40552),
            .in2(N__38280),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_18_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_15_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_15_18_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_LC_15_18_1  (
            .in0(_gnd_net_),
            .in1(N__40666),
            .in2(N__38284),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_24 ),
            .carryout(\current_shift_inst.un10_control_input_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_15_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_15_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_LC_15_18_2  (
            .in0(_gnd_net_),
            .in1(N__40540),
            .in2(N__38281),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_25 ),
            .carryout(\current_shift_inst.un10_control_input_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_15_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_15_18_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_LC_15_18_3  (
            .in0(_gnd_net_),
            .in1(N__40546),
            .in2(N__38285),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_26 ),
            .carryout(\current_shift_inst.un10_control_input_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_15_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_15_18_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_LC_15_18_4  (
            .in0(_gnd_net_),
            .in1(N__40615),
            .in2(N__38282),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_27 ),
            .carryout(\current_shift_inst.un10_control_input_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_15_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_15_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_15_18_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_LC_15_18_5  (
            .in0(_gnd_net_),
            .in1(N__40729),
            .in2(N__38286),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_28 ),
            .carryout(\current_shift_inst.un10_control_input_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_15_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_15_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_15_18_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_LC_15_18_6  (
            .in0(_gnd_net_),
            .in1(N__43186),
            .in2(N__38283),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_29 ),
            .carryout(\current_shift_inst.un10_control_input_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_15_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_15_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_15_18_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_15_18_7  (
            .in0(_gnd_net_),
            .in1(N__46749),
            .in2(_gnd_net_),
            .in3(N__37996),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_15_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_15_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_LC_15_19_0  (
            .in0(_gnd_net_),
            .in1(N__37993),
            .in2(N__37974),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_19_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_15_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_15_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_LC_15_19_1  (
            .in0(_gnd_net_),
            .in1(N__40387),
            .in2(N__40425),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_15_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_15_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_LC_15_19_2  (
            .in0(_gnd_net_),
            .in1(N__37951),
            .in2(N__46255),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_LC_15_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_LC_15_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s1_c_LC_15_19_3  (
            .in0(_gnd_net_),
            .in1(N__40477),
            .in2(N__46258),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_LC_15_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_LC_15_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_LC_15_19_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s1_c_LC_15_19_4  (
            .in0(_gnd_net_),
            .in1(N__40717),
            .in2(N__46256),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_LC_15_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_LC_15_19_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s1_c_LC_15_19_5  (
            .in0(_gnd_net_),
            .in1(N__40660),
            .in2(N__46259),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_15_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_15_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_15_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_15_19_6  (
            .in0(_gnd_net_),
            .in1(N__47062),
            .in2(N__46257),
            .in3(N__38464),
            .lcout(\current_shift_inst.un38_control_input_0_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_15_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_15_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_15_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_15_19_7  (
            .in0(_gnd_net_),
            .in1(N__47383),
            .in2(N__46260),
            .in3(N__38452),
            .lcout(\current_shift_inst.un38_control_input_0_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_15_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_15_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_15_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_15_20_0  (
            .in0(_gnd_net_),
            .in1(N__40627),
            .in2(N__46325),
            .in3(N__38437),
            .lcout(\current_shift_inst.un38_control_input_0_s1_8 ),
            .ltout(),
            .carryin(bfn_15_20_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_15_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_15_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_15_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_15_20_1  (
            .in0(_gnd_net_),
            .in1(N__40579),
            .in2(N__46329),
            .in3(N__38422),
            .lcout(\current_shift_inst.un38_control_input_0_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_15_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_15_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_15_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_15_20_2  (
            .in0(_gnd_net_),
            .in1(N__40735),
            .in2(N__46326),
            .in3(N__38404),
            .lcout(\current_shift_inst.un38_control_input_0_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_15_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_15_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_15_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_15_20_3  (
            .in0(_gnd_net_),
            .in1(N__40723),
            .in2(N__46330),
            .in3(N__38401),
            .lcout(\current_shift_inst.un38_control_input_0_s1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_15_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_15_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_15_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_15_20_4  (
            .in0(_gnd_net_),
            .in1(N__40561),
            .in2(N__46327),
            .in3(N__38599),
            .lcout(\current_shift_inst.un38_control_input_0_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_15_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_15_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_15_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_15_20_5  (
            .in0(_gnd_net_),
            .in1(N__40621),
            .in2(N__46331),
            .in3(N__38596),
            .lcout(\current_shift_inst.un38_control_input_0_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_15_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_15_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_15_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_15_20_6  (
            .in0(_gnd_net_),
            .in1(N__40687),
            .in2(N__46328),
            .in3(N__38578),
            .lcout(\current_shift_inst.un38_control_input_0_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_15_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_15_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_15_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_15_20_7  (
            .in0(_gnd_net_),
            .in1(N__40753),
            .in2(N__46332),
            .in3(N__38560),
            .lcout(\current_shift_inst.un38_control_input_0_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_15_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_15_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_15_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_15_21_0  (
            .in0(_gnd_net_),
            .in1(N__41263),
            .in2(N__46366),
            .in3(N__38542),
            .lcout(\current_shift_inst.un38_control_input_0_s1_16 ),
            .ltout(),
            .carryin(bfn_15_21_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_15_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_15_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_15_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_15_21_1  (
            .in0(_gnd_net_),
            .in1(N__40699),
            .in2(N__46273),
            .in3(N__38524),
            .lcout(\current_shift_inst.un38_control_input_0_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_15_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_15_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_15_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_15_21_2  (
            .in0(_gnd_net_),
            .in1(N__40813),
            .in2(N__46367),
            .in3(N__38506),
            .lcout(\current_shift_inst.un38_control_input_0_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_15_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_15_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_15_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_15_21_3  (
            .in0(_gnd_net_),
            .in1(N__40693),
            .in2(N__46274),
            .in3(N__38488),
            .lcout(\current_shift_inst.un38_control_input_0_s1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_15_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_15_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_15_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_15_21_4  (
            .in0(_gnd_net_),
            .in1(N__40801),
            .in2(N__46368),
            .in3(N__38737),
            .lcout(\current_shift_inst.un38_control_input_0_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_15_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_15_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_15_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_15_21_5  (
            .in0(_gnd_net_),
            .in1(N__41275),
            .in2(N__46275),
            .in3(N__38719),
            .lcout(\current_shift_inst.un38_control_input_0_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_15_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_15_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_15_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_15_21_6  (
            .in0(_gnd_net_),
            .in1(N__40795),
            .in2(N__46369),
            .in3(N__38704),
            .lcout(\current_shift_inst.un38_control_input_0_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_15_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_15_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_15_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_15_21_7  (
            .in0(_gnd_net_),
            .in1(N__40807),
            .in2(N__46276),
            .in3(N__38686),
            .lcout(\current_shift_inst.un38_control_input_0_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_15_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_15_22_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_15_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_15_22_0  (
            .in0(_gnd_net_),
            .in1(N__40639),
            .in2(N__46375),
            .in3(N__38671),
            .lcout(\current_shift_inst.un38_control_input_0_s1_24 ),
            .ltout(),
            .carryin(bfn_15_22_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_15_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_15_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_15_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_15_22_1  (
            .in0(_gnd_net_),
            .in1(N__40759),
            .in2(N__46370),
            .in3(N__38659),
            .lcout(\current_shift_inst.un38_control_input_0_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_15_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_15_22_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_15_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_15_22_2  (
            .in0(_gnd_net_),
            .in1(N__40765),
            .in2(N__46376),
            .in3(N__38647),
            .lcout(\current_shift_inst.un38_control_input_0_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_15_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_15_22_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_15_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_15_22_3  (
            .in0(_gnd_net_),
            .in1(N__41269),
            .in2(N__46371),
            .in3(N__38632),
            .lcout(\current_shift_inst.un38_control_input_0_s1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_15_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_15_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_15_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_15_22_4  (
            .in0(_gnd_net_),
            .in1(N__46283),
            .in2(N__40747),
            .in3(N__38617),
            .lcout(\current_shift_inst.un38_control_input_0_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_15_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_15_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_15_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_15_22_5  (
            .in0(_gnd_net_),
            .in1(N__40789),
            .in2(N__46372),
            .in3(N__39085),
            .lcout(\current_shift_inst.un38_control_input_0_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIJ39T_LC_15_22_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIJ39T_LC_15_22_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIJ39T_LC_15_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s1_c_RNIJ39T_LC_15_22_6  (
            .in0(_gnd_net_),
            .in1(N__40776),
            .in2(N__46377),
            .in3(N__39070),
            .lcout(\current_shift_inst.un38_control_input_0_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_RNO_2_25_LC_15_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_RNO_2_25_LC_15_22_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_RNO_2_25_LC_15_22_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \current_shift_inst.control_input_RNO_2_25_LC_15_22_7  (
            .in0(N__46800),
            .in1(N__46315),
            .in2(_gnd_net_),
            .in3(N__39067),
            .lcout(\current_shift_inst.un38_control_input_0_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_15_25_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_15_25_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_15_25_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_15_25_0  (
            .in0(N__39048),
            .in1(N__39018),
            .in2(N__38991),
            .in3(N__38961),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_15_26_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_15_26_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_15_26_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_15_26_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38911),
            .lcout(\delay_measurement_inst.elapsed_time_hc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50140),
            .ce(N__38812),
            .sr(N__49717));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_15_26_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_15_26_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_15_26_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_15_26_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38863),
            .lcout(\delay_measurement_inst.elapsed_time_hc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50140),
            .ce(N__38812),
            .sr(N__49717));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_1_3_LC_15_27_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_1_3_LC_15_27_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_1_3_LC_15_27_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto30_1_3_LC_15_27_1  (
            .in0(_gnd_net_),
            .in1(N__41244),
            .in2(_gnd_net_),
            .in3(N__41256),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un1_startlto30_1Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_1_LC_15_27_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_1_LC_15_27_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_1_LC_15_27_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto30_1_LC_15_27_2  (
            .in0(N__40902),
            .in1(N__41232),
            .in2(N__38791),
            .in3(N__38788),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto30Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_16_2_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_16_2_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_16_2_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_16_2_2  (
            .in0(_gnd_net_),
            .in1(N__39134),
            .in2(_gnd_net_),
            .in3(N__39115),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_304_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.start_timer_tr_LC_16_3_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_tr_LC_16_3_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.start_timer_tr_LC_16_3_1 .LUT_INIT=16'b1100110001100110;
    LogicCell40 \delay_measurement_inst.start_timer_tr_LC_16_3_1  (
            .in0(N__39189),
            .in1(N__39207),
            .in2(_gnd_net_),
            .in3(N__39167),
            .lcout(\delay_measurement_inst.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50272),
            .ce(),
            .sr(N__49603));
    defparam \delay_measurement_inst.prev_tr_sig_LC_16_3_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.prev_tr_sig_LC_16_3_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.prev_tr_sig_LC_16_3_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.prev_tr_sig_LC_16_3_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39190),
            .lcout(\delay_measurement_inst.prev_tr_sigZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50272),
            .ce(),
            .sr(N__49603));
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_16_3_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_16_3_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_16_3_4 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_LC_16_3_4  (
            .in0(N__39151),
            .in1(N__39138),
            .in2(_gnd_net_),
            .in3(N__39118),
            .lcout(\delay_measurement_inst.delay_tr_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50272),
            .ce(),
            .sr(N__49603));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_4_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_4_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_4_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39116),
            .lcout(\delay_measurement_inst.delay_tr_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_16_4_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_16_4_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_16_4_5 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_16_4_5  (
            .in0(N__39150),
            .in1(N__39139),
            .in2(_gnd_net_),
            .in3(N__39117),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_305_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_16_5_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_16_5_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_16_5_1 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_0_LC_16_5_1  (
            .in0(N__45112),
            .in1(N__45340),
            .in2(_gnd_net_),
            .in3(N__39268),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50263),
            .ce(),
            .sr(N__49608));
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_16_6_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_16_6_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_16_6_1 .LUT_INIT=16'b0011000011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_4_LC_16_6_1  (
            .in0(N__45136),
            .in1(N__45303),
            .in2(N__44935),
            .in3(N__39613),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50257),
            .ce(),
            .sr(N__49609));
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_16_6_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_16_6_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_16_6_6 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_2_LC_16_6_6  (
            .in0(N__45301),
            .in1(N__45137),
            .in2(_gnd_net_),
            .in3(N__39658),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50257),
            .ce(),
            .sr(N__49609));
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_16_6_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_16_6_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_16_6_7 .LUT_INIT=16'b0011000011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_22_LC_16_6_7  (
            .in0(N__45135),
            .in1(N__45302),
            .in2(N__44934),
            .in3(N__39862),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50257),
            .ce(),
            .sr(N__49609));
    defparam \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_16_7_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_16_7_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_16_7_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_16_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39425),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_16_7_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_16_7_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_16_7_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_16_7_1  (
            .in0(N__40854),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_16_7_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_16_7_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_16_7_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_16_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39377),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_16_7_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_16_7_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_16_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_16_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39331),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_16_7_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_16_7_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_16_7_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_16_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41428),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_16_8_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_16_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_16_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_16_8_0  (
            .in0(_gnd_net_),
            .in1(N__39309),
            .in2(N__39310),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_8_0_),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_0_LC_16_8_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_0_LC_16_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_0_LC_16_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_0_LC_16_8_1  (
            .in0(_gnd_net_),
            .in1(N__39292),
            .in2(N__39285),
            .in3(N__39259),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_16_8_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_16_8_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_16_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_16_8_2  (
            .in0(_gnd_net_),
            .in1(N__39256),
            .in2(N__39250),
            .in3(N__39226),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_16_8_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_16_8_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_16_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_16_8_3  (
            .in0(_gnd_net_),
            .in1(N__39673),
            .in2(N__39667),
            .in3(N__39649),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_16_8_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_16_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_16_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_16_8_4  (
            .in0(_gnd_net_),
            .in1(N__39646),
            .in2(N__39640),
            .in3(N__39631),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_16_8_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_16_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_16_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_16_8_5  (
            .in0(_gnd_net_),
            .in1(N__39628),
            .in2(N__39622),
            .in3(N__39604),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_16_8_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_16_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_16_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_16_8_6  (
            .in0(_gnd_net_),
            .in1(N__39601),
            .in2(N__39595),
            .in3(N__39580),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_16_8_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_16_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_16_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_16_8_7  (
            .in0(_gnd_net_),
            .in1(N__39577),
            .in2(N__39571),
            .in3(N__39553),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_16_9_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_16_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_16_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_16_9_0  (
            .in0(_gnd_net_),
            .in1(N__39550),
            .in2(N__44152),
            .in3(N__39541),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(bfn_16_9_0_),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_16_9_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_16_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_16_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_16_9_1  (
            .in0(_gnd_net_),
            .in1(N__39538),
            .in2(N__41473),
            .in3(N__39532),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_7 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_16_9_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_16_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_16_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_16_9_2  (
            .in0(_gnd_net_),
            .in1(N__39529),
            .in2(N__39517),
            .in3(N__39496),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_16_9_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_16_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_16_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_16_9_3  (
            .in0(_gnd_net_),
            .in1(N__43825),
            .in2(N__44218),
            .in3(N__39814),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_16_9_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_16_9_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_16_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_16_9_4  (
            .in0(_gnd_net_),
            .in1(N__39811),
            .in2(N__39805),
            .in3(N__39796),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_16_9_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_16_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_16_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_16_9_5  (
            .in0(_gnd_net_),
            .in1(N__39793),
            .in2(N__41629),
            .in3(N__39787),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_16_9_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_16_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_16_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_16_9_6  (
            .in0(_gnd_net_),
            .in1(N__44227),
            .in2(N__44095),
            .in3(N__39772),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_16_9_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_16_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_16_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_16_9_7  (
            .in0(_gnd_net_),
            .in1(N__41530),
            .in2(N__41482),
            .in3(N__39757),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_16_10_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_16_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_16_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_16_10_0  (
            .in0(_gnd_net_),
            .in1(N__39754),
            .in2(N__39748),
            .in3(N__39724),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(bfn_16_10_0_),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_16_10_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_16_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_16_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_16_10_1  (
            .in0(_gnd_net_),
            .in1(N__39721),
            .in2(N__39715),
            .in3(N__39694),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_16_10_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_16_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_16_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_16_10_2  (
            .in0(_gnd_net_),
            .in1(N__41812),
            .in2(N__39691),
            .in3(N__39676),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_16_10_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_16_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_16_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_16_10_3  (
            .in0(_gnd_net_),
            .in1(N__39925),
            .in2(N__40351),
            .in3(N__39919),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_16_10_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_16_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_16_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_16_10_4  (
            .in0(_gnd_net_),
            .in1(N__40339),
            .in2(N__39916),
            .in3(N__39907),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_16_10_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_16_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_16_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_16_10_5  (
            .in0(_gnd_net_),
            .in1(N__40288),
            .in2(N__39952),
            .in3(N__39904),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_16_10_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_16_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_16_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_16_10_6  (
            .in0(_gnd_net_),
            .in1(N__41398),
            .in2(N__39901),
            .in3(N__39886),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_16_10_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_16_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_16_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_16_10_7  (
            .in0(_gnd_net_),
            .in1(N__39883),
            .in2(N__39877),
            .in3(N__39853),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_16_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_16_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_16_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_16_11_0  (
            .in0(_gnd_net_),
            .in1(N__39850),
            .in2(N__44407),
            .in3(N__39844),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ),
            .ltout(),
            .carryin(bfn_16_11_0_),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_16_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_16_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_16_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_16_11_1  (
            .in0(_gnd_net_),
            .in1(N__39841),
            .in2(N__44533),
            .in3(N__39826),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_16_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_16_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_16_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_16_11_2  (
            .in0(_gnd_net_),
            .in1(N__39823),
            .in2(N__40828),
            .in3(N__39817),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_16_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_16_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_16_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_16_11_3  (
            .in0(_gnd_net_),
            .in1(N__40087),
            .in2(N__44593),
            .in3(N__40081),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_16_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_16_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_16_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_16_11_4  (
            .in0(_gnd_net_),
            .in1(N__40078),
            .in2(N__40066),
            .in3(N__40045),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_16_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_16_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_16_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_16_11_5  (
            .in0(_gnd_net_),
            .in1(N__39935),
            .in2(N__44473),
            .in3(N__40042),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_16_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_16_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_16_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_16_11_6  (
            .in0(_gnd_net_),
            .in1(N__39958),
            .in2(N__39940),
            .in3(N__40030),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_16_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_16_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_16_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_16_11_7  (
            .in0(_gnd_net_),
            .in1(N__39939),
            .in2(N__40027),
            .in3(N__40003),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_16_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_16_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_16_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_16_12_0  (
            .in0(N__43998),
            .in1(N__44852),
            .in2(_gnd_net_),
            .in3(N__40000),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_16_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_16_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_16_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_16_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39997),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_16_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_16_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_16_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_16_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40240),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIGNK3_26_LC_16_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIGNK3_26_LC_16_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIGNK3_26_LC_16_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIGNK3_26_LC_16_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43997),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_i_0_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_16_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_16_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_16_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_16_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40182),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_16_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_16_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_16_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_16_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40117),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNICIEQ_24_LC_16_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNICIEQ_24_LC_16_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNICIEQ_24_LC_16_13_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNICIEQ_24_LC_16_13_0  (
            .in0(N__43996),
            .in1(N__40326),
            .in2(N__40258),
            .in3(N__40300),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNICIEQZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_16_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_16_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_16_13_2 .LUT_INIT=16'b0101000011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_20_LC_16_13_2  (
            .in0(N__45249),
            .in1(N__45132),
            .in2(N__44923),
            .in3(N__40279),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50213),
            .ce(),
            .sr(N__49631));
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_16_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_16_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_16_13_3 .LUT_INIT=16'b0011000011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_18_LC_16_13_3  (
            .in0(N__45130),
            .in1(N__45250),
            .in2(N__44911),
            .in3(N__40216),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50213),
            .ce(),
            .sr(N__49631));
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_16_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_16_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_16_13_5 .LUT_INIT=16'b0011000011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_19_LC_16_13_5  (
            .in0(N__45131),
            .in1(N__45251),
            .in2(N__44912),
            .in3(N__40159),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50213),
            .ce(),
            .sr(N__49631));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_16_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_16_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_16_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_16_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40372),
            .lcout(\current_shift_inst.un4_control_input_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_16_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_16_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_16_14_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_16_14_2  (
            .in0(N__46682),
            .in1(N__47478),
            .in2(N__46374),
            .in3(N__42576),
            .lcout(\current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_16_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_16_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_16_14_3 .LUT_INIT=16'b1000101110001011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_16_14_3  (
            .in0(N__42577),
            .in1(N__46681),
            .in2(N__47482),
            .in3(N__46301),
            .lcout(\current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_16_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_16_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_16_14_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_16_14_4  (
            .in0(N__47223),
            .in1(N__47477),
            .in2(_gnd_net_),
            .in3(N__42575),
            .lcout(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_16_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_16_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_16_14_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_16_14_5  (
            .in0(N__47226),
            .in1(N__47829),
            .in2(_gnd_net_),
            .in3(N__47399),
            .lcout(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_16_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_16_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_16_14_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_16_14_6  (
            .in0(N__47224),
            .in1(N__47901),
            .in2(_gnd_net_),
            .in3(N__42551),
            .lcout(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_14_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_14_7  (
            .in0(N__47225),
            .in1(N__47449),
            .in2(_gnd_net_),
            .in3(N__45563),
            .lcout(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_16_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_16_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_16_15_0 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_16_15_0  (
            .in0(N__46679),
            .in1(N__42591),
            .in2(N__40426),
            .in3(N__40374),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_16_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_16_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_16_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_16_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48778),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50203),
            .ce(N__48267),
            .sr(N__49646));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_16_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_16_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_16_15_3 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_16_15_3  (
            .in0(N__40375),
            .in1(N__46678),
            .in2(N__42595),
            .in3(N__40424),
            .lcout(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_16_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_16_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_16_15_4 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_16_15_4  (
            .in0(N__47265),
            .in1(N__42590),
            .in2(_gnd_net_),
            .in3(N__40373),
            .lcout(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_16_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_16_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_16_15_7 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_16_15_7  (
            .in0(N__43280),
            .in1(N__46680),
            .in2(_gnd_net_),
            .in3(N__48426),
            .lcout(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_16_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_16_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_16_16_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_16_16_0  (
            .in0(N__47586),
            .in1(N__47280),
            .in2(_gnd_net_),
            .in3(N__42869),
            .lcout(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_16_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_16_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_16_16_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_16_16_1  (
            .in0(N__47277),
            .in1(N__47795),
            .in2(_gnd_net_),
            .in3(N__42986),
            .lcout(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_16_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_16_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_16_16_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_16_16_2  (
            .in0(N__47630),
            .in1(N__47279),
            .in2(_gnd_net_),
            .in3(N__42899),
            .lcout(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_16_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_16_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_16_16_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_16_16_3  (
            .in0(N__47281),
            .in1(N__48188),
            .in2(_gnd_net_),
            .in3(N__42806),
            .lcout(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_16_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_16_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_16_16_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_16_16_4  (
            .in0(N__47267),
            .in1(N__47673),
            .in2(_gnd_net_),
            .in3(N__47111),
            .lcout(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_16_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_16_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_16_16_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_16_16_5  (
            .in0(N__48233),
            .in1(N__47268),
            .in2(_gnd_net_),
            .in3(N__42839),
            .lcout(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_16_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_16_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_16_16_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_16_16_6  (
            .in0(N__47266),
            .in1(N__47709),
            .in2(_gnd_net_),
            .in3(N__42929),
            .lcout(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_16_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_16_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_16_16_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_16_16_7  (
            .in0(N__47278),
            .in1(N__47750),
            .in2(_gnd_net_),
            .in3(N__42959),
            .lcout(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_16_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_16_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_16_17_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_16_17_0  (
            .in0(N__47273),
            .in1(N__48018),
            .in2(_gnd_net_),
            .in3(N__43127),
            .lcout(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_16_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_16_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_16_17_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_16_17_1  (
            .in0(N__47269),
            .in1(N__48144),
            .in2(_gnd_net_),
            .in3(N__45503),
            .lcout(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_16_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_16_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_16_17_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_16_17_2  (
            .in0(N__47272),
            .in1(N__48099),
            .in2(_gnd_net_),
            .in3(N__43364),
            .lcout(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_16_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_16_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_16_17_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_16_17_3  (
            .in0(N__47270),
            .in1(N__48578),
            .in2(_gnd_net_),
            .in3(N__43041),
            .lcout(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_16_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_16_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_16_17_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_16_17_4  (
            .in0(N__46704),
            .in1(N__48019),
            .in2(N__46324),
            .in3(N__43128),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_16_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_16_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_16_17_5 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_16_17_5  (
            .in0(N__46702),
            .in1(N__42960),
            .in2(N__46229),
            .in3(N__47751),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_16_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_16_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_16_17_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_16_17_6  (
            .in0(N__48537),
            .in1(N__47271),
            .in2(_gnd_net_),
            .in3(N__43163),
            .lcout(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_16_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_16_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_16_17_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_16_17_7  (
            .in0(N__46703),
            .in1(N__47631),
            .in2(N__46230),
            .in3(N__42900),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_18_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_18_0  (
            .in0(N__47275),
            .in1(N__48498),
            .in2(_gnd_net_),
            .in3(N__43016),
            .lcout(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_16_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_16_18_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_16_18_1  (
            .in0(N__46690),
            .in1(N__48381),
            .in2(_gnd_net_),
            .in3(N__43313),
            .lcout(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_16_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_16_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_16_18_2 .LUT_INIT=16'b1000101110001011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_16_18_2  (
            .in0(N__43107),
            .in1(N__46691),
            .in2(N__47986),
            .in3(N__46152),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_16_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_16_18_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_16_18_3  (
            .in0(N__46689),
            .in1(N__48465),
            .in2(_gnd_net_),
            .in3(N__43694),
            .lcout(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_16_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_16_18_4 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_16_18_4  (
            .in0(N__42559),
            .in1(N__46688),
            .in2(N__46290),
            .in3(N__47900),
            .lcout(\current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_16_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_16_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_16_18_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_16_18_5  (
            .in0(N__47276),
            .in1(N__47981),
            .in2(_gnd_net_),
            .in3(N__43106),
            .lcout(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_16_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_16_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_16_18_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_16_18_6  (
            .in0(N__47274),
            .in1(N__47952),
            .in2(_gnd_net_),
            .in3(N__43076),
            .lcout(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_16_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_16_18_7 .LUT_INIT=16'b1000101110001011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_16_18_7  (
            .in0(N__43017),
            .in1(N__46799),
            .in2(N__48502),
            .in3(N__46098),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_16_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_16_19_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_16_19_0  (
            .in0(N__46692),
            .in1(N__47796),
            .in2(N__46293),
            .in3(N__43000),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_16_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_16_19_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_16_19_1  (
            .in0(N__46687),
            .in1(N__47585),
            .in2(N__46320),
            .in3(N__42876),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_16_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_16_19_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_16_19_2  (
            .in0(N__48341),
            .in1(N__46684),
            .in2(_gnd_net_),
            .in3(N__43241),
            .lcout(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_16_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_16_19_3 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_16_19_3  (
            .in0(N__43242),
            .in1(N__46694),
            .in2(N__46319),
            .in3(N__48342),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_16_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_16_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_16_19_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_16_19_4  (
            .in0(N__46693),
            .in1(N__47708),
            .in2(N__46291),
            .in3(N__42940),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_16_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_16_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_16_19_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_16_19_5  (
            .in0(N__46685),
            .in1(N__48302),
            .in2(_gnd_net_),
            .in3(N__43217),
            .lcout(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_16_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_16_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_16_19_6 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_16_19_6  (
            .in0(N__47116),
            .in1(N__46686),
            .in2(N__46292),
            .in3(N__47672),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNID8O11_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_16_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_16_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_16_19_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_16_19_7  (
            .in0(N__46683),
            .in1(N__47447),
            .in2(N__46321),
            .in3(N__45574),
            .lcout(\current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_16_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_16_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_16_20_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_16_20_0  (
            .in0(N__46813),
            .in1(N__48307),
            .in2(N__46296),
            .in3(N__43224),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_16_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_16_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_16_20_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_16_20_2  (
            .in0(N__46810),
            .in1(N__48100),
            .in2(N__46297),
            .in3(N__43375),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_16_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_16_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_16_20_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_16_20_3  (
            .in0(N__46701),
            .in1(N__48017),
            .in2(N__46334),
            .in3(N__43132),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJO221_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_16_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_16_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_16_20_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_16_20_4  (
            .in0(N__46809),
            .in1(N__48234),
            .in2(N__46294),
            .in3(N__42850),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_16_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_16_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_16_20_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_16_20_5  (
            .in0(N__46700),
            .in1(N__48056),
            .in2(N__46333),
            .in3(N__45441),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI25021_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_16_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_16_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_16_20_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_16_20_6  (
            .in0(N__46812),
            .in1(N__48538),
            .in2(N__46295),
            .in3(N__43171),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_16_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_16_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_16_20_7 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_16_20_7  (
            .in0(N__47985),
            .in1(N__46811),
            .in2(N__46335),
            .in3(N__43111),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_16_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_16_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_16_21_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_16_21_0  (
            .in0(N__46697),
            .in1(N__48579),
            .in2(N__46302),
            .in3(N__43053),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_16_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_16_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_16_21_2 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_16_21_2  (
            .in0(N__43225),
            .in1(N__46817),
            .in2(N__46303),
            .in3(N__48303),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIF4PE_LC_16_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIF4PE_LC_16_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIF4PE_LC_16_21_3 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIF4PE_LC_16_21_3  (
            .in0(_gnd_net_),
            .in1(N__46699),
            .in2(_gnd_net_),
            .in3(N__43198),
            .lcout(\current_shift_inst.un4_control_input_0_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_16_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_16_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_16_21_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_16_21_4  (
            .in0(N__46698),
            .in1(N__48419),
            .in2(N__46305),
            .in3(N__43287),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_16_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_16_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_16_21_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_16_21_5  (
            .in0(N__46816),
            .in1(N__48466),
            .in2(N__46323),
            .in3(N__43705),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_16_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_16_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_16_21_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_16_21_6  (
            .in0(N__46695),
            .in1(N__48189),
            .in2(N__46304),
            .in3(N__42820),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_16_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_16_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_16_21_7 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_16_21_7  (
            .in0(N__47948),
            .in1(N__46696),
            .in2(N__46322),
            .in3(N__43090),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_16_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_16_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_16_22_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_16_22_5  (
            .in0(N__46815),
            .in1(N__48382),
            .in2(N__46378),
            .in3(N__43324),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_16_22_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_16_22_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_16_22_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_16_22_6  (
            .in0(N__46814),
            .in1(N__48145),
            .in2(N__46373),
            .in3(N__45517),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISST11_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_29_LC_16_26_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_29_LC_16_26_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_29_LC_16_26_5 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_29_LC_16_26_5  (
            .in0(N__41187),
            .in1(N__41257),
            .in2(_gnd_net_),
            .in3(N__41050),
            .lcout(measured_delay_hc_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50146),
            .ce(),
            .sr(N__49710));
    defparam \delay_measurement_inst.delay_hc_reg_30_LC_16_27_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_30_LC_16_27_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_30_LC_16_27_0 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_30_LC_16_27_0  (
            .in0(N__41042),
            .in1(_gnd_net_),
            .in2(N__41221),
            .in3(N__41245),
            .lcout(measured_delay_hc_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50141),
            .ce(),
            .sr(N__49718));
    defparam \delay_measurement_inst.delay_hc_reg_27_LC_16_27_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_27_LC_16_27_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_27_LC_16_27_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_27_LC_16_27_1  (
            .in0(N__41233),
            .in1(N__41214),
            .in2(_gnd_net_),
            .in3(N__41040),
            .lcout(measured_delay_hc_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50141),
            .ce(),
            .sr(N__49718));
    defparam \delay_measurement_inst.delay_hc_reg_28_LC_16_27_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_28_LC_16_27_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_28_LC_16_27_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_28_LC_16_27_3  (
            .in0(N__40903),
            .in1(N__41215),
            .in2(_gnd_net_),
            .in3(N__41041),
            .lcout(measured_delay_hc_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50141),
            .ce(),
            .sr(N__49718));
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_17_5_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_17_5_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_17_5_6 .LUT_INIT=16'b0001000111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_3_LC_17_5_6  (
            .in0(N__45138),
            .in1(N__45339),
            .in2(_gnd_net_),
            .in3(N__40891),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50268),
            .ce(),
            .sr(N__49607));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_17_6_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_17_6_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_17_6_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_17_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41319),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_17_7_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_17_7_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_17_7_7 .LUT_INIT=16'b0011000011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_21_LC_17_7_7  (
            .in0(N__45134),
            .in1(N__45281),
            .in2(N__44883),
            .in3(N__41584),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50258),
            .ce(),
            .sr(N__49610));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIOTCP_18_LC_17_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIOTCP_18_LC_17_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIOTCP_18_LC_17_8_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIOTCP_18_LC_17_8_0  (
            .in0(N__44083),
            .in1(N__41571),
            .in2(N__41524),
            .in3(N__41542),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIOTCPZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_17_8_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_17_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_17_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_17_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41519),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_17_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_17_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_17_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_17_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43612),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_17_8_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_17_8_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_17_8_7 .LUT_INIT=16'b0000000111110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_8_LC_17_8_7  (
            .in0(N__45133),
            .in1(N__44768),
            .in2(N__45321),
            .in3(N__41464),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50253),
            .ce(),
            .sr(N__49613));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIGNFQ_25_LC_17_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIGNFQ_25_LC_17_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIGNFQ_25_LC_17_9_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIGNFQ_25_LC_17_9_0  (
            .in0(N__44082),
            .in1(N__41391),
            .in2(N__41453),
            .in3(N__41410),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIGNFQZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIFMK3_25_LC_17_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIFMK3_25_LC_17_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIFMK3_25_LC_17_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIFMK3_25_LC_17_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41390),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_17_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_17_9_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_17_9_5 .LUT_INIT=16'b0011000011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_25_LC_17_9_5  (
            .in0(N__45046),
            .in1(N__45322),
            .in2(N__44810),
            .in3(N__41353),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50247),
            .ce(),
            .sr(N__49614));
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_17_9_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_17_9_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_17_9_7 .LUT_INIT=16'b0011000011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_26_LC_17_9_7  (
            .in0(N__45047),
            .in1(N__45323),
            .in2(N__44811),
            .in3(N__41284),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50247),
            .ce(),
            .sr(N__49614));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI9BAQ_21_LC_17_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI9BAQ_21_LC_17_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI9BAQ_21_LC_17_10_0 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI9BAQ_21_LC_17_10_0  (
            .in0(N__41854),
            .in1(N__44077),
            .in2(N__41778),
            .in3(N__41841),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNI9BAQZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_17_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_17_10_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_17_10_2 .LUT_INIT=16'b0011000011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_17_LC_17_10_2  (
            .in0(N__45126),
            .in1(N__45305),
            .in2(N__44866),
            .in3(N__41806),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50241),
            .ce(),
            .sr(N__49617));
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_17_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_17_10_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_17_10_4 .LUT_INIT=16'b0011000011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_11_LC_17_10_4  (
            .in0(N__45125),
            .in1(N__45304),
            .in2(N__44865),
            .in3(N__41746),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50241),
            .ce(),
            .sr(N__49617));
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_17_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_17_10_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_17_10_6 .LUT_INIT=16'b0101010111011100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_12_LC_17_10_6  (
            .in0(N__41680),
            .in1(N__44799),
            .in2(N__45139),
            .in3(N__45306),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50241),
            .ce(),
            .sr(N__49617));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_17_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_17_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_17_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_17_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41640),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_11_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_11_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_11_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_11_0  (
            .in0(N__42780),
            .in1(N__50321),
            .in2(_gnd_net_),
            .in3(N__41617),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_17_11_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .clk(N__50235),
            .ce(N__42623),
            .sr(N__49618));
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_11_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_11_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_11_1  (
            .in0(N__42776),
            .in1(N__44327),
            .in2(_gnd_net_),
            .in3(N__41614),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .clk(N__50235),
            .ce(N__42623),
            .sr(N__49618));
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_11_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_11_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_11_2  (
            .in0(N__42781),
            .in1(N__41603),
            .in2(_gnd_net_),
            .in3(N__41587),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .clk(N__50235),
            .ce(N__42623),
            .sr(N__49618));
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_11_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_11_3  (
            .in0(N__42777),
            .in1(N__42083),
            .in2(_gnd_net_),
            .in3(N__42067),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .clk(N__50235),
            .ce(N__42623),
            .sr(N__49618));
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_11_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_11_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_11_4  (
            .in0(N__42782),
            .in1(N__42062),
            .in2(_gnd_net_),
            .in3(N__42046),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .clk(N__50235),
            .ce(N__42623),
            .sr(N__49618));
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_11_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_11_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_11_5  (
            .in0(N__42778),
            .in1(N__42036),
            .in2(_gnd_net_),
            .in3(N__42022),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .clk(N__50235),
            .ce(N__42623),
            .sr(N__49618));
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_11_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_11_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_11_6  (
            .in0(N__42783),
            .in1(N__42011),
            .in2(_gnd_net_),
            .in3(N__41995),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .clk(N__50235),
            .ce(N__42623),
            .sr(N__49618));
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_11_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_11_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_11_7  (
            .in0(N__42779),
            .in1(N__41984),
            .in2(_gnd_net_),
            .in3(N__41968),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .clk(N__50235),
            .ce(N__42623),
            .sr(N__49618));
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_12_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_12_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_12_0  (
            .in0(N__42775),
            .in1(N__41960),
            .in2(_gnd_net_),
            .in3(N__41941),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_17_12_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .clk(N__50230),
            .ce(N__42639),
            .sr(N__49622));
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_12_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_12_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_12_1  (
            .in0(N__42771),
            .in1(N__41927),
            .in2(_gnd_net_),
            .in3(N__41911),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .clk(N__50230),
            .ce(N__42639),
            .sr(N__49622));
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_12_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_12_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_12_2  (
            .in0(N__42772),
            .in1(N__41900),
            .in2(_gnd_net_),
            .in3(N__41884),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .clk(N__50230),
            .ce(N__42639),
            .sr(N__49622));
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_12_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_12_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_12_3  (
            .in0(N__42768),
            .in1(N__41873),
            .in2(_gnd_net_),
            .in3(N__41857),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .clk(N__50230),
            .ce(N__42639),
            .sr(N__49622));
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_12_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_12_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_12_4  (
            .in0(N__42773),
            .in1(N__42294),
            .in2(_gnd_net_),
            .in3(N__42280),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .clk(N__50230),
            .ce(N__42639),
            .sr(N__49622));
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_12_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_12_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_12_5  (
            .in0(N__42769),
            .in1(N__42275),
            .in2(_gnd_net_),
            .in3(N__42259),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .clk(N__50230),
            .ce(N__42639),
            .sr(N__49622));
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_12_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_12_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_12_6  (
            .in0(N__42774),
            .in1(N__42248),
            .in2(_gnd_net_),
            .in3(N__42232),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .clk(N__50230),
            .ce(N__42639),
            .sr(N__49622));
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_12_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_12_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_12_7  (
            .in0(N__42770),
            .in1(N__42221),
            .in2(_gnd_net_),
            .in3(N__42205),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .clk(N__50230),
            .ce(N__42639),
            .sr(N__49622));
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_13_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_13_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_13_0  (
            .in0(N__42764),
            .in1(N__42191),
            .in2(_gnd_net_),
            .in3(N__42175),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_17_13_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .clk(N__50223),
            .ce(N__42638),
            .sr(N__49626));
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_13_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_13_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_13_1  (
            .in0(N__42784),
            .in1(N__42167),
            .in2(_gnd_net_),
            .in3(N__42148),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .clk(N__50223),
            .ce(N__42638),
            .sr(N__49626));
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_13_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_13_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_13_2  (
            .in0(N__42765),
            .in1(N__42137),
            .in2(_gnd_net_),
            .in3(N__42121),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .clk(N__50223),
            .ce(N__42638),
            .sr(N__49626));
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_13_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_13_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_13_3  (
            .in0(N__42785),
            .in1(N__42110),
            .in2(_gnd_net_),
            .in3(N__42094),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .clk(N__50223),
            .ce(N__42638),
            .sr(N__49626));
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_13_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_13_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_13_4  (
            .in0(N__42766),
            .in1(N__42524),
            .in2(_gnd_net_),
            .in3(N__42508),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .clk(N__50223),
            .ce(N__42638),
            .sr(N__49626));
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_13_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_13_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_13_5  (
            .in0(N__42786),
            .in1(N__42503),
            .in2(_gnd_net_),
            .in3(N__42487),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .clk(N__50223),
            .ce(N__42638),
            .sr(N__49626));
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_13_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_13_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_13_6  (
            .in0(N__42767),
            .in1(N__42476),
            .in2(_gnd_net_),
            .in3(N__42460),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .clk(N__50223),
            .ce(N__42638),
            .sr(N__49626));
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_13_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_13_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_13_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_13_7  (
            .in0(N__42787),
            .in1(N__42449),
            .in2(_gnd_net_),
            .in3(N__42433),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .clk(N__50223),
            .ce(N__42638),
            .sr(N__49626));
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_14_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_14_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_14_0  (
            .in0(N__42758),
            .in1(N__42425),
            .in2(_gnd_net_),
            .in3(N__42406),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_17_14_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .clk(N__50214),
            .ce(N__42640),
            .sr(N__49632));
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_14_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_14_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_14_1  (
            .in0(N__42762),
            .in1(N__42392),
            .in2(_gnd_net_),
            .in3(N__42376),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .clk(N__50214),
            .ce(N__42640),
            .sr(N__49632));
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_14_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_14_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_14_2  (
            .in0(N__42759),
            .in1(N__42365),
            .in2(_gnd_net_),
            .in3(N__42349),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .clk(N__50214),
            .ce(N__42640),
            .sr(N__49632));
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_14_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_14_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_14_3  (
            .in0(N__42763),
            .in1(N__42338),
            .in2(_gnd_net_),
            .in3(N__42322),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .clk(N__50214),
            .ce(N__42640),
            .sr(N__49632));
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_14_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_14_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_14_4  (
            .in0(N__42760),
            .in1(N__42318),
            .in2(_gnd_net_),
            .in3(N__42304),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ),
            .clk(N__50214),
            .ce(N__42640),
            .sr(N__49632));
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_14_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_14_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_14_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_14_5  (
            .in0(N__42654),
            .in1(N__42761),
            .in2(_gnd_net_),
            .in3(N__42658),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50214),
            .ce(N__42640),
            .sr(N__49632));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_17_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_17_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_17_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_17_15_0  (
            .in0(_gnd_net_),
            .in1(N__42601),
            .in2(N__45390),
            .in3(N__45386),
            .lcout(\current_shift_inst.un4_control_input1_2 ),
            .ltout(),
            .carryin(bfn_17_15_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_17_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_17_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_17_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_17_15_1  (
            .in0(_gnd_net_),
            .in1(N__47356),
            .in2(_gnd_net_),
            .in3(N__42580),
            .lcout(\current_shift_inst.un4_control_input1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_1 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_17_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_17_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_17_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_17_15_2  (
            .in0(_gnd_net_),
            .in1(N__46825),
            .in2(_gnd_net_),
            .in3(N__42565),
            .lcout(\current_shift_inst.un4_control_input1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_2 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_17_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_17_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_17_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_17_15_3  (
            .in0(_gnd_net_),
            .in1(N__47344),
            .in2(_gnd_net_),
            .in3(N__42562),
            .lcout(\current_shift_inst.un4_control_input1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_3 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_17_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_17_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_17_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_17_15_4  (
            .in0(_gnd_net_),
            .in1(N__47338),
            .in2(_gnd_net_),
            .in3(N__42535),
            .lcout(\current_shift_inst.un4_control_input1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_4 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_17_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_17_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_17_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_17_15_5  (
            .in0(_gnd_net_),
            .in1(N__47350),
            .in2(_gnd_net_),
            .in3(N__42532),
            .lcout(\current_shift_inst.un4_control_input1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_5 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_17_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_17_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_17_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_17_15_6  (
            .in0(_gnd_net_),
            .in1(N__47362),
            .in2(_gnd_net_),
            .in3(N__42529),
            .lcout(\current_shift_inst.un4_control_input1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_6 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_17_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_17_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_17_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_17_15_7  (
            .in0(_gnd_net_),
            .in1(N__47287),
            .in2(_gnd_net_),
            .in3(N__42973),
            .lcout(\current_shift_inst.un4_control_input1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_7 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_17_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_17_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_17_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_17_16_0  (
            .in0(_gnd_net_),
            .in1(N__47320),
            .in2(_gnd_net_),
            .in3(N__42943),
            .lcout(\current_shift_inst.un4_control_input1_10 ),
            .ltout(),
            .carryin(bfn_17_16_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_17_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_17_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_17_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_17_16_1  (
            .in0(_gnd_net_),
            .in1(N__47533),
            .in2(_gnd_net_),
            .in3(N__42913),
            .lcout(\current_shift_inst.un4_control_input1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_9 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_17_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_17_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_17_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_17_16_2  (
            .in0(_gnd_net_),
            .in1(N__47332),
            .in2(_gnd_net_),
            .in3(N__42910),
            .lcout(\current_shift_inst.un4_control_input1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_10 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_17_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_17_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_17_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_17_16_3  (
            .in0(_gnd_net_),
            .in1(N__47527),
            .in2(_gnd_net_),
            .in3(N__42883),
            .lcout(\current_shift_inst.un4_control_input1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_11 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_17_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_17_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_17_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_17_16_4  (
            .in0(_gnd_net_),
            .in1(N__47326),
            .in2(_gnd_net_),
            .in3(N__42853),
            .lcout(\current_shift_inst.un4_control_input1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_12 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_17_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_17_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_17_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_17_16_5  (
            .in0(_gnd_net_),
            .in1(N__47551),
            .in2(_gnd_net_),
            .in3(N__42823),
            .lcout(\current_shift_inst.un4_control_input1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_13 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_17_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_17_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_17_16_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_17_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__47371),
            .in3(N__42793),
            .lcout(\current_shift_inst.un4_control_input1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_14 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_17_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_17_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_17_16_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_17_16_7  (
            .in0(_gnd_net_),
            .in1(N__47545),
            .in2(_gnd_net_),
            .in3(N__42790),
            .lcout(\current_shift_inst.un4_control_input1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_15 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_17_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_17_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_17_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_17_17_0  (
            .in0(_gnd_net_),
            .in1(N__43399),
            .in2(_gnd_net_),
            .in3(N__43138),
            .lcout(\current_shift_inst.un4_control_input1_18 ),
            .ltout(),
            .carryin(bfn_17_17_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_17_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_17_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_17_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_17_17_1  (
            .in0(_gnd_net_),
            .in1(N__43177),
            .in2(_gnd_net_),
            .in3(N__43135),
            .lcout(\current_shift_inst.un4_control_input1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_17 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_17_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_17_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_17_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_17_17_2  (
            .in0(_gnd_net_),
            .in1(N__43342),
            .in2(_gnd_net_),
            .in3(N__43114),
            .lcout(\current_shift_inst.un4_control_input1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_18 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_17_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_17_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_17_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_17_17_3  (
            .in0(_gnd_net_),
            .in1(N__43384),
            .in2(_gnd_net_),
            .in3(N__43093),
            .lcout(\current_shift_inst.un4_control_input1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_19 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_17_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_17_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_17_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_17_17_4  (
            .in0(_gnd_net_),
            .in1(N__43417),
            .in2(_gnd_net_),
            .in3(N__43063),
            .lcout(\current_shift_inst.un4_control_input1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_20 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_17_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_17_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_17_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_17_17_5  (
            .in0(_gnd_net_),
            .in1(N__43408),
            .in2(_gnd_net_),
            .in3(N__43030),
            .lcout(\current_shift_inst.un4_control_input1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_21 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_17_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_17_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_17_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_17_17_6  (
            .in0(_gnd_net_),
            .in1(N__47539),
            .in2(_gnd_net_),
            .in3(N__43027),
            .lcout(\current_shift_inst.un4_control_input1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_22 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_17_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_17_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_17_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_17_17_7  (
            .in0(_gnd_net_),
            .in1(N__43333),
            .in2(_gnd_net_),
            .in3(N__43003),
            .lcout(\current_shift_inst.un4_control_input1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_23 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_17_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_17_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_17_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_17_18_0  (
            .in0(_gnd_net_),
            .in1(N__43390),
            .in2(_gnd_net_),
            .in3(N__43291),
            .lcout(\current_shift_inst.un4_control_input1_26 ),
            .ltout(),
            .carryin(bfn_17_18_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_17_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_17_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_17_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_17_18_1  (
            .in0(_gnd_net_),
            .in1(N__43726),
            .in2(_gnd_net_),
            .in3(N__43258),
            .lcout(\current_shift_inst.un4_control_input1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_25 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_17_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_17_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_17_18_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_17_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__44281),
            .in3(N__43255),
            .lcout(\current_shift_inst.un4_control_input1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_26 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_17_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_17_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_17_18_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_17_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43717),
            .in3(N__43228),
            .lcout(\current_shift_inst.un4_control_input1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_27 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_17_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_17_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_17_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_17_18_4  (
            .in0(_gnd_net_),
            .in1(N__43672),
            .in2(_gnd_net_),
            .in3(N__43204),
            .lcout(\current_shift_inst.un4_control_input1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_28 ),
            .carryout(\current_shift_inst.un4_control_input1_31 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_17_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_17_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_17_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_17_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43201),
            .lcout(\current_shift_inst.un4_control_input1_31_THRU_CO ),
            .ltout(\current_shift_inst.un4_control_input1_31_THRU_CO_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_17_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_17_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_17_18_6 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_17_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43189),
            .in3(N__46801),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_17_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_17_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_17_18_7 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_17_18_7  (
            .in0(_gnd_net_),
            .in1(N__48049),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_17_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_17_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_17_19_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_17_19_0  (
            .in0(N__46803),
            .in1(N__48529),
            .in2(N__46418),
            .in3(N__43170),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_17_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_17_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_17_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_17_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47926),
            .lcout(\current_shift_inst.un4_control_input_1_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_17_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_17_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_17_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_17_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48559),
            .lcout(\current_shift_inst.un4_control_input_1_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_17_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_17_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_17_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_17_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48085),
            .lcout(\current_shift_inst.un4_control_input_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_17_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_17_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_17_19_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_17_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48451),
            .lcout(\current_shift_inst.un4_control_input_1_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_17_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_17_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_17_19_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_17_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47967),
            .lcout(\current_shift_inst.un4_control_input_1_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_17_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_17_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_17_19_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_17_19_6  (
            .in0(N__48086),
            .in1(N__46802),
            .in2(N__46419),
            .in3(N__43371),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_17_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_17_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_17_19_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_17_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48005),
            .lcout(\current_shift_inst.un4_control_input_1_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_17_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_17_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_17_20_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_17_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48485),
            .lcout(\current_shift_inst.un4_control_input_1_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_17_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_17_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_17_20_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_17_20_4  (
            .in0(N__48373),
            .in1(N__46819),
            .in2(N__46420),
            .in3(N__43320),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_17_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_17_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_17_20_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_17_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48403),
            .lcout(\current_shift_inst.un4_control_input_1_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_17_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_17_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_17_20_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_17_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48326),
            .lcout(\current_shift_inst.un4_control_input_1_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_17_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_17_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_17_20_7 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_17_20_7  (
            .in0(N__46818),
            .in1(N__43701),
            .in2(N__46379),
            .in3(N__48455),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_21_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48284),
            .lcout(\current_shift_inst.un4_control_input_1_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_17_28_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_17_28_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_17_28_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIUKI8_LC_17_28_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43663),
            .lcout(\current_shift_inst.timer_s1.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_18_7_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_18_7_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_18_7_4 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_18_7_4  (
            .in0(_gnd_net_),
            .in1(N__44178),
            .in2(_gnd_net_),
            .in3(N__43452),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_18_7_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_18_7_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_18_7_5 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_18_7_5  (
            .in0(N__43616),
            .in1(N__43590),
            .in2(N__43540),
            .in3(N__43537),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_18_8_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_18_8_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_18_8_2 .LUT_INIT=16'b0000000111001111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_5_LC_18_8_2  (
            .in0(N__45122),
            .in1(N__45297),
            .in2(N__44832),
            .in3(N__43486),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50259),
            .ce(),
            .sr(N__49611));
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_18_8_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_18_8_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_18_8_3 .LUT_INIT=16'b0000000110101111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_7_LC_18_8_3  (
            .in0(N__45296),
            .in1(N__45123),
            .in2(N__44833),
            .in3(N__43429),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50259),
            .ce(),
            .sr(N__49611));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIKOBP_17_LC_18_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIKOBP_17_LC_18_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIKOBP_17_LC_18_9_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIKOBP_17_LC_18_9_0  (
            .in0(N__44265),
            .in1(N__44081),
            .in2(N__44140),
            .in3(N__44236),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIKOBPZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_18_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_18_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_18_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_18_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43785),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_18_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_18_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_18_9_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_18_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44179),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_18_9_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_18_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_18_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_18_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44135),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI898P_14_LC_18_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI898P_14_LC_18_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI898P_14_LC_18_10_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI898P_14_LC_18_10_0  (
            .in0(N__44080),
            .in1(N__43872),
            .in2(N__43793),
            .in3(N__43837),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNI898PZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_18_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_18_10_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_18_10_2 .LUT_INIT=16'b0011000011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_10_LC_18_10_2  (
            .in0(N__45118),
            .in1(N__45309),
            .in2(N__44806),
            .in3(N__43813),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50248),
            .ce(),
            .sr(N__49615));
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_18_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_18_10_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_18_10_3 .LUT_INIT=16'b0101000011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_28_LC_18_10_3  (
            .in0(N__45307),
            .in1(N__45120),
            .in2(N__44808),
            .in3(N__43750),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50248),
            .ce(),
            .sr(N__49615));
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_18_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_18_10_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_18_10_6 .LUT_INIT=16'b0011000011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_23_LC_18_10_6  (
            .in0(N__45119),
            .in1(N__45310),
            .in2(N__44807),
            .in3(N__43738),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50248),
            .ce(),
            .sr(N__49615));
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_18_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_18_10_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_18_10_7 .LUT_INIT=16'b0101000011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_31_LC_18_10_7  (
            .in0(N__45308),
            .in1(N__45121),
            .in2(N__44809),
            .in3(N__44947),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50248),
            .ce(),
            .sr(N__49615));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_18_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_18_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_18_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_18_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44625),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_18_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_18_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_18_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_18_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44577),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_18_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_18_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_18_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_18_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44489),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_18_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_18_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_18_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_18_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44431),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2P9P1_20_LC_18_12_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2P9P1_20_LC_18_12_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2P9P1_20_LC_18_12_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2P9P1_20_LC_18_12_0  (
            .in0(N__44395),
            .in1(N__44383),
            .in2(N__44371),
            .in3(N__44356),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_18_12_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_18_12_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_18_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_18_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44331),
            .lcout(\delay_measurement_inst.elapsed_time_tr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50236),
            .ce(N__49815),
            .sr(N__49619));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_18_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_18_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_18_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_18_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48374),
            .lcout(\current_shift_inst.un4_control_input_1_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_18_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_18_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_18_13_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_18_13_2  (
            .in0(N__46756),
            .in1(N__47448),
            .in2(N__46423),
            .in3(N__45570),
            .lcout(\current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_18_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_18_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_18_13_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_18_13_3  (
            .in0(N__47863),
            .in1(N__46757),
            .in2(N__46421),
            .in3(N__47080),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_18_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_18_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_18_13_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_18_13_4  (
            .in0(N__46758),
            .in1(N__48143),
            .in2(N__46422),
            .in3(N__45516),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISST11_0_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_18_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_18_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_18_13_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_18_13_5  (
            .in0(N__47862),
            .in1(N__47215),
            .in2(_gnd_net_),
            .in3(N__47079),
            .lcout(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_RNO_1_25_LC_18_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_RNO_1_25_LC_18_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_RNO_1_25_LC_18_14_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.control_input_RNO_1_25_LC_18_14_2  (
            .in0(_gnd_net_),
            .in1(N__46798),
            .in2(_gnd_net_),
            .in3(N__46339),
            .lcout(\current_shift_inst.un38_control_input_axb_31_s0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_18_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_18_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_18_14_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_18_14_3  (
            .in0(N__47219),
            .in1(N__48057),
            .in2(_gnd_net_),
            .in3(N__45440),
            .lcout(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_18_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_18_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_18_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_18_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47300),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_1 ),
            .ltout(\current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_18_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_18_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_18_14_5 .LUT_INIT=16'b0000111101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_18_14_5  (
            .in0(N__47301),
            .in1(_gnd_net_),
            .in2(N__45367),
            .in3(N__47188),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_18_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_18_14_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_18_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_18_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48845),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50224),
            .ce(N__48268),
            .sr(N__49627));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_18_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_18_14_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_18_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_18_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48814),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50224),
            .ce(N__48268),
            .sr(N__49627));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_18_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_18_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_18_15_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_18_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47785),
            .lcout(\current_shift_inst.un4_control_input_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_18_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_18_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_18_15_2 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_18_15_2  (
            .in0(N__47192),
            .in1(N__47136),
            .in2(_gnd_net_),
            .in3(N__47508),
            .lcout(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_18_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_18_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_18_15_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_18_15_3  (
            .in0(N__46706),
            .in1(N__47674),
            .in2(N__46408),
            .in3(N__47112),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_18_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_18_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_18_15_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_18_15_5  (
            .in0(N__46705),
            .in1(N__47861),
            .in2(N__46407),
            .in3(N__47078),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_18_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_18_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_18_15_6 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_18_15_6  (
            .in0(N__47050),
            .in1(N__47035),
            .in2(_gnd_net_),
            .in3(N__46965),
            .lcout(\current_shift_inst.control_input_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_18_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_18_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_18_15_7 .LUT_INIT=16'b0011000000111111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_18_15_7  (
            .in0(_gnd_net_),
            .in1(N__47011),
            .in2(N__46991),
            .in3(N__46849),
            .lcout(\current_shift_inst.control_input_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_18_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_18_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_18_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_18_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47469),
            .lcout(\current_shift_inst.un4_control_input_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_18_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_18_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_18_16_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_18_16_1  (
            .in0(N__46796),
            .in1(N__47822),
            .in2(N__46406),
            .in3(N__47400),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_18_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_18_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_18_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_18_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48175),
            .lcout(\current_shift_inst.un4_control_input_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_18_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_18_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_18_16_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_18_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47821),
            .lcout(\current_shift_inst.un4_control_input_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_18_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_18_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_18_16_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_18_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47507),
            .lcout(\current_shift_inst.un4_control_input_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_18_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_18_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_18_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_18_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47860),
            .lcout(\current_shift_inst.un4_control_input_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_18_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_18_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_18_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_18_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47437),
            .lcout(\current_shift_inst.un4_control_input_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_18_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_18_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_18_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_18_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47893),
            .lcout(\current_shift_inst.un4_control_input_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_18_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_18_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_18_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_18_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47665),
            .lcout(\current_shift_inst.un4_control_input_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_18_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_18_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_18_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_18_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47578),
            .lcout(\current_shift_inst.un4_control_input_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_18_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_18_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_18_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_18_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47732),
            .lcout(\current_shift_inst.un4_control_input_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_18_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_18_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_18_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_18_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48220),
            .lcout(\current_shift_inst.un4_control_input_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_18_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_18_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_18_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_18_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48133),
            .lcout(\current_shift_inst.un4_control_input_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_18_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_18_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_18_17_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_18_17_5  (
            .in0(N__48530),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_18_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_18_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_18_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_18_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47701),
            .lcout(\current_shift_inst.un4_control_input_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_18_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_18_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_18_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_18_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47620),
            .lcout(\current_shift_inst.un4_control_input_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_18_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_18_18_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_18_18_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_18_18_0  (
            .in0(_gnd_net_),
            .in1(N__48741),
            .in2(N__48810),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_3 ),
            .ltout(),
            .carryin(bfn_18_18_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .clk(N__50195),
            .ce(N__48266),
            .sr(N__49651));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_18_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_18_18_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_18_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_18_18_1  (
            .in0(_gnd_net_),
            .in1(N__48717),
            .in2(N__48774),
            .in3(N__47452),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .clk(N__50195),
            .ce(N__48266),
            .sr(N__49651));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_18_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_18_18_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_18_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_18_18_2  (
            .in0(_gnd_net_),
            .in1(N__48742),
            .in2(N__48696),
            .in3(N__47410),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .clk(N__50195),
            .ce(N__48266),
            .sr(N__49651));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_18_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_18_18_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_18_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_18_18_3  (
            .in0(_gnd_net_),
            .in1(N__48718),
            .in2(N__48670),
            .in3(N__47866),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .clk(N__50195),
            .ce(N__48266),
            .sr(N__49651));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_18_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_18_18_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_18_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_18_18_4  (
            .in0(_gnd_net_),
            .in1(N__48636),
            .in2(N__48697),
            .in3(N__47836),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .clk(N__50195),
            .ce(N__48266),
            .sr(N__49651));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_18_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_18_18_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_18_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_18_18_5  (
            .in0(_gnd_net_),
            .in1(N__48666),
            .in2(N__48615),
            .in3(N__47803),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .clk(N__50195),
            .ce(N__48266),
            .sr(N__49651));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_18_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_18_18_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_18_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_18_18_6  (
            .in0(_gnd_net_),
            .in1(N__48637),
            .in2(N__49066),
            .in3(N__47758),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .clk(N__50195),
            .ce(N__48266),
            .sr(N__49651));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_18_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_18_18_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_18_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_18_18_7  (
            .in0(_gnd_net_),
            .in1(N__49038),
            .in2(N__48616),
            .in3(N__47716),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .clk(N__50195),
            .ce(N__48266),
            .sr(N__49651));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_18_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_18_19_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_18_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_18_19_0  (
            .in0(_gnd_net_),
            .in1(N__49065),
            .in2(N__49014),
            .in3(N__47677),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_11 ),
            .ltout(),
            .carryin(bfn_18_19_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .clk(N__50188),
            .ce(N__48265),
            .sr(N__49655));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_18_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_18_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_18_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_18_19_1  (
            .in0(_gnd_net_),
            .in1(N__49039),
            .in2(N__48987),
            .in3(N__47638),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .clk(N__50188),
            .ce(N__48265),
            .sr(N__49655));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_18_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_18_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_18_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_18_19_2  (
            .in0(_gnd_net_),
            .in1(N__48960),
            .in2(N__49015),
            .in3(N__47593),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .clk(N__50188),
            .ce(N__48265),
            .sr(N__49655));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_18_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_18_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_18_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_18_19_3  (
            .in0(_gnd_net_),
            .in1(N__48933),
            .in2(N__48988),
            .in3(N__47554),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .clk(N__50188),
            .ce(N__48265),
            .sr(N__49655));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_18_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_18_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_18_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_18_19_4  (
            .in0(_gnd_net_),
            .in1(N__48961),
            .in2(N__48906),
            .in3(N__48193),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .clk(N__50188),
            .ce(N__48265),
            .sr(N__49655));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_18_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_18_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_18_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_18_19_5  (
            .in0(_gnd_net_),
            .in1(N__48876),
            .in2(N__48937),
            .in3(N__48148),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .clk(N__50188),
            .ce(N__48265),
            .sr(N__49655));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_18_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_18_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_18_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_18_19_6  (
            .in0(_gnd_net_),
            .in1(N__49311),
            .in2(N__48907),
            .in3(N__48103),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .clk(N__50188),
            .ce(N__48265),
            .sr(N__49655));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_18_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_18_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_18_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_18_19_7  (
            .in0(_gnd_net_),
            .in1(N__48877),
            .in2(N__49285),
            .in3(N__48067),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .clk(N__50188),
            .ce(N__48265),
            .sr(N__49655));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_18_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_18_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_18_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_18_20_0  (
            .in0(_gnd_net_),
            .in1(N__49312),
            .in2(N__49254),
            .in3(N__48022),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_19 ),
            .ltout(),
            .carryin(bfn_18_20_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .clk(N__50182),
            .ce(N__48263),
            .sr(N__49661));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_18_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_18_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_18_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_18_20_1  (
            .in0(_gnd_net_),
            .in1(N__49284),
            .in2(N__49224),
            .in3(N__47989),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .clk(N__50182),
            .ce(N__48263),
            .sr(N__49661));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_18_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_18_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_18_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_18_20_2  (
            .in0(_gnd_net_),
            .in1(N__49194),
            .in2(N__49255),
            .in3(N__47956),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .clk(N__50182),
            .ce(N__48263),
            .sr(N__49661));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_18_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_18_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_18_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_18_20_3  (
            .in0(_gnd_net_),
            .in1(N__49170),
            .in2(N__49225),
            .in3(N__47908),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .clk(N__50182),
            .ce(N__48263),
            .sr(N__49661));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_18_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_18_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_18_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_18_20_4  (
            .in0(_gnd_net_),
            .in1(N__49195),
            .in2(N__49146),
            .in3(N__48541),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .clk(N__50182),
            .ce(N__48263),
            .sr(N__49661));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_18_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_18_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_18_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_18_20_5  (
            .in0(_gnd_net_),
            .in1(N__49171),
            .in2(N__49119),
            .in3(N__48505),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .clk(N__50182),
            .ce(N__48263),
            .sr(N__49661));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_18_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_18_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_18_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_18_20_6  (
            .in0(_gnd_net_),
            .in1(N__49092),
            .in2(N__49147),
            .in3(N__48469),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .clk(N__50182),
            .ce(N__48263),
            .sr(N__49661));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_18_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_18_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_18_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_18_20_7  (
            .in0(_gnd_net_),
            .in1(N__50631),
            .in2(N__49120),
            .in3(N__48430),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .clk(N__50182),
            .ce(N__48263),
            .sr(N__49661));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_18_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_18_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_18_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_18_21_0  (
            .in0(_gnd_net_),
            .in1(N__49093),
            .in2(N__50604),
            .in3(N__48385),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_27 ),
            .ltout(),
            .carryin(bfn_18_21_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .clk(N__50177),
            .ce(N__48262),
            .sr(N__49666));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_18_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_18_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_18_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_18_21_1  (
            .in0(_gnd_net_),
            .in1(N__50632),
            .in2(N__50577),
            .in3(N__48346),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .clk(N__50177),
            .ce(N__48262),
            .sr(N__49666));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_18_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_18_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_18_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_18_21_2  (
            .in0(_gnd_net_),
            .in1(N__50551),
            .in2(N__50605),
            .in3(N__48310),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .clk(N__50177),
            .ce(N__48262),
            .sr(N__49666));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_18_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_18_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_18_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_18_21_3  (
            .in0(_gnd_net_),
            .in1(N__50407),
            .in2(N__50578),
            .in3(N__48271),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ),
            .clk(N__50177),
            .ce(N__48262),
            .sr(N__49666));
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_18_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_18_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_18_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_18_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48238),
            .lcout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.counter_0_LC_18_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_0_LC_18_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_0_LC_18_22_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_0_LC_18_22_0  (
            .in0(N__50520),
            .in1(N__48797),
            .in2(_gnd_net_),
            .in3(N__48781),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_18_22_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_0 ),
            .clk(N__50172),
            .ce(N__50389),
            .sr(N__49673));
    defparam \current_shift_inst.timer_s1.counter_1_LC_18_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_1_LC_18_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_1_LC_18_22_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_1_LC_18_22_1  (
            .in0(N__50504),
            .in1(N__48764),
            .in2(_gnd_net_),
            .in3(N__48745),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_0 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_1 ),
            .clk(N__50172),
            .ce(N__50389),
            .sr(N__49673));
    defparam \current_shift_inst.timer_s1.counter_2_LC_18_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_2_LC_18_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_2_LC_18_22_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_2_LC_18_22_2  (
            .in0(N__50521),
            .in1(N__48735),
            .in2(_gnd_net_),
            .in3(N__48721),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_1 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_2 ),
            .clk(N__50172),
            .ce(N__50389),
            .sr(N__49673));
    defparam \current_shift_inst.timer_s1.counter_3_LC_18_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_3_LC_18_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_3_LC_18_22_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_3_LC_18_22_3  (
            .in0(N__50505),
            .in1(N__48716),
            .in2(_gnd_net_),
            .in3(N__48700),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_3 ),
            .clk(N__50172),
            .ce(N__50389),
            .sr(N__49673));
    defparam \current_shift_inst.timer_s1.counter_4_LC_18_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_4_LC_18_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_4_LC_18_22_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_4_LC_18_22_4  (
            .in0(N__50522),
            .in1(N__48689),
            .in2(_gnd_net_),
            .in3(N__48673),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_4 ),
            .clk(N__50172),
            .ce(N__50389),
            .sr(N__49673));
    defparam \current_shift_inst.timer_s1.counter_5_LC_18_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_5_LC_18_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_5_LC_18_22_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_5_LC_18_22_5  (
            .in0(N__50506),
            .in1(N__48662),
            .in2(_gnd_net_),
            .in3(N__48640),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_5 ),
            .clk(N__50172),
            .ce(N__50389),
            .sr(N__49673));
    defparam \current_shift_inst.timer_s1.counter_6_LC_18_22_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_6_LC_18_22_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_6_LC_18_22_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_6_LC_18_22_6  (
            .in0(N__50523),
            .in1(N__48635),
            .in2(_gnd_net_),
            .in3(N__48619),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_6 ),
            .clk(N__50172),
            .ce(N__50389),
            .sr(N__49673));
    defparam \current_shift_inst.timer_s1.counter_7_LC_18_22_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_7_LC_18_22_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_7_LC_18_22_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_7_LC_18_22_7  (
            .in0(N__50507),
            .in1(N__48603),
            .in2(_gnd_net_),
            .in3(N__48589),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_7 ),
            .clk(N__50172),
            .ce(N__50389),
            .sr(N__49673));
    defparam \current_shift_inst.timer_s1.counter_8_LC_18_23_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_8_LC_18_23_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_8_LC_18_23_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_8_LC_18_23_0  (
            .in0(N__50511),
            .in1(N__49061),
            .in2(_gnd_net_),
            .in3(N__49042),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_18_23_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_8 ),
            .clk(N__50166),
            .ce(N__50385),
            .sr(N__49680));
    defparam \current_shift_inst.timer_s1.counter_9_LC_18_23_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_9_LC_18_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_9_LC_18_23_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_9_LC_18_23_1  (
            .in0(N__50515),
            .in1(N__49037),
            .in2(_gnd_net_),
            .in3(N__49018),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_9 ),
            .clk(N__50166),
            .ce(N__50385),
            .sr(N__49680));
    defparam \current_shift_inst.timer_s1.counter_10_LC_18_23_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_10_LC_18_23_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_10_LC_18_23_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_10_LC_18_23_2  (
            .in0(N__50508),
            .in1(N__49007),
            .in2(_gnd_net_),
            .in3(N__48991),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_9 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_10 ),
            .clk(N__50166),
            .ce(N__50385),
            .sr(N__49680));
    defparam \current_shift_inst.timer_s1.counter_11_LC_18_23_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_11_LC_18_23_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_11_LC_18_23_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_11_LC_18_23_3  (
            .in0(N__50512),
            .in1(N__48980),
            .in2(_gnd_net_),
            .in3(N__48964),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_11 ),
            .clk(N__50166),
            .ce(N__50385),
            .sr(N__49680));
    defparam \current_shift_inst.timer_s1.counter_12_LC_18_23_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_12_LC_18_23_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_12_LC_18_23_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_12_LC_18_23_4  (
            .in0(N__50509),
            .in1(N__48954),
            .in2(_gnd_net_),
            .in3(N__48940),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_12 ),
            .clk(N__50166),
            .ce(N__50385),
            .sr(N__49680));
    defparam \current_shift_inst.timer_s1.counter_13_LC_18_23_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_13_LC_18_23_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_13_LC_18_23_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_13_LC_18_23_5  (
            .in0(N__50513),
            .in1(N__48926),
            .in2(_gnd_net_),
            .in3(N__48910),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_13 ),
            .clk(N__50166),
            .ce(N__50385),
            .sr(N__49680));
    defparam \current_shift_inst.timer_s1.counter_14_LC_18_23_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_14_LC_18_23_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_14_LC_18_23_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_14_LC_18_23_6  (
            .in0(N__50510),
            .in1(N__48894),
            .in2(_gnd_net_),
            .in3(N__48880),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_14 ),
            .clk(N__50166),
            .ce(N__50385),
            .sr(N__49680));
    defparam \current_shift_inst.timer_s1.counter_15_LC_18_23_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_15_LC_18_23_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_15_LC_18_23_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_15_LC_18_23_7  (
            .in0(N__50514),
            .in1(N__48875),
            .in2(_gnd_net_),
            .in3(N__48859),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_15 ),
            .clk(N__50166),
            .ce(N__50385),
            .sr(N__49680));
    defparam \current_shift_inst.timer_s1.counter_16_LC_18_24_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_16_LC_18_24_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_16_LC_18_24_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_16_LC_18_24_0  (
            .in0(N__50524),
            .in1(N__49304),
            .in2(_gnd_net_),
            .in3(N__49288),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_18_24_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_16 ),
            .clk(N__50162),
            .ce(N__50384),
            .sr(N__49687));
    defparam \current_shift_inst.timer_s1.counter_17_LC_18_24_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_17_LC_18_24_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_17_LC_18_24_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_17_LC_18_24_1  (
            .in0(N__50516),
            .in1(N__49274),
            .in2(_gnd_net_),
            .in3(N__49258),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_17 ),
            .clk(N__50162),
            .ce(N__50384),
            .sr(N__49687));
    defparam \current_shift_inst.timer_s1.counter_18_LC_18_24_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_18_LC_18_24_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_18_LC_18_24_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_18_LC_18_24_2  (
            .in0(N__50525),
            .in1(N__49242),
            .in2(_gnd_net_),
            .in3(N__49228),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_17 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_18 ),
            .clk(N__50162),
            .ce(N__50384),
            .sr(N__49687));
    defparam \current_shift_inst.timer_s1.counter_19_LC_18_24_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_19_LC_18_24_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_19_LC_18_24_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_19_LC_18_24_3  (
            .in0(N__50517),
            .in1(N__49212),
            .in2(_gnd_net_),
            .in3(N__49198),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_19 ),
            .clk(N__50162),
            .ce(N__50384),
            .sr(N__49687));
    defparam \current_shift_inst.timer_s1.counter_20_LC_18_24_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_20_LC_18_24_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_20_LC_18_24_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_20_LC_18_24_4  (
            .in0(N__50526),
            .in1(N__49188),
            .in2(_gnd_net_),
            .in3(N__49174),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_20 ),
            .clk(N__50162),
            .ce(N__50384),
            .sr(N__49687));
    defparam \current_shift_inst.timer_s1.counter_21_LC_18_24_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_21_LC_18_24_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_21_LC_18_24_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_21_LC_18_24_5  (
            .in0(N__50518),
            .in1(N__49164),
            .in2(_gnd_net_),
            .in3(N__49150),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_21 ),
            .clk(N__50162),
            .ce(N__50384),
            .sr(N__49687));
    defparam \current_shift_inst.timer_s1.counter_22_LC_18_24_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_22_LC_18_24_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_22_LC_18_24_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_22_LC_18_24_6  (
            .in0(N__50527),
            .in1(N__49139),
            .in2(_gnd_net_),
            .in3(N__49123),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_22 ),
            .clk(N__50162),
            .ce(N__50384),
            .sr(N__49687));
    defparam \current_shift_inst.timer_s1.counter_23_LC_18_24_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_23_LC_18_24_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_23_LC_18_24_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_23_LC_18_24_7  (
            .in0(N__50519),
            .in1(N__49112),
            .in2(_gnd_net_),
            .in3(N__49096),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_23 ),
            .clk(N__50162),
            .ce(N__50384),
            .sr(N__49687));
    defparam \current_shift_inst.timer_s1.counter_24_LC_18_25_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_24_LC_18_25_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_24_LC_18_25_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_24_LC_18_25_0  (
            .in0(N__50528),
            .in1(N__49085),
            .in2(_gnd_net_),
            .in3(N__49069),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_18_25_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_24 ),
            .clk(N__50159),
            .ce(N__50383),
            .sr(N__49692));
    defparam \current_shift_inst.timer_s1.counter_25_LC_18_25_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_25_LC_18_25_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_25_LC_18_25_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_25_LC_18_25_1  (
            .in0(N__50532),
            .in1(N__50624),
            .in2(_gnd_net_),
            .in3(N__50608),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_25 ),
            .clk(N__50159),
            .ce(N__50383),
            .sr(N__49692));
    defparam \current_shift_inst.timer_s1.counter_26_LC_18_25_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_26_LC_18_25_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_26_LC_18_25_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_26_LC_18_25_2  (
            .in0(N__50529),
            .in1(N__50597),
            .in2(_gnd_net_),
            .in3(N__50581),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_25 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_26 ),
            .clk(N__50159),
            .ce(N__50383),
            .sr(N__49692));
    defparam \current_shift_inst.timer_s1.counter_27_LC_18_25_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_27_LC_18_25_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_27_LC_18_25_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_27_LC_18_25_3  (
            .in0(N__50533),
            .in1(N__50570),
            .in2(_gnd_net_),
            .in3(N__50554),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_27 ),
            .clk(N__50159),
            .ce(N__50383),
            .sr(N__49692));
    defparam \current_shift_inst.timer_s1.counter_28_LC_18_25_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_28_LC_18_25_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_28_LC_18_25_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_28_LC_18_25_4  (
            .in0(N__50530),
            .in1(N__50550),
            .in2(_gnd_net_),
            .in3(N__50536),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_28 ),
            .clk(N__50159),
            .ce(N__50383),
            .sr(N__49692));
    defparam \current_shift_inst.timer_s1.counter_29_LC_18_25_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.counter_29_LC_18_25_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_29_LC_18_25_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \current_shift_inst.timer_s1.counter_29_LC_18_25_5  (
            .in0(N__50403),
            .in1(N__50531),
            .in2(_gnd_net_),
            .in3(N__50410),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50159),
            .ce(N__50383),
            .sr(N__49692));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_20_12_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_20_12_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_20_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_20_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50332),
            .lcout(\delay_measurement_inst.elapsed_time_tr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50249),
            .ce(N__49816),
            .sr(N__49620));
endmodule // MAIN
