-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jul 24 2025 22:26:30

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "MAIN" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of MAIN
entity MAIN is
port (
    s3_phy : out std_logic;
    il_min_comp2 : in std_logic;
    il_max_comp1 : in std_logic;
    s1_phy : out std_logic;
    reset : in std_logic;
    il_min_comp1 : in std_logic;
    delay_tr_input : in std_logic;
    s4_phy : out std_logic;
    rgb_g : out std_logic;
    start_stop : in std_logic;
    s2_phy : out std_logic;
    rgb_r : out std_logic;
    rgb_b : out std_logic;
    pwm_output : out std_logic;
    il_max_comp2 : in std_logic;
    delay_hc_input : in std_logic);
end MAIN;

-- Architecture of MAIN
-- View name is \INTERFACE\
architecture \INTERFACE\ of MAIN is

signal \N__48680\ : std_logic;
signal \N__48679\ : std_logic;
signal \N__48678\ : std_logic;
signal \N__48669\ : std_logic;
signal \N__48668\ : std_logic;
signal \N__48667\ : std_logic;
signal \N__48660\ : std_logic;
signal \N__48659\ : std_logic;
signal \N__48658\ : std_logic;
signal \N__48651\ : std_logic;
signal \N__48650\ : std_logic;
signal \N__48649\ : std_logic;
signal \N__48642\ : std_logic;
signal \N__48641\ : std_logic;
signal \N__48640\ : std_logic;
signal \N__48633\ : std_logic;
signal \N__48632\ : std_logic;
signal \N__48631\ : std_logic;
signal \N__48624\ : std_logic;
signal \N__48623\ : std_logic;
signal \N__48622\ : std_logic;
signal \N__48615\ : std_logic;
signal \N__48614\ : std_logic;
signal \N__48613\ : std_logic;
signal \N__48606\ : std_logic;
signal \N__48605\ : std_logic;
signal \N__48604\ : std_logic;
signal \N__48597\ : std_logic;
signal \N__48596\ : std_logic;
signal \N__48595\ : std_logic;
signal \N__48588\ : std_logic;
signal \N__48587\ : std_logic;
signal \N__48586\ : std_logic;
signal \N__48579\ : std_logic;
signal \N__48578\ : std_logic;
signal \N__48577\ : std_logic;
signal \N__48570\ : std_logic;
signal \N__48569\ : std_logic;
signal \N__48568\ : std_logic;
signal \N__48551\ : std_logic;
signal \N__48550\ : std_logic;
signal \N__48547\ : std_logic;
signal \N__48544\ : std_logic;
signal \N__48543\ : std_logic;
signal \N__48538\ : std_logic;
signal \N__48535\ : std_logic;
signal \N__48532\ : std_logic;
signal \N__48529\ : std_logic;
signal \N__48524\ : std_logic;
signal \N__48521\ : std_logic;
signal \N__48520\ : std_logic;
signal \N__48517\ : std_logic;
signal \N__48514\ : std_logic;
signal \N__48509\ : std_logic;
signal \N__48506\ : std_logic;
signal \N__48505\ : std_logic;
signal \N__48504\ : std_logic;
signal \N__48499\ : std_logic;
signal \N__48496\ : std_logic;
signal \N__48495\ : std_logic;
signal \N__48494\ : std_logic;
signal \N__48491\ : std_logic;
signal \N__48488\ : std_logic;
signal \N__48485\ : std_logic;
signal \N__48482\ : std_logic;
signal \N__48479\ : std_logic;
signal \N__48472\ : std_logic;
signal \N__48467\ : std_logic;
signal \N__48466\ : std_logic;
signal \N__48463\ : std_logic;
signal \N__48460\ : std_logic;
signal \N__48459\ : std_logic;
signal \N__48454\ : std_logic;
signal \N__48451\ : std_logic;
signal \N__48446\ : std_logic;
signal \N__48443\ : std_logic;
signal \N__48442\ : std_logic;
signal \N__48439\ : std_logic;
signal \N__48438\ : std_logic;
signal \N__48435\ : std_logic;
signal \N__48432\ : std_logic;
signal \N__48429\ : std_logic;
signal \N__48426\ : std_logic;
signal \N__48423\ : std_logic;
signal \N__48420\ : std_logic;
signal \N__48417\ : std_logic;
signal \N__48410\ : std_logic;
signal \N__48409\ : std_logic;
signal \N__48406\ : std_logic;
signal \N__48403\ : std_logic;
signal \N__48402\ : std_logic;
signal \N__48397\ : std_logic;
signal \N__48394\ : std_logic;
signal \N__48389\ : std_logic;
signal \N__48388\ : std_logic;
signal \N__48385\ : std_logic;
signal \N__48382\ : std_logic;
signal \N__48377\ : std_logic;
signal \N__48374\ : std_logic;
signal \N__48373\ : std_logic;
signal \N__48370\ : std_logic;
signal \N__48367\ : std_logic;
signal \N__48366\ : std_logic;
signal \N__48361\ : std_logic;
signal \N__48358\ : std_logic;
signal \N__48357\ : std_logic;
signal \N__48352\ : std_logic;
signal \N__48349\ : std_logic;
signal \N__48346\ : std_logic;
signal \N__48343\ : std_logic;
signal \N__48338\ : std_logic;
signal \N__48335\ : std_logic;
signal \N__48334\ : std_logic;
signal \N__48331\ : std_logic;
signal \N__48328\ : std_logic;
signal \N__48327\ : std_logic;
signal \N__48322\ : std_logic;
signal \N__48319\ : std_logic;
signal \N__48318\ : std_logic;
signal \N__48313\ : std_logic;
signal \N__48310\ : std_logic;
signal \N__48307\ : std_logic;
signal \N__48304\ : std_logic;
signal \N__48299\ : std_logic;
signal \N__48296\ : std_logic;
signal \N__48293\ : std_logic;
signal \N__48290\ : std_logic;
signal \N__48287\ : std_logic;
signal \N__48284\ : std_logic;
signal \N__48283\ : std_logic;
signal \N__48282\ : std_logic;
signal \N__48281\ : std_logic;
signal \N__48280\ : std_logic;
signal \N__48279\ : std_logic;
signal \N__48278\ : std_logic;
signal \N__48275\ : std_logic;
signal \N__48274\ : std_logic;
signal \N__48273\ : std_logic;
signal \N__48270\ : std_logic;
signal \N__48267\ : std_logic;
signal \N__48266\ : std_logic;
signal \N__48265\ : std_logic;
signal \N__48262\ : std_logic;
signal \N__48261\ : std_logic;
signal \N__48260\ : std_logic;
signal \N__48259\ : std_logic;
signal \N__48258\ : std_logic;
signal \N__48257\ : std_logic;
signal \N__48254\ : std_logic;
signal \N__48253\ : std_logic;
signal \N__48252\ : std_logic;
signal \N__48247\ : std_logic;
signal \N__48240\ : std_logic;
signal \N__48231\ : std_logic;
signal \N__48228\ : std_logic;
signal \N__48223\ : std_logic;
signal \N__48220\ : std_logic;
signal \N__48217\ : std_logic;
signal \N__48216\ : std_logic;
signal \N__48215\ : std_logic;
signal \N__48212\ : std_logic;
signal \N__48211\ : std_logic;
signal \N__48208\ : std_logic;
signal \N__48203\ : std_logic;
signal \N__48196\ : std_logic;
signal \N__48191\ : std_logic;
signal \N__48178\ : std_logic;
signal \N__48173\ : std_logic;
signal \N__48168\ : std_logic;
signal \N__48165\ : std_logic;
signal \N__48162\ : std_logic;
signal \N__48155\ : std_logic;
signal \N__48154\ : std_logic;
signal \N__48151\ : std_logic;
signal \N__48148\ : std_logic;
signal \N__48147\ : std_logic;
signal \N__48144\ : std_logic;
signal \N__48141\ : std_logic;
signal \N__48138\ : std_logic;
signal \N__48133\ : std_logic;
signal \N__48130\ : std_logic;
signal \N__48125\ : std_logic;
signal \N__48122\ : std_logic;
signal \N__48121\ : std_logic;
signal \N__48120\ : std_logic;
signal \N__48119\ : std_logic;
signal \N__48114\ : std_logic;
signal \N__48111\ : std_logic;
signal \N__48108\ : std_logic;
signal \N__48107\ : std_logic;
signal \N__48106\ : std_logic;
signal \N__48103\ : std_logic;
signal \N__48100\ : std_logic;
signal \N__48097\ : std_logic;
signal \N__48092\ : std_logic;
signal \N__48091\ : std_logic;
signal \N__48090\ : std_logic;
signal \N__48081\ : std_logic;
signal \N__48080\ : std_logic;
signal \N__48075\ : std_logic;
signal \N__48072\ : std_logic;
signal \N__48069\ : std_logic;
signal \N__48066\ : std_logic;
signal \N__48059\ : std_logic;
signal \N__48056\ : std_logic;
signal \N__48055\ : std_logic;
signal \N__48054\ : std_logic;
signal \N__48051\ : std_logic;
signal \N__48048\ : std_logic;
signal \N__48045\ : std_logic;
signal \N__48044\ : std_logic;
signal \N__48041\ : std_logic;
signal \N__48038\ : std_logic;
signal \N__48035\ : std_logic;
signal \N__48032\ : std_logic;
signal \N__48027\ : std_logic;
signal \N__48024\ : std_logic;
signal \N__48021\ : std_logic;
signal \N__48018\ : std_logic;
signal \N__48013\ : std_logic;
signal \N__48008\ : std_logic;
signal \N__48007\ : std_logic;
signal \N__48006\ : std_logic;
signal \N__48005\ : std_logic;
signal \N__48004\ : std_logic;
signal \N__48003\ : std_logic;
signal \N__48002\ : std_logic;
signal \N__48001\ : std_logic;
signal \N__48000\ : std_logic;
signal \N__47999\ : std_logic;
signal \N__47998\ : std_logic;
signal \N__47997\ : std_logic;
signal \N__47996\ : std_logic;
signal \N__47995\ : std_logic;
signal \N__47994\ : std_logic;
signal \N__47993\ : std_logic;
signal \N__47992\ : std_logic;
signal \N__47991\ : std_logic;
signal \N__47990\ : std_logic;
signal \N__47989\ : std_logic;
signal \N__47988\ : std_logic;
signal \N__47987\ : std_logic;
signal \N__47986\ : std_logic;
signal \N__47985\ : std_logic;
signal \N__47984\ : std_logic;
signal \N__47983\ : std_logic;
signal \N__47982\ : std_logic;
signal \N__47981\ : std_logic;
signal \N__47980\ : std_logic;
signal \N__47979\ : std_logic;
signal \N__47978\ : std_logic;
signal \N__47977\ : std_logic;
signal \N__47976\ : std_logic;
signal \N__47975\ : std_logic;
signal \N__47974\ : std_logic;
signal \N__47973\ : std_logic;
signal \N__47972\ : std_logic;
signal \N__47971\ : std_logic;
signal \N__47970\ : std_logic;
signal \N__47969\ : std_logic;
signal \N__47968\ : std_logic;
signal \N__47967\ : std_logic;
signal \N__47966\ : std_logic;
signal \N__47965\ : std_logic;
signal \N__47964\ : std_logic;
signal \N__47963\ : std_logic;
signal \N__47962\ : std_logic;
signal \N__47961\ : std_logic;
signal \N__47960\ : std_logic;
signal \N__47959\ : std_logic;
signal \N__47958\ : std_logic;
signal \N__47957\ : std_logic;
signal \N__47956\ : std_logic;
signal \N__47955\ : std_logic;
signal \N__47954\ : std_logic;
signal \N__47953\ : std_logic;
signal \N__47952\ : std_logic;
signal \N__47951\ : std_logic;
signal \N__47950\ : std_logic;
signal \N__47949\ : std_logic;
signal \N__47948\ : std_logic;
signal \N__47947\ : std_logic;
signal \N__47946\ : std_logic;
signal \N__47945\ : std_logic;
signal \N__47944\ : std_logic;
signal \N__47943\ : std_logic;
signal \N__47942\ : std_logic;
signal \N__47941\ : std_logic;
signal \N__47940\ : std_logic;
signal \N__47939\ : std_logic;
signal \N__47938\ : std_logic;
signal \N__47937\ : std_logic;
signal \N__47936\ : std_logic;
signal \N__47935\ : std_logic;
signal \N__47934\ : std_logic;
signal \N__47933\ : std_logic;
signal \N__47932\ : std_logic;
signal \N__47931\ : std_logic;
signal \N__47930\ : std_logic;
signal \N__47929\ : std_logic;
signal \N__47928\ : std_logic;
signal \N__47927\ : std_logic;
signal \N__47926\ : std_logic;
signal \N__47925\ : std_logic;
signal \N__47924\ : std_logic;
signal \N__47923\ : std_logic;
signal \N__47922\ : std_logic;
signal \N__47921\ : std_logic;
signal \N__47920\ : std_logic;
signal \N__47919\ : std_logic;
signal \N__47918\ : std_logic;
signal \N__47917\ : std_logic;
signal \N__47916\ : std_logic;
signal \N__47915\ : std_logic;
signal \N__47914\ : std_logic;
signal \N__47913\ : std_logic;
signal \N__47912\ : std_logic;
signal \N__47911\ : std_logic;
signal \N__47910\ : std_logic;
signal \N__47909\ : std_logic;
signal \N__47908\ : std_logic;
signal \N__47907\ : std_logic;
signal \N__47906\ : std_logic;
signal \N__47905\ : std_logic;
signal \N__47904\ : std_logic;
signal \N__47903\ : std_logic;
signal \N__47902\ : std_logic;
signal \N__47901\ : std_logic;
signal \N__47900\ : std_logic;
signal \N__47899\ : std_logic;
signal \N__47898\ : std_logic;
signal \N__47897\ : std_logic;
signal \N__47896\ : std_logic;
signal \N__47895\ : std_logic;
signal \N__47894\ : std_logic;
signal \N__47893\ : std_logic;
signal \N__47892\ : std_logic;
signal \N__47891\ : std_logic;
signal \N__47890\ : std_logic;
signal \N__47889\ : std_logic;
signal \N__47888\ : std_logic;
signal \N__47887\ : std_logic;
signal \N__47886\ : std_logic;
signal \N__47885\ : std_logic;
signal \N__47884\ : std_logic;
signal \N__47883\ : std_logic;
signal \N__47882\ : std_logic;
signal \N__47881\ : std_logic;
signal \N__47880\ : std_logic;
signal \N__47879\ : std_logic;
signal \N__47878\ : std_logic;
signal \N__47877\ : std_logic;
signal \N__47876\ : std_logic;
signal \N__47875\ : std_logic;
signal \N__47874\ : std_logic;
signal \N__47873\ : std_logic;
signal \N__47872\ : std_logic;
signal \N__47871\ : std_logic;
signal \N__47870\ : std_logic;
signal \N__47869\ : std_logic;
signal \N__47868\ : std_logic;
signal \N__47867\ : std_logic;
signal \N__47866\ : std_logic;
signal \N__47865\ : std_logic;
signal \N__47864\ : std_logic;
signal \N__47863\ : std_logic;
signal \N__47862\ : std_logic;
signal \N__47861\ : std_logic;
signal \N__47860\ : std_logic;
signal \N__47859\ : std_logic;
signal \N__47858\ : std_logic;
signal \N__47857\ : std_logic;
signal \N__47856\ : std_logic;
signal \N__47855\ : std_logic;
signal \N__47854\ : std_logic;
signal \N__47853\ : std_logic;
signal \N__47852\ : std_logic;
signal \N__47851\ : std_logic;
signal \N__47850\ : std_logic;
signal \N__47849\ : std_logic;
signal \N__47848\ : std_logic;
signal \N__47847\ : std_logic;
signal \N__47522\ : std_logic;
signal \N__47519\ : std_logic;
signal \N__47518\ : std_logic;
signal \N__47515\ : std_logic;
signal \N__47512\ : std_logic;
signal \N__47511\ : std_logic;
signal \N__47508\ : std_logic;
signal \N__47505\ : std_logic;
signal \N__47502\ : std_logic;
signal \N__47499\ : std_logic;
signal \N__47496\ : std_logic;
signal \N__47493\ : std_logic;
signal \N__47492\ : std_logic;
signal \N__47491\ : std_logic;
signal \N__47490\ : std_logic;
signal \N__47483\ : std_logic;
signal \N__47480\ : std_logic;
signal \N__47477\ : std_logic;
signal \N__47474\ : std_logic;
signal \N__47465\ : std_logic;
signal \N__47464\ : std_logic;
signal \N__47463\ : std_logic;
signal \N__47462\ : std_logic;
signal \N__47461\ : std_logic;
signal \N__47460\ : std_logic;
signal \N__47459\ : std_logic;
signal \N__47456\ : std_logic;
signal \N__47453\ : std_logic;
signal \N__47450\ : std_logic;
signal \N__47447\ : std_logic;
signal \N__47444\ : std_logic;
signal \N__47441\ : std_logic;
signal \N__47438\ : std_logic;
signal \N__47435\ : std_logic;
signal \N__47432\ : std_logic;
signal \N__47429\ : std_logic;
signal \N__47426\ : std_logic;
signal \N__47423\ : std_logic;
signal \N__47422\ : std_logic;
signal \N__47421\ : std_logic;
signal \N__47418\ : std_logic;
signal \N__47417\ : std_logic;
signal \N__47416\ : std_logic;
signal \N__47415\ : std_logic;
signal \N__47414\ : std_logic;
signal \N__47413\ : std_logic;
signal \N__47412\ : std_logic;
signal \N__47411\ : std_logic;
signal \N__47410\ : std_logic;
signal \N__47409\ : std_logic;
signal \N__47408\ : std_logic;
signal \N__47407\ : std_logic;
signal \N__47406\ : std_logic;
signal \N__47405\ : std_logic;
signal \N__47404\ : std_logic;
signal \N__47403\ : std_logic;
signal \N__47402\ : std_logic;
signal \N__47401\ : std_logic;
signal \N__47400\ : std_logic;
signal \N__47399\ : std_logic;
signal \N__47398\ : std_logic;
signal \N__47397\ : std_logic;
signal \N__47396\ : std_logic;
signal \N__47395\ : std_logic;
signal \N__47394\ : std_logic;
signal \N__47393\ : std_logic;
signal \N__47392\ : std_logic;
signal \N__47391\ : std_logic;
signal \N__47390\ : std_logic;
signal \N__47389\ : std_logic;
signal \N__47388\ : std_logic;
signal \N__47387\ : std_logic;
signal \N__47386\ : std_logic;
signal \N__47385\ : std_logic;
signal \N__47384\ : std_logic;
signal \N__47383\ : std_logic;
signal \N__47382\ : std_logic;
signal \N__47381\ : std_logic;
signal \N__47380\ : std_logic;
signal \N__47379\ : std_logic;
signal \N__47378\ : std_logic;
signal \N__47377\ : std_logic;
signal \N__47376\ : std_logic;
signal \N__47375\ : std_logic;
signal \N__47374\ : std_logic;
signal \N__47373\ : std_logic;
signal \N__47372\ : std_logic;
signal \N__47371\ : std_logic;
signal \N__47370\ : std_logic;
signal \N__47369\ : std_logic;
signal \N__47368\ : std_logic;
signal \N__47367\ : std_logic;
signal \N__47366\ : std_logic;
signal \N__47365\ : std_logic;
signal \N__47364\ : std_logic;
signal \N__47363\ : std_logic;
signal \N__47362\ : std_logic;
signal \N__47361\ : std_logic;
signal \N__47360\ : std_logic;
signal \N__47359\ : std_logic;
signal \N__47358\ : std_logic;
signal \N__47357\ : std_logic;
signal \N__47356\ : std_logic;
signal \N__47355\ : std_logic;
signal \N__47354\ : std_logic;
signal \N__47353\ : std_logic;
signal \N__47352\ : std_logic;
signal \N__47351\ : std_logic;
signal \N__47350\ : std_logic;
signal \N__47349\ : std_logic;
signal \N__47348\ : std_logic;
signal \N__47347\ : std_logic;
signal \N__47346\ : std_logic;
signal \N__47345\ : std_logic;
signal \N__47344\ : std_logic;
signal \N__47343\ : std_logic;
signal \N__47342\ : std_logic;
signal \N__47341\ : std_logic;
signal \N__47340\ : std_logic;
signal \N__47339\ : std_logic;
signal \N__47338\ : std_logic;
signal \N__47337\ : std_logic;
signal \N__47336\ : std_logic;
signal \N__47335\ : std_logic;
signal \N__47332\ : std_logic;
signal \N__47331\ : std_logic;
signal \N__47330\ : std_logic;
signal \N__47329\ : std_logic;
signal \N__47328\ : std_logic;
signal \N__47327\ : std_logic;
signal \N__47326\ : std_logic;
signal \N__47325\ : std_logic;
signal \N__47324\ : std_logic;
signal \N__47323\ : std_logic;
signal \N__47322\ : std_logic;
signal \N__47321\ : std_logic;
signal \N__47320\ : std_logic;
signal \N__47319\ : std_logic;
signal \N__47318\ : std_logic;
signal \N__47317\ : std_logic;
signal \N__47316\ : std_logic;
signal \N__47315\ : std_logic;
signal \N__47314\ : std_logic;
signal \N__47313\ : std_logic;
signal \N__47312\ : std_logic;
signal \N__47311\ : std_logic;
signal \N__47310\ : std_logic;
signal \N__47309\ : std_logic;
signal \N__47308\ : std_logic;
signal \N__47307\ : std_logic;
signal \N__47306\ : std_logic;
signal \N__47305\ : std_logic;
signal \N__47304\ : std_logic;
signal \N__47303\ : std_logic;
signal \N__47302\ : std_logic;
signal \N__47301\ : std_logic;
signal \N__47300\ : std_logic;
signal \N__47299\ : std_logic;
signal \N__47298\ : std_logic;
signal \N__47297\ : std_logic;
signal \N__47296\ : std_logic;
signal \N__47295\ : std_logic;
signal \N__47294\ : std_logic;
signal \N__47293\ : std_logic;
signal \N__47292\ : std_logic;
signal \N__47291\ : std_logic;
signal \N__47290\ : std_logic;
signal \N__47289\ : std_logic;
signal \N__47288\ : std_logic;
signal \N__47287\ : std_logic;
signal \N__47286\ : std_logic;
signal \N__47283\ : std_logic;
signal \N__47280\ : std_logic;
signal \N__47279\ : std_logic;
signal \N__47278\ : std_logic;
signal \N__47277\ : std_logic;
signal \N__47276\ : std_logic;
signal \N__47275\ : std_logic;
signal \N__47274\ : std_logic;
signal \N__47273\ : std_logic;
signal \N__47272\ : std_logic;
signal \N__46979\ : std_logic;
signal \N__46976\ : std_logic;
signal \N__46973\ : std_logic;
signal \N__46970\ : std_logic;
signal \N__46969\ : std_logic;
signal \N__46966\ : std_logic;
signal \N__46963\ : std_logic;
signal \N__46960\ : std_logic;
signal \N__46957\ : std_logic;
signal \N__46954\ : std_logic;
signal \N__46951\ : std_logic;
signal \N__46946\ : std_logic;
signal \N__46945\ : std_logic;
signal \N__46942\ : std_logic;
signal \N__46941\ : std_logic;
signal \N__46938\ : std_logic;
signal \N__46935\ : std_logic;
signal \N__46932\ : std_logic;
signal \N__46929\ : std_logic;
signal \N__46924\ : std_logic;
signal \N__46919\ : std_logic;
signal \N__46916\ : std_logic;
signal \N__46915\ : std_logic;
signal \N__46914\ : std_logic;
signal \N__46911\ : std_logic;
signal \N__46906\ : std_logic;
signal \N__46903\ : std_logic;
signal \N__46900\ : std_logic;
signal \N__46897\ : std_logic;
signal \N__46894\ : std_logic;
signal \N__46889\ : std_logic;
signal \N__46888\ : std_logic;
signal \N__46885\ : std_logic;
signal \N__46884\ : std_logic;
signal \N__46881\ : std_logic;
signal \N__46878\ : std_logic;
signal \N__46875\ : std_logic;
signal \N__46872\ : std_logic;
signal \N__46867\ : std_logic;
signal \N__46864\ : std_logic;
signal \N__46861\ : std_logic;
signal \N__46858\ : std_logic;
signal \N__46855\ : std_logic;
signal \N__46850\ : std_logic;
signal \N__46849\ : std_logic;
signal \N__46846\ : std_logic;
signal \N__46843\ : std_logic;
signal \N__46840\ : std_logic;
signal \N__46837\ : std_logic;
signal \N__46834\ : std_logic;
signal \N__46831\ : std_logic;
signal \N__46828\ : std_logic;
signal \N__46823\ : std_logic;
signal \N__46822\ : std_logic;
signal \N__46819\ : std_logic;
signal \N__46816\ : std_logic;
signal \N__46815\ : std_logic;
signal \N__46812\ : std_logic;
signal \N__46809\ : std_logic;
signal \N__46806\ : std_logic;
signal \N__46803\ : std_logic;
signal \N__46798\ : std_logic;
signal \N__46795\ : std_logic;
signal \N__46792\ : std_logic;
signal \N__46787\ : std_logic;
signal \N__46786\ : std_logic;
signal \N__46783\ : std_logic;
signal \N__46780\ : std_logic;
signal \N__46777\ : std_logic;
signal \N__46774\ : std_logic;
signal \N__46771\ : std_logic;
signal \N__46768\ : std_logic;
signal \N__46763\ : std_logic;
signal \N__46760\ : std_logic;
signal \N__46759\ : std_logic;
signal \N__46758\ : std_logic;
signal \N__46755\ : std_logic;
signal \N__46752\ : std_logic;
signal \N__46749\ : std_logic;
signal \N__46742\ : std_logic;
signal \N__46739\ : std_logic;
signal \N__46736\ : std_logic;
signal \N__46735\ : std_logic;
signal \N__46734\ : std_logic;
signal \N__46731\ : std_logic;
signal \N__46728\ : std_logic;
signal \N__46725\ : std_logic;
signal \N__46722\ : std_logic;
signal \N__46719\ : std_logic;
signal \N__46716\ : std_logic;
signal \N__46713\ : std_logic;
signal \N__46710\ : std_logic;
signal \N__46707\ : std_logic;
signal \N__46700\ : std_logic;
signal \N__46699\ : std_logic;
signal \N__46696\ : std_logic;
signal \N__46693\ : std_logic;
signal \N__46690\ : std_logic;
signal \N__46687\ : std_logic;
signal \N__46682\ : std_logic;
signal \N__46679\ : std_logic;
signal \N__46678\ : std_logic;
signal \N__46675\ : std_logic;
signal \N__46674\ : std_logic;
signal \N__46671\ : std_logic;
signal \N__46668\ : std_logic;
signal \N__46665\ : std_logic;
signal \N__46662\ : std_logic;
signal \N__46655\ : std_logic;
signal \N__46652\ : std_logic;
signal \N__46649\ : std_logic;
signal \N__46648\ : std_logic;
signal \N__46647\ : std_logic;
signal \N__46644\ : std_logic;
signal \N__46641\ : std_logic;
signal \N__46638\ : std_logic;
signal \N__46637\ : std_logic;
signal \N__46630\ : std_logic;
signal \N__46627\ : std_logic;
signal \N__46622\ : std_logic;
signal \N__46619\ : std_logic;
signal \N__46616\ : std_logic;
signal \N__46615\ : std_logic;
signal \N__46614\ : std_logic;
signal \N__46611\ : std_logic;
signal \N__46608\ : std_logic;
signal \N__46605\ : std_logic;
signal \N__46598\ : std_logic;
signal \N__46595\ : std_logic;
signal \N__46592\ : std_logic;
signal \N__46591\ : std_logic;
signal \N__46588\ : std_logic;
signal \N__46585\ : std_logic;
signal \N__46582\ : std_logic;
signal \N__46579\ : std_logic;
signal \N__46576\ : std_logic;
signal \N__46573\ : std_logic;
signal \N__46568\ : std_logic;
signal \N__46565\ : std_logic;
signal \N__46564\ : std_logic;
signal \N__46563\ : std_logic;
signal \N__46560\ : std_logic;
signal \N__46557\ : std_logic;
signal \N__46554\ : std_logic;
signal \N__46547\ : std_logic;
signal \N__46544\ : std_logic;
signal \N__46541\ : std_logic;
signal \N__46540\ : std_logic;
signal \N__46539\ : std_logic;
signal \N__46538\ : std_logic;
signal \N__46537\ : std_logic;
signal \N__46536\ : std_logic;
signal \N__46535\ : std_logic;
signal \N__46534\ : std_logic;
signal \N__46525\ : std_logic;
signal \N__46516\ : std_logic;
signal \N__46513\ : std_logic;
signal \N__46510\ : std_logic;
signal \N__46507\ : std_logic;
signal \N__46504\ : std_logic;
signal \N__46499\ : std_logic;
signal \N__46498\ : std_logic;
signal \N__46497\ : std_logic;
signal \N__46490\ : std_logic;
signal \N__46489\ : std_logic;
signal \N__46488\ : std_logic;
signal \N__46487\ : std_logic;
signal \N__46484\ : std_logic;
signal \N__46477\ : std_logic;
signal \N__46472\ : std_logic;
signal \N__46469\ : std_logic;
signal \N__46468\ : std_logic;
signal \N__46467\ : std_logic;
signal \N__46464\ : std_logic;
signal \N__46461\ : std_logic;
signal \N__46458\ : std_logic;
signal \N__46455\ : std_logic;
signal \N__46452\ : std_logic;
signal \N__46449\ : std_logic;
signal \N__46444\ : std_logic;
signal \N__46441\ : std_logic;
signal \N__46438\ : std_logic;
signal \N__46433\ : std_logic;
signal \N__46432\ : std_logic;
signal \N__46429\ : std_logic;
signal \N__46426\ : std_logic;
signal \N__46423\ : std_logic;
signal \N__46422\ : std_logic;
signal \N__46419\ : std_logic;
signal \N__46416\ : std_logic;
signal \N__46413\ : std_logic;
signal \N__46410\ : std_logic;
signal \N__46405\ : std_logic;
signal \N__46402\ : std_logic;
signal \N__46399\ : std_logic;
signal \N__46394\ : std_logic;
signal \N__46391\ : std_logic;
signal \N__46388\ : std_logic;
signal \N__46385\ : std_logic;
signal \N__46382\ : std_logic;
signal \N__46379\ : std_logic;
signal \N__46376\ : std_logic;
signal \N__46375\ : std_logic;
signal \N__46372\ : std_logic;
signal \N__46369\ : std_logic;
signal \N__46364\ : std_logic;
signal \N__46363\ : std_logic;
signal \N__46358\ : std_logic;
signal \N__46355\ : std_logic;
signal \N__46352\ : std_logic;
signal \N__46349\ : std_logic;
signal \N__46348\ : std_logic;
signal \N__46345\ : std_logic;
signal \N__46342\ : std_logic;
signal \N__46341\ : std_logic;
signal \N__46340\ : std_logic;
signal \N__46337\ : std_logic;
signal \N__46334\ : std_logic;
signal \N__46329\ : std_logic;
signal \N__46322\ : std_logic;
signal \N__46319\ : std_logic;
signal \N__46318\ : std_logic;
signal \N__46317\ : std_logic;
signal \N__46314\ : std_logic;
signal \N__46313\ : std_logic;
signal \N__46312\ : std_logic;
signal \N__46309\ : std_logic;
signal \N__46306\ : std_logic;
signal \N__46303\ : std_logic;
signal \N__46298\ : std_logic;
signal \N__46295\ : std_logic;
signal \N__46288\ : std_logic;
signal \N__46285\ : std_logic;
signal \N__46282\ : std_logic;
signal \N__46277\ : std_logic;
signal \N__46276\ : std_logic;
signal \N__46275\ : std_logic;
signal \N__46274\ : std_logic;
signal \N__46273\ : std_logic;
signal \N__46272\ : std_logic;
signal \N__46269\ : std_logic;
signal \N__46266\ : std_logic;
signal \N__46263\ : std_logic;
signal \N__46260\ : std_logic;
signal \N__46255\ : std_logic;
signal \N__46254\ : std_logic;
signal \N__46251\ : std_logic;
signal \N__46248\ : std_logic;
signal \N__46241\ : std_logic;
signal \N__46238\ : std_logic;
signal \N__46235\ : std_logic;
signal \N__46232\ : std_logic;
signal \N__46229\ : std_logic;
signal \N__46226\ : std_logic;
signal \N__46217\ : std_logic;
signal \N__46214\ : std_logic;
signal \N__46213\ : std_logic;
signal \N__46210\ : std_logic;
signal \N__46207\ : std_logic;
signal \N__46206\ : std_logic;
signal \N__46205\ : std_logic;
signal \N__46204\ : std_logic;
signal \N__46201\ : std_logic;
signal \N__46198\ : std_logic;
signal \N__46191\ : std_logic;
signal \N__46184\ : std_logic;
signal \N__46183\ : std_logic;
signal \N__46182\ : std_logic;
signal \N__46181\ : std_logic;
signal \N__46180\ : std_logic;
signal \N__46179\ : std_logic;
signal \N__46178\ : std_logic;
signal \N__46177\ : std_logic;
signal \N__46174\ : std_logic;
signal \N__46173\ : std_logic;
signal \N__46170\ : std_logic;
signal \N__46167\ : std_logic;
signal \N__46164\ : std_logic;
signal \N__46161\ : std_logic;
signal \N__46156\ : std_logic;
signal \N__46155\ : std_logic;
signal \N__46152\ : std_logic;
signal \N__46149\ : std_logic;
signal \N__46146\ : std_logic;
signal \N__46143\ : std_logic;
signal \N__46140\ : std_logic;
signal \N__46137\ : std_logic;
signal \N__46132\ : std_logic;
signal \N__46127\ : std_logic;
signal \N__46120\ : std_logic;
signal \N__46115\ : std_logic;
signal \N__46110\ : std_logic;
signal \N__46105\ : std_logic;
signal \N__46102\ : std_logic;
signal \N__46099\ : std_logic;
signal \N__46096\ : std_logic;
signal \N__46091\ : std_logic;
signal \N__46090\ : std_logic;
signal \N__46087\ : std_logic;
signal \N__46084\ : std_logic;
signal \N__46081\ : std_logic;
signal \N__46078\ : std_logic;
signal \N__46075\ : std_logic;
signal \N__46072\ : std_logic;
signal \N__46067\ : std_logic;
signal \N__46064\ : std_logic;
signal \N__46061\ : std_logic;
signal \N__46060\ : std_logic;
signal \N__46057\ : std_logic;
signal \N__46054\ : std_logic;
signal \N__46051\ : std_logic;
signal \N__46048\ : std_logic;
signal \N__46043\ : std_logic;
signal \N__46040\ : std_logic;
signal \N__46037\ : std_logic;
signal \N__46034\ : std_logic;
signal \N__46031\ : std_logic;
signal \N__46030\ : std_logic;
signal \N__46029\ : std_logic;
signal \N__46028\ : std_logic;
signal \N__46025\ : std_logic;
signal \N__46022\ : std_logic;
signal \N__46021\ : std_logic;
signal \N__46018\ : std_logic;
signal \N__46015\ : std_logic;
signal \N__46012\ : std_logic;
signal \N__46009\ : std_logic;
signal \N__46006\ : std_logic;
signal \N__46003\ : std_logic;
signal \N__46000\ : std_logic;
signal \N__45993\ : std_logic;
signal \N__45986\ : std_logic;
signal \N__45983\ : std_logic;
signal \N__45980\ : std_logic;
signal \N__45977\ : std_logic;
signal \N__45974\ : std_logic;
signal \N__45971\ : std_logic;
signal \N__45968\ : std_logic;
signal \N__45965\ : std_logic;
signal \N__45964\ : std_logic;
signal \N__45961\ : std_logic;
signal \N__45958\ : std_logic;
signal \N__45953\ : std_logic;
signal \N__45950\ : std_logic;
signal \N__45949\ : std_logic;
signal \N__45946\ : std_logic;
signal \N__45943\ : std_logic;
signal \N__45940\ : std_logic;
signal \N__45937\ : std_logic;
signal \N__45934\ : std_logic;
signal \N__45931\ : std_logic;
signal \N__45926\ : std_logic;
signal \N__45925\ : std_logic;
signal \N__45922\ : std_logic;
signal \N__45919\ : std_logic;
signal \N__45916\ : std_logic;
signal \N__45913\ : std_logic;
signal \N__45912\ : std_logic;
signal \N__45909\ : std_logic;
signal \N__45906\ : std_logic;
signal \N__45903\ : std_logic;
signal \N__45896\ : std_logic;
signal \N__45893\ : std_logic;
signal \N__45890\ : std_logic;
signal \N__45889\ : std_logic;
signal \N__45886\ : std_logic;
signal \N__45883\ : std_logic;
signal \N__45878\ : std_logic;
signal \N__45875\ : std_logic;
signal \N__45872\ : std_logic;
signal \N__45869\ : std_logic;
signal \N__45866\ : std_logic;
signal \N__45863\ : std_logic;
signal \N__45860\ : std_logic;
signal \N__45859\ : std_logic;
signal \N__45856\ : std_logic;
signal \N__45853\ : std_logic;
signal \N__45850\ : std_logic;
signal \N__45845\ : std_logic;
signal \N__45842\ : std_logic;
signal \N__45839\ : std_logic;
signal \N__45836\ : std_logic;
signal \N__45833\ : std_logic;
signal \N__45832\ : std_logic;
signal \N__45829\ : std_logic;
signal \N__45826\ : std_logic;
signal \N__45823\ : std_logic;
signal \N__45818\ : std_logic;
signal \N__45815\ : std_logic;
signal \N__45812\ : std_logic;
signal \N__45809\ : std_logic;
signal \N__45806\ : std_logic;
signal \N__45805\ : std_logic;
signal \N__45802\ : std_logic;
signal \N__45799\ : std_logic;
signal \N__45796\ : std_logic;
signal \N__45791\ : std_logic;
signal \N__45788\ : std_logic;
signal \N__45785\ : std_logic;
signal \N__45782\ : std_logic;
signal \N__45779\ : std_logic;
signal \N__45778\ : std_logic;
signal \N__45775\ : std_logic;
signal \N__45772\ : std_logic;
signal \N__45769\ : std_logic;
signal \N__45764\ : std_logic;
signal \N__45761\ : std_logic;
signal \N__45758\ : std_logic;
signal \N__45755\ : std_logic;
signal \N__45752\ : std_logic;
signal \N__45751\ : std_logic;
signal \N__45748\ : std_logic;
signal \N__45745\ : std_logic;
signal \N__45742\ : std_logic;
signal \N__45737\ : std_logic;
signal \N__45734\ : std_logic;
signal \N__45731\ : std_logic;
signal \N__45728\ : std_logic;
signal \N__45725\ : std_logic;
signal \N__45724\ : std_logic;
signal \N__45721\ : std_logic;
signal \N__45718\ : std_logic;
signal \N__45713\ : std_logic;
signal \N__45712\ : std_logic;
signal \N__45709\ : std_logic;
signal \N__45708\ : std_logic;
signal \N__45705\ : std_logic;
signal \N__45702\ : std_logic;
signal \N__45699\ : std_logic;
signal \N__45696\ : std_logic;
signal \N__45695\ : std_logic;
signal \N__45694\ : std_logic;
signal \N__45693\ : std_logic;
signal \N__45686\ : std_logic;
signal \N__45683\ : std_logic;
signal \N__45680\ : std_logic;
signal \N__45677\ : std_logic;
signal \N__45668\ : std_logic;
signal \N__45665\ : std_logic;
signal \N__45662\ : std_logic;
signal \N__45659\ : std_logic;
signal \N__45656\ : std_logic;
signal \N__45653\ : std_logic;
signal \N__45650\ : std_logic;
signal \N__45647\ : std_logic;
signal \N__45644\ : std_logic;
signal \N__45643\ : std_logic;
signal \N__45640\ : std_logic;
signal \N__45637\ : std_logic;
signal \N__45632\ : std_logic;
signal \N__45629\ : std_logic;
signal \N__45626\ : std_logic;
signal \N__45623\ : std_logic;
signal \N__45620\ : std_logic;
signal \N__45617\ : std_logic;
signal \N__45614\ : std_logic;
signal \N__45611\ : std_logic;
signal \N__45610\ : std_logic;
signal \N__45607\ : std_logic;
signal \N__45604\ : std_logic;
signal \N__45599\ : std_logic;
signal \N__45596\ : std_logic;
signal \N__45593\ : std_logic;
signal \N__45590\ : std_logic;
signal \N__45587\ : std_logic;
signal \N__45584\ : std_logic;
signal \N__45581\ : std_logic;
signal \N__45578\ : std_logic;
signal \N__45577\ : std_logic;
signal \N__45574\ : std_logic;
signal \N__45571\ : std_logic;
signal \N__45568\ : std_logic;
signal \N__45563\ : std_logic;
signal \N__45560\ : std_logic;
signal \N__45557\ : std_logic;
signal \N__45554\ : std_logic;
signal \N__45551\ : std_logic;
signal \N__45548\ : std_logic;
signal \N__45547\ : std_logic;
signal \N__45544\ : std_logic;
signal \N__45541\ : std_logic;
signal \N__45536\ : std_logic;
signal \N__45533\ : std_logic;
signal \N__45530\ : std_logic;
signal \N__45527\ : std_logic;
signal \N__45524\ : std_logic;
signal \N__45521\ : std_logic;
signal \N__45518\ : std_logic;
signal \N__45515\ : std_logic;
signal \N__45514\ : std_logic;
signal \N__45511\ : std_logic;
signal \N__45508\ : std_logic;
signal \N__45505\ : std_logic;
signal \N__45500\ : std_logic;
signal \N__45497\ : std_logic;
signal \N__45494\ : std_logic;
signal \N__45491\ : std_logic;
signal \N__45488\ : std_logic;
signal \N__45487\ : std_logic;
signal \N__45484\ : std_logic;
signal \N__45481\ : std_logic;
signal \N__45478\ : std_logic;
signal \N__45473\ : std_logic;
signal \N__45470\ : std_logic;
signal \N__45467\ : std_logic;
signal \N__45464\ : std_logic;
signal \N__45461\ : std_logic;
signal \N__45460\ : std_logic;
signal \N__45457\ : std_logic;
signal \N__45454\ : std_logic;
signal \N__45451\ : std_logic;
signal \N__45446\ : std_logic;
signal \N__45443\ : std_logic;
signal \N__45440\ : std_logic;
signal \N__45437\ : std_logic;
signal \N__45436\ : std_logic;
signal \N__45435\ : std_logic;
signal \N__45430\ : std_logic;
signal \N__45427\ : std_logic;
signal \N__45424\ : std_logic;
signal \N__45419\ : std_logic;
signal \N__45416\ : std_logic;
signal \N__45415\ : std_logic;
signal \N__45412\ : std_logic;
signal \N__45409\ : std_logic;
signal \N__45406\ : std_logic;
signal \N__45401\ : std_logic;
signal \N__45398\ : std_logic;
signal \N__45395\ : std_logic;
signal \N__45392\ : std_logic;
signal \N__45389\ : std_logic;
signal \N__45388\ : std_logic;
signal \N__45387\ : std_logic;
signal \N__45384\ : std_logic;
signal \N__45381\ : std_logic;
signal \N__45378\ : std_logic;
signal \N__45377\ : std_logic;
signal \N__45374\ : std_logic;
signal \N__45373\ : std_logic;
signal \N__45370\ : std_logic;
signal \N__45367\ : std_logic;
signal \N__45364\ : std_logic;
signal \N__45361\ : std_logic;
signal \N__45358\ : std_logic;
signal \N__45347\ : std_logic;
signal \N__45344\ : std_logic;
signal \N__45341\ : std_logic;
signal \N__45338\ : std_logic;
signal \N__45335\ : std_logic;
signal \N__45332\ : std_logic;
signal \N__45329\ : std_logic;
signal \N__45328\ : std_logic;
signal \N__45327\ : std_logic;
signal \N__45324\ : std_logic;
signal \N__45321\ : std_logic;
signal \N__45318\ : std_logic;
signal \N__45315\ : std_logic;
signal \N__45310\ : std_logic;
signal \N__45305\ : std_logic;
signal \N__45302\ : std_logic;
signal \N__45299\ : std_logic;
signal \N__45296\ : std_logic;
signal \N__45295\ : std_logic;
signal \N__45292\ : std_logic;
signal \N__45289\ : std_logic;
signal \N__45284\ : std_logic;
signal \N__45281\ : std_logic;
signal \N__45278\ : std_logic;
signal \N__45275\ : std_logic;
signal \N__45272\ : std_logic;
signal \N__45269\ : std_logic;
signal \N__45266\ : std_logic;
signal \N__45263\ : std_logic;
signal \N__45260\ : std_logic;
signal \N__45257\ : std_logic;
signal \N__45254\ : std_logic;
signal \N__45253\ : std_logic;
signal \N__45250\ : std_logic;
signal \N__45247\ : std_logic;
signal \N__45242\ : std_logic;
signal \N__45239\ : std_logic;
signal \N__45236\ : std_logic;
signal \N__45233\ : std_logic;
signal \N__45230\ : std_logic;
signal \N__45227\ : std_logic;
signal \N__45224\ : std_logic;
signal \N__45221\ : std_logic;
signal \N__45220\ : std_logic;
signal \N__45217\ : std_logic;
signal \N__45214\ : std_logic;
signal \N__45209\ : std_logic;
signal \N__45206\ : std_logic;
signal \N__45203\ : std_logic;
signal \N__45200\ : std_logic;
signal \N__45197\ : std_logic;
signal \N__45194\ : std_logic;
signal \N__45191\ : std_logic;
signal \N__45188\ : std_logic;
signal \N__45187\ : std_logic;
signal \N__45184\ : std_logic;
signal \N__45181\ : std_logic;
signal \N__45176\ : std_logic;
signal \N__45173\ : std_logic;
signal \N__45170\ : std_logic;
signal \N__45167\ : std_logic;
signal \N__45164\ : std_logic;
signal \N__45161\ : std_logic;
signal \N__45158\ : std_logic;
signal \N__45155\ : std_logic;
signal \N__45152\ : std_logic;
signal \N__45151\ : std_logic;
signal \N__45148\ : std_logic;
signal \N__45145\ : std_logic;
signal \N__45140\ : std_logic;
signal \N__45139\ : std_logic;
signal \N__45136\ : std_logic;
signal \N__45133\ : std_logic;
signal \N__45132\ : std_logic;
signal \N__45127\ : std_logic;
signal \N__45124\ : std_logic;
signal \N__45121\ : std_logic;
signal \N__45116\ : std_logic;
signal \N__45113\ : std_logic;
signal \N__45110\ : std_logic;
signal \N__45107\ : std_logic;
signal \N__45106\ : std_logic;
signal \N__45101\ : std_logic;
signal \N__45100\ : std_logic;
signal \N__45097\ : std_logic;
signal \N__45094\ : std_logic;
signal \N__45091\ : std_logic;
signal \N__45086\ : std_logic;
signal \N__45083\ : std_logic;
signal \N__45080\ : std_logic;
signal \N__45077\ : std_logic;
signal \N__45074\ : std_logic;
signal \N__45073\ : std_logic;
signal \N__45070\ : std_logic;
signal \N__45067\ : std_logic;
signal \N__45066\ : std_logic;
signal \N__45061\ : std_logic;
signal \N__45058\ : std_logic;
signal \N__45055\ : std_logic;
signal \N__45050\ : std_logic;
signal \N__45047\ : std_logic;
signal \N__45044\ : std_logic;
signal \N__45041\ : std_logic;
signal \N__45038\ : std_logic;
signal \N__45037\ : std_logic;
signal \N__45034\ : std_logic;
signal \N__45031\ : std_logic;
signal \N__45028\ : std_logic;
signal \N__45027\ : std_logic;
signal \N__45022\ : std_logic;
signal \N__45019\ : std_logic;
signal \N__45016\ : std_logic;
signal \N__45011\ : std_logic;
signal \N__45008\ : std_logic;
signal \N__45005\ : std_logic;
signal \N__45002\ : std_logic;
signal \N__45001\ : std_logic;
signal \N__45000\ : std_logic;
signal \N__44995\ : std_logic;
signal \N__44992\ : std_logic;
signal \N__44989\ : std_logic;
signal \N__44984\ : std_logic;
signal \N__44981\ : std_logic;
signal \N__44978\ : std_logic;
signal \N__44975\ : std_logic;
signal \N__44972\ : std_logic;
signal \N__44971\ : std_logic;
signal \N__44968\ : std_logic;
signal \N__44967\ : std_logic;
signal \N__44964\ : std_logic;
signal \N__44961\ : std_logic;
signal \N__44958\ : std_logic;
signal \N__44955\ : std_logic;
signal \N__44948\ : std_logic;
signal \N__44945\ : std_logic;
signal \N__44942\ : std_logic;
signal \N__44939\ : std_logic;
signal \N__44936\ : std_logic;
signal \N__44933\ : std_logic;
signal \N__44932\ : std_logic;
signal \N__44931\ : std_logic;
signal \N__44928\ : std_logic;
signal \N__44925\ : std_logic;
signal \N__44922\ : std_logic;
signal \N__44919\ : std_logic;
signal \N__44916\ : std_logic;
signal \N__44909\ : std_logic;
signal \N__44906\ : std_logic;
signal \N__44903\ : std_logic;
signal \N__44900\ : std_logic;
signal \N__44897\ : std_logic;
signal \N__44894\ : std_logic;
signal \N__44893\ : std_logic;
signal \N__44890\ : std_logic;
signal \N__44887\ : std_logic;
signal \N__44884\ : std_logic;
signal \N__44879\ : std_logic;
signal \N__44878\ : std_logic;
signal \N__44875\ : std_logic;
signal \N__44872\ : std_logic;
signal \N__44871\ : std_logic;
signal \N__44866\ : std_logic;
signal \N__44863\ : std_logic;
signal \N__44860\ : std_logic;
signal \N__44855\ : std_logic;
signal \N__44852\ : std_logic;
signal \N__44849\ : std_logic;
signal \N__44846\ : std_logic;
signal \N__44845\ : std_logic;
signal \N__44842\ : std_logic;
signal \N__44839\ : std_logic;
signal \N__44836\ : std_logic;
signal \N__44835\ : std_logic;
signal \N__44830\ : std_logic;
signal \N__44827\ : std_logic;
signal \N__44824\ : std_logic;
signal \N__44819\ : std_logic;
signal \N__44816\ : std_logic;
signal \N__44815\ : std_logic;
signal \N__44812\ : std_logic;
signal \N__44809\ : std_logic;
signal \N__44808\ : std_logic;
signal \N__44803\ : std_logic;
signal \N__44800\ : std_logic;
signal \N__44797\ : std_logic;
signal \N__44792\ : std_logic;
signal \N__44789\ : std_logic;
signal \N__44788\ : std_logic;
signal \N__44785\ : std_logic;
signal \N__44782\ : std_logic;
signal \N__44781\ : std_logic;
signal \N__44776\ : std_logic;
signal \N__44773\ : std_logic;
signal \N__44770\ : std_logic;
signal \N__44765\ : std_logic;
signal \N__44762\ : std_logic;
signal \N__44761\ : std_logic;
signal \N__44760\ : std_logic;
signal \N__44755\ : std_logic;
signal \N__44752\ : std_logic;
signal \N__44749\ : std_logic;
signal \N__44744\ : std_logic;
signal \N__44741\ : std_logic;
signal \N__44740\ : std_logic;
signal \N__44739\ : std_logic;
signal \N__44734\ : std_logic;
signal \N__44731\ : std_logic;
signal \N__44728\ : std_logic;
signal \N__44723\ : std_logic;
signal \N__44720\ : std_logic;
signal \N__44719\ : std_logic;
signal \N__44716\ : std_logic;
signal \N__44715\ : std_logic;
signal \N__44712\ : std_logic;
signal \N__44709\ : std_logic;
signal \N__44706\ : std_logic;
signal \N__44701\ : std_logic;
signal \N__44696\ : std_logic;
signal \N__44693\ : std_logic;
signal \N__44692\ : std_logic;
signal \N__44689\ : std_logic;
signal \N__44688\ : std_logic;
signal \N__44685\ : std_logic;
signal \N__44682\ : std_logic;
signal \N__44679\ : std_logic;
signal \N__44676\ : std_logic;
signal \N__44669\ : std_logic;
signal \N__44666\ : std_logic;
signal \N__44663\ : std_logic;
signal \N__44660\ : std_logic;
signal \N__44659\ : std_logic;
signal \N__44656\ : std_logic;
signal \N__44653\ : std_logic;
signal \N__44652\ : std_logic;
signal \N__44647\ : std_logic;
signal \N__44644\ : std_logic;
signal \N__44641\ : std_logic;
signal \N__44636\ : std_logic;
signal \N__44633\ : std_logic;
signal \N__44630\ : std_logic;
signal \N__44627\ : std_logic;
signal \N__44626\ : std_logic;
signal \N__44623\ : std_logic;
signal \N__44620\ : std_logic;
signal \N__44619\ : std_logic;
signal \N__44614\ : std_logic;
signal \N__44611\ : std_logic;
signal \N__44608\ : std_logic;
signal \N__44603\ : std_logic;
signal \N__44600\ : std_logic;
signal \N__44599\ : std_logic;
signal \N__44596\ : std_logic;
signal \N__44593\ : std_logic;
signal \N__44592\ : std_logic;
signal \N__44587\ : std_logic;
signal \N__44584\ : std_logic;
signal \N__44581\ : std_logic;
signal \N__44576\ : std_logic;
signal \N__44573\ : std_logic;
signal \N__44572\ : std_logic;
signal \N__44567\ : std_logic;
signal \N__44566\ : std_logic;
signal \N__44563\ : std_logic;
signal \N__44560\ : std_logic;
signal \N__44557\ : std_logic;
signal \N__44552\ : std_logic;
signal \N__44549\ : std_logic;
signal \N__44548\ : std_logic;
signal \N__44543\ : std_logic;
signal \N__44542\ : std_logic;
signal \N__44539\ : std_logic;
signal \N__44536\ : std_logic;
signal \N__44533\ : std_logic;
signal \N__44528\ : std_logic;
signal \N__44525\ : std_logic;
signal \N__44524\ : std_logic;
signal \N__44521\ : std_logic;
signal \N__44518\ : std_logic;
signal \N__44515\ : std_logic;
signal \N__44514\ : std_logic;
signal \N__44509\ : std_logic;
signal \N__44506\ : std_logic;
signal \N__44503\ : std_logic;
signal \N__44498\ : std_logic;
signal \N__44495\ : std_logic;
signal \N__44494\ : std_logic;
signal \N__44491\ : std_logic;
signal \N__44488\ : std_logic;
signal \N__44483\ : std_logic;
signal \N__44482\ : std_logic;
signal \N__44479\ : std_logic;
signal \N__44476\ : std_logic;
signal \N__44473\ : std_logic;
signal \N__44468\ : std_logic;
signal \N__44465\ : std_logic;
signal \N__44462\ : std_logic;
signal \N__44461\ : std_logic;
signal \N__44458\ : std_logic;
signal \N__44457\ : std_logic;
signal \N__44454\ : std_logic;
signal \N__44451\ : std_logic;
signal \N__44448\ : std_logic;
signal \N__44445\ : std_logic;
signal \N__44438\ : std_logic;
signal \N__44435\ : std_logic;
signal \N__44432\ : std_logic;
signal \N__44431\ : std_logic;
signal \N__44430\ : std_logic;
signal \N__44427\ : std_logic;
signal \N__44424\ : std_logic;
signal \N__44421\ : std_logic;
signal \N__44414\ : std_logic;
signal \N__44411\ : std_logic;
signal \N__44410\ : std_logic;
signal \N__44407\ : std_logic;
signal \N__44404\ : std_logic;
signal \N__44401\ : std_logic;
signal \N__44400\ : std_logic;
signal \N__44395\ : std_logic;
signal \N__44392\ : std_logic;
signal \N__44389\ : std_logic;
signal \N__44384\ : std_logic;
signal \N__44381\ : std_logic;
signal \N__44378\ : std_logic;
signal \N__44375\ : std_logic;
signal \N__44374\ : std_logic;
signal \N__44373\ : std_logic;
signal \N__44370\ : std_logic;
signal \N__44367\ : std_logic;
signal \N__44364\ : std_logic;
signal \N__44357\ : std_logic;
signal \N__44356\ : std_logic;
signal \N__44355\ : std_logic;
signal \N__44352\ : std_logic;
signal \N__44349\ : std_logic;
signal \N__44346\ : std_logic;
signal \N__44341\ : std_logic;
signal \N__44336\ : std_logic;
signal \N__44333\ : std_logic;
signal \N__44332\ : std_logic;
signal \N__44331\ : std_logic;
signal \N__44330\ : std_logic;
signal \N__44329\ : std_logic;
signal \N__44328\ : std_logic;
signal \N__44315\ : std_logic;
signal \N__44312\ : std_logic;
signal \N__44309\ : std_logic;
signal \N__44306\ : std_logic;
signal \N__44305\ : std_logic;
signal \N__44302\ : std_logic;
signal \N__44299\ : std_logic;
signal \N__44298\ : std_logic;
signal \N__44293\ : std_logic;
signal \N__44290\ : std_logic;
signal \N__44285\ : std_logic;
signal \N__44284\ : std_logic;
signal \N__44281\ : std_logic;
signal \N__44278\ : std_logic;
signal \N__44277\ : std_logic;
signal \N__44274\ : std_logic;
signal \N__44271\ : std_logic;
signal \N__44268\ : std_logic;
signal \N__44261\ : std_logic;
signal \N__44258\ : std_logic;
signal \N__44257\ : std_logic;
signal \N__44254\ : std_logic;
signal \N__44251\ : std_logic;
signal \N__44250\ : std_logic;
signal \N__44247\ : std_logic;
signal \N__44244\ : std_logic;
signal \N__44241\ : std_logic;
signal \N__44236\ : std_logic;
signal \N__44233\ : std_logic;
signal \N__44228\ : std_logic;
signal \N__44227\ : std_logic;
signal \N__44224\ : std_logic;
signal \N__44221\ : std_logic;
signal \N__44220\ : std_logic;
signal \N__44217\ : std_logic;
signal \N__44214\ : std_logic;
signal \N__44211\ : std_logic;
signal \N__44204\ : std_logic;
signal \N__44201\ : std_logic;
signal \N__44200\ : std_logic;
signal \N__44197\ : std_logic;
signal \N__44194\ : std_logic;
signal \N__44189\ : std_logic;
signal \N__44186\ : std_logic;
signal \N__44185\ : std_logic;
signal \N__44184\ : std_logic;
signal \N__44183\ : std_logic;
signal \N__44182\ : std_logic;
signal \N__44181\ : std_logic;
signal \N__44178\ : std_logic;
signal \N__44175\ : std_logic;
signal \N__44168\ : std_logic;
signal \N__44165\ : std_logic;
signal \N__44156\ : std_logic;
signal \N__44153\ : std_logic;
signal \N__44150\ : std_logic;
signal \N__44149\ : std_logic;
signal \N__44146\ : std_logic;
signal \N__44145\ : std_logic;
signal \N__44142\ : std_logic;
signal \N__44139\ : std_logic;
signal \N__44138\ : std_logic;
signal \N__44135\ : std_logic;
signal \N__44134\ : std_logic;
signal \N__44133\ : std_logic;
signal \N__44130\ : std_logic;
signal \N__44127\ : std_logic;
signal \N__44124\ : std_logic;
signal \N__44121\ : std_logic;
signal \N__44118\ : std_logic;
signal \N__44115\ : std_logic;
signal \N__44112\ : std_logic;
signal \N__44107\ : std_logic;
signal \N__44102\ : std_logic;
signal \N__44099\ : std_logic;
signal \N__44090\ : std_logic;
signal \N__44087\ : std_logic;
signal \N__44084\ : std_logic;
signal \N__44081\ : std_logic;
signal \N__44080\ : std_logic;
signal \N__44079\ : std_logic;
signal \N__44078\ : std_logic;
signal \N__44075\ : std_logic;
signal \N__44072\ : std_logic;
signal \N__44071\ : std_logic;
signal \N__44068\ : std_logic;
signal \N__44067\ : std_logic;
signal \N__44064\ : std_logic;
signal \N__44061\ : std_logic;
signal \N__44058\ : std_logic;
signal \N__44055\ : std_logic;
signal \N__44052\ : std_logic;
signal \N__44049\ : std_logic;
signal \N__44046\ : std_logic;
signal \N__44043\ : std_logic;
signal \N__44040\ : std_logic;
signal \N__44037\ : std_logic;
signal \N__44032\ : std_logic;
signal \N__44021\ : std_logic;
signal \N__44020\ : std_logic;
signal \N__44017\ : std_logic;
signal \N__44016\ : std_logic;
signal \N__44015\ : std_logic;
signal \N__44014\ : std_logic;
signal \N__44013\ : std_logic;
signal \N__44010\ : std_logic;
signal \N__44007\ : std_logic;
signal \N__44000\ : std_logic;
signal \N__43997\ : std_logic;
signal \N__43994\ : std_logic;
signal \N__43991\ : std_logic;
signal \N__43988\ : std_logic;
signal \N__43985\ : std_logic;
signal \N__43982\ : std_logic;
signal \N__43977\ : std_logic;
signal \N__43970\ : std_logic;
signal \N__43967\ : std_logic;
signal \N__43964\ : std_logic;
signal \N__43963\ : std_logic;
signal \N__43960\ : std_logic;
signal \N__43957\ : std_logic;
signal \N__43956\ : std_logic;
signal \N__43951\ : std_logic;
signal \N__43950\ : std_logic;
signal \N__43947\ : std_logic;
signal \N__43944\ : std_logic;
signal \N__43943\ : std_logic;
signal \N__43940\ : std_logic;
signal \N__43935\ : std_logic;
signal \N__43932\ : std_logic;
signal \N__43929\ : std_logic;
signal \N__43928\ : std_logic;
signal \N__43925\ : std_logic;
signal \N__43922\ : std_logic;
signal \N__43919\ : std_logic;
signal \N__43916\ : std_logic;
signal \N__43907\ : std_logic;
signal \N__43904\ : std_logic;
signal \N__43901\ : std_logic;
signal \N__43900\ : std_logic;
signal \N__43897\ : std_logic;
signal \N__43896\ : std_logic;
signal \N__43893\ : std_logic;
signal \N__43890\ : std_logic;
signal \N__43887\ : std_logic;
signal \N__43880\ : std_logic;
signal \N__43879\ : std_logic;
signal \N__43876\ : std_logic;
signal \N__43875\ : std_logic;
signal \N__43872\ : std_logic;
signal \N__43869\ : std_logic;
signal \N__43866\ : std_logic;
signal \N__43859\ : std_logic;
signal \N__43856\ : std_logic;
signal \N__43855\ : std_logic;
signal \N__43854\ : std_logic;
signal \N__43853\ : std_logic;
signal \N__43852\ : std_logic;
signal \N__43849\ : std_logic;
signal \N__43846\ : std_logic;
signal \N__43845\ : std_logic;
signal \N__43844\ : std_logic;
signal \N__43843\ : std_logic;
signal \N__43842\ : std_logic;
signal \N__43841\ : std_logic;
signal \N__43840\ : std_logic;
signal \N__43839\ : std_logic;
signal \N__43836\ : std_logic;
signal \N__43835\ : std_logic;
signal \N__43834\ : std_logic;
signal \N__43833\ : std_logic;
signal \N__43830\ : std_logic;
signal \N__43829\ : std_logic;
signal \N__43828\ : std_logic;
signal \N__43827\ : std_logic;
signal \N__43826\ : std_logic;
signal \N__43825\ : std_logic;
signal \N__43824\ : std_logic;
signal \N__43823\ : std_logic;
signal \N__43822\ : std_logic;
signal \N__43819\ : std_logic;
signal \N__43816\ : std_logic;
signal \N__43799\ : std_logic;
signal \N__43796\ : std_logic;
signal \N__43791\ : std_logic;
signal \N__43790\ : std_logic;
signal \N__43787\ : std_logic;
signal \N__43784\ : std_logic;
signal \N__43767\ : std_logic;
signal \N__43764\ : std_logic;
signal \N__43755\ : std_logic;
signal \N__43750\ : std_logic;
signal \N__43747\ : std_logic;
signal \N__43740\ : std_logic;
signal \N__43733\ : std_logic;
signal \N__43732\ : std_logic;
signal \N__43729\ : std_logic;
signal \N__43728\ : std_logic;
signal \N__43725\ : std_logic;
signal \N__43724\ : std_logic;
signal \N__43723\ : std_logic;
signal \N__43722\ : std_logic;
signal \N__43721\ : std_logic;
signal \N__43720\ : std_logic;
signal \N__43715\ : std_logic;
signal \N__43714\ : std_logic;
signal \N__43713\ : std_logic;
signal \N__43712\ : std_logic;
signal \N__43711\ : std_logic;
signal \N__43710\ : std_logic;
signal \N__43707\ : std_logic;
signal \N__43704\ : std_logic;
signal \N__43703\ : std_logic;
signal \N__43702\ : std_logic;
signal \N__43701\ : std_logic;
signal \N__43700\ : std_logic;
signal \N__43697\ : std_logic;
signal \N__43694\ : std_logic;
signal \N__43691\ : std_logic;
signal \N__43688\ : std_logic;
signal \N__43685\ : std_logic;
signal \N__43682\ : std_logic;
signal \N__43681\ : std_logic;
signal \N__43678\ : std_logic;
signal \N__43675\ : std_logic;
signal \N__43672\ : std_logic;
signal \N__43669\ : std_logic;
signal \N__43668\ : std_logic;
signal \N__43667\ : std_logic;
signal \N__43666\ : std_logic;
signal \N__43665\ : std_logic;
signal \N__43664\ : std_logic;
signal \N__43661\ : std_logic;
signal \N__43660\ : std_logic;
signal \N__43657\ : std_logic;
signal \N__43640\ : std_logic;
signal \N__43635\ : std_logic;
signal \N__43618\ : std_logic;
signal \N__43613\ : std_logic;
signal \N__43610\ : std_logic;
signal \N__43607\ : std_logic;
signal \N__43600\ : std_logic;
signal \N__43589\ : std_logic;
signal \N__43588\ : std_logic;
signal \N__43587\ : std_logic;
signal \N__43586\ : std_logic;
signal \N__43585\ : std_logic;
signal \N__43584\ : std_logic;
signal \N__43583\ : std_logic;
signal \N__43580\ : std_logic;
signal \N__43577\ : std_logic;
signal \N__43574\ : std_logic;
signal \N__43573\ : std_logic;
signal \N__43572\ : std_logic;
signal \N__43571\ : std_logic;
signal \N__43570\ : std_logic;
signal \N__43569\ : std_logic;
signal \N__43568\ : std_logic;
signal \N__43565\ : std_logic;
signal \N__43564\ : std_logic;
signal \N__43561\ : std_logic;
signal \N__43560\ : std_logic;
signal \N__43559\ : std_logic;
signal \N__43558\ : std_logic;
signal \N__43557\ : std_logic;
signal \N__43556\ : std_logic;
signal \N__43555\ : std_logic;
signal \N__43554\ : std_logic;
signal \N__43553\ : std_logic;
signal \N__43550\ : std_logic;
signal \N__43547\ : std_logic;
signal \N__43540\ : std_logic;
signal \N__43529\ : std_logic;
signal \N__43526\ : std_logic;
signal \N__43521\ : std_logic;
signal \N__43520\ : std_logic;
signal \N__43519\ : std_logic;
signal \N__43516\ : std_logic;
signal \N__43499\ : std_logic;
signal \N__43494\ : std_logic;
signal \N__43485\ : std_logic;
signal \N__43480\ : std_logic;
signal \N__43477\ : std_logic;
signal \N__43470\ : std_logic;
signal \N__43463\ : std_logic;
signal \N__43460\ : std_logic;
signal \N__43457\ : std_logic;
signal \N__43456\ : std_logic;
signal \N__43453\ : std_logic;
signal \N__43450\ : std_logic;
signal \N__43445\ : std_logic;
signal \N__43442\ : std_logic;
signal \N__43441\ : std_logic;
signal \N__43440\ : std_logic;
signal \N__43439\ : std_logic;
signal \N__43438\ : std_logic;
signal \N__43437\ : std_logic;
signal \N__43436\ : std_logic;
signal \N__43435\ : std_logic;
signal \N__43434\ : std_logic;
signal \N__43431\ : std_logic;
signal \N__43424\ : std_logic;
signal \N__43413\ : std_logic;
signal \N__43412\ : std_logic;
signal \N__43411\ : std_logic;
signal \N__43410\ : std_logic;
signal \N__43409\ : std_logic;
signal \N__43408\ : std_logic;
signal \N__43407\ : std_logic;
signal \N__43406\ : std_logic;
signal \N__43403\ : std_logic;
signal \N__43400\ : std_logic;
signal \N__43397\ : std_logic;
signal \N__43382\ : std_logic;
signal \N__43373\ : std_logic;
signal \N__43370\ : std_logic;
signal \N__43367\ : std_logic;
signal \N__43364\ : std_logic;
signal \N__43361\ : std_logic;
signal \N__43358\ : std_logic;
signal \N__43355\ : std_logic;
signal \N__43354\ : std_logic;
signal \N__43353\ : std_logic;
signal \N__43352\ : std_logic;
signal \N__43349\ : std_logic;
signal \N__43348\ : std_logic;
signal \N__43345\ : std_logic;
signal \N__43342\ : std_logic;
signal \N__43339\ : std_logic;
signal \N__43336\ : std_logic;
signal \N__43333\ : std_logic;
signal \N__43330\ : std_logic;
signal \N__43325\ : std_logic;
signal \N__43318\ : std_logic;
signal \N__43315\ : std_logic;
signal \N__43310\ : std_logic;
signal \N__43309\ : std_logic;
signal \N__43304\ : std_logic;
signal \N__43303\ : std_logic;
signal \N__43302\ : std_logic;
signal \N__43301\ : std_logic;
signal \N__43300\ : std_logic;
signal \N__43299\ : std_logic;
signal \N__43298\ : std_logic;
signal \N__43297\ : std_logic;
signal \N__43296\ : std_logic;
signal \N__43293\ : std_logic;
signal \N__43290\ : std_logic;
signal \N__43281\ : std_logic;
signal \N__43274\ : std_logic;
signal \N__43265\ : std_logic;
signal \N__43264\ : std_logic;
signal \N__43263\ : std_logic;
signal \N__43260\ : std_logic;
signal \N__43257\ : std_logic;
signal \N__43254\ : std_logic;
signal \N__43249\ : std_logic;
signal \N__43244\ : std_logic;
signal \N__43243\ : std_logic;
signal \N__43238\ : std_logic;
signal \N__43237\ : std_logic;
signal \N__43236\ : std_logic;
signal \N__43233\ : std_logic;
signal \N__43228\ : std_logic;
signal \N__43223\ : std_logic;
signal \N__43222\ : std_logic;
signal \N__43219\ : std_logic;
signal \N__43218\ : std_logic;
signal \N__43215\ : std_logic;
signal \N__43212\ : std_logic;
signal \N__43209\ : std_logic;
signal \N__43206\ : std_logic;
signal \N__43203\ : std_logic;
signal \N__43200\ : std_logic;
signal \N__43197\ : std_logic;
signal \N__43190\ : std_logic;
signal \N__43189\ : std_logic;
signal \N__43188\ : std_logic;
signal \N__43187\ : std_logic;
signal \N__43186\ : std_logic;
signal \N__43185\ : std_logic;
signal \N__43176\ : std_logic;
signal \N__43171\ : std_logic;
signal \N__43166\ : std_logic;
signal \N__43165\ : std_logic;
signal \N__43164\ : std_logic;
signal \N__43163\ : std_logic;
signal \N__43162\ : std_logic;
signal \N__43161\ : std_logic;
signal \N__43160\ : std_logic;
signal \N__43157\ : std_logic;
signal \N__43154\ : std_logic;
signal \N__43143\ : std_logic;
signal \N__43136\ : std_logic;
signal \N__43133\ : std_logic;
signal \N__43130\ : std_logic;
signal \N__43127\ : std_logic;
signal \N__43124\ : std_logic;
signal \N__43123\ : std_logic;
signal \N__43120\ : std_logic;
signal \N__43117\ : std_logic;
signal \N__43112\ : std_logic;
signal \N__43111\ : std_logic;
signal \N__43110\ : std_logic;
signal \N__43107\ : std_logic;
signal \N__43104\ : std_logic;
signal \N__43103\ : std_logic;
signal \N__43100\ : std_logic;
signal \N__43095\ : std_logic;
signal \N__43094\ : std_logic;
signal \N__43091\ : std_logic;
signal \N__43088\ : std_logic;
signal \N__43085\ : std_logic;
signal \N__43082\ : std_logic;
signal \N__43079\ : std_logic;
signal \N__43076\ : std_logic;
signal \N__43071\ : std_logic;
signal \N__43064\ : std_logic;
signal \N__43063\ : std_logic;
signal \N__43062\ : std_logic;
signal \N__43061\ : std_logic;
signal \N__43058\ : std_logic;
signal \N__43055\ : std_logic;
signal \N__43050\ : std_logic;
signal \N__43043\ : std_logic;
signal \N__43040\ : std_logic;
signal \N__43037\ : std_logic;
signal \N__43034\ : std_logic;
signal \N__43033\ : std_logic;
signal \N__43032\ : std_logic;
signal \N__43029\ : std_logic;
signal \N__43024\ : std_logic;
signal \N__43023\ : std_logic;
signal \N__43022\ : std_logic;
signal \N__43019\ : std_logic;
signal \N__43016\ : std_logic;
signal \N__43015\ : std_logic;
signal \N__43010\ : std_logic;
signal \N__43007\ : std_logic;
signal \N__43004\ : std_logic;
signal \N__43001\ : std_logic;
signal \N__42998\ : std_logic;
signal \N__42989\ : std_logic;
signal \N__42988\ : std_logic;
signal \N__42985\ : std_logic;
signal \N__42982\ : std_logic;
signal \N__42981\ : std_logic;
signal \N__42980\ : std_logic;
signal \N__42977\ : std_logic;
signal \N__42974\ : std_logic;
signal \N__42971\ : std_logic;
signal \N__42968\ : std_logic;
signal \N__42965\ : std_logic;
signal \N__42956\ : std_logic;
signal \N__42953\ : std_logic;
signal \N__42950\ : std_logic;
signal \N__42947\ : std_logic;
signal \N__42944\ : std_logic;
signal \N__42941\ : std_logic;
signal \N__42938\ : std_logic;
signal \N__42935\ : std_logic;
signal \N__42932\ : std_logic;
signal \N__42929\ : std_logic;
signal \N__42926\ : std_logic;
signal \N__42923\ : std_logic;
signal \N__42920\ : std_logic;
signal \N__42917\ : std_logic;
signal \N__42914\ : std_logic;
signal \N__42911\ : std_logic;
signal \N__42908\ : std_logic;
signal \N__42905\ : std_logic;
signal \N__42904\ : std_logic;
signal \N__42903\ : std_logic;
signal \N__42900\ : std_logic;
signal \N__42897\ : std_logic;
signal \N__42894\ : std_logic;
signal \N__42893\ : std_logic;
signal \N__42892\ : std_logic;
signal \N__42891\ : std_logic;
signal \N__42888\ : std_logic;
signal \N__42885\ : std_logic;
signal \N__42882\ : std_logic;
signal \N__42877\ : std_logic;
signal \N__42874\ : std_logic;
signal \N__42863\ : std_logic;
signal \N__42862\ : std_logic;
signal \N__42861\ : std_logic;
signal \N__42856\ : std_logic;
signal \N__42853\ : std_logic;
signal \N__42850\ : std_logic;
signal \N__42847\ : std_logic;
signal \N__42844\ : std_logic;
signal \N__42841\ : std_logic;
signal \N__42838\ : std_logic;
signal \N__42835\ : std_logic;
signal \N__42832\ : std_logic;
signal \N__42827\ : std_logic;
signal \N__42824\ : std_logic;
signal \N__42823\ : std_logic;
signal \N__42818\ : std_logic;
signal \N__42817\ : std_logic;
signal \N__42814\ : std_logic;
signal \N__42813\ : std_logic;
signal \N__42812\ : std_logic;
signal \N__42809\ : std_logic;
signal \N__42806\ : std_logic;
signal \N__42803\ : std_logic;
signal \N__42800\ : std_logic;
signal \N__42797\ : std_logic;
signal \N__42794\ : std_logic;
signal \N__42785\ : std_logic;
signal \N__42782\ : std_logic;
signal \N__42781\ : std_logic;
signal \N__42778\ : std_logic;
signal \N__42775\ : std_logic;
signal \N__42774\ : std_logic;
signal \N__42771\ : std_logic;
signal \N__42768\ : std_logic;
signal \N__42765\ : std_logic;
signal \N__42762\ : std_logic;
signal \N__42755\ : std_logic;
signal \N__42752\ : std_logic;
signal \N__42749\ : std_logic;
signal \N__42746\ : std_logic;
signal \N__42743\ : std_logic;
signal \N__42740\ : std_logic;
signal \N__42739\ : std_logic;
signal \N__42738\ : std_logic;
signal \N__42737\ : std_logic;
signal \N__42736\ : std_logic;
signal \N__42735\ : std_logic;
signal \N__42734\ : std_logic;
signal \N__42733\ : std_logic;
signal \N__42724\ : std_logic;
signal \N__42723\ : std_logic;
signal \N__42722\ : std_logic;
signal \N__42721\ : std_logic;
signal \N__42720\ : std_logic;
signal \N__42719\ : std_logic;
signal \N__42718\ : std_logic;
signal \N__42717\ : std_logic;
signal \N__42716\ : std_logic;
signal \N__42715\ : std_logic;
signal \N__42714\ : std_logic;
signal \N__42713\ : std_logic;
signal \N__42712\ : std_logic;
signal \N__42711\ : std_logic;
signal \N__42710\ : std_logic;
signal \N__42709\ : std_logic;
signal \N__42708\ : std_logic;
signal \N__42707\ : std_logic;
signal \N__42706\ : std_logic;
signal \N__42705\ : std_logic;
signal \N__42704\ : std_logic;
signal \N__42703\ : std_logic;
signal \N__42702\ : std_logic;
signal \N__42693\ : std_logic;
signal \N__42690\ : std_logic;
signal \N__42681\ : std_logic;
signal \N__42672\ : std_logic;
signal \N__42663\ : std_logic;
signal \N__42654\ : std_logic;
signal \N__42649\ : std_logic;
signal \N__42640\ : std_logic;
signal \N__42633\ : std_logic;
signal \N__42626\ : std_logic;
signal \N__42621\ : std_logic;
signal \N__42616\ : std_logic;
signal \N__42613\ : std_logic;
signal \N__42610\ : std_logic;
signal \N__42607\ : std_logic;
signal \N__42602\ : std_logic;
signal \N__42599\ : std_logic;
signal \N__42596\ : std_logic;
signal \N__42595\ : std_logic;
signal \N__42592\ : std_logic;
signal \N__42591\ : std_logic;
signal \N__42590\ : std_logic;
signal \N__42587\ : std_logic;
signal \N__42584\ : std_logic;
signal \N__42581\ : std_logic;
signal \N__42578\ : std_logic;
signal \N__42575\ : std_logic;
signal \N__42572\ : std_logic;
signal \N__42569\ : std_logic;
signal \N__42566\ : std_logic;
signal \N__42563\ : std_logic;
signal \N__42560\ : std_logic;
signal \N__42557\ : std_logic;
signal \N__42554\ : std_logic;
signal \N__42551\ : std_logic;
signal \N__42548\ : std_logic;
signal \N__42545\ : std_logic;
signal \N__42542\ : std_logic;
signal \N__42533\ : std_logic;
signal \N__42530\ : std_logic;
signal \N__42527\ : std_logic;
signal \N__42524\ : std_logic;
signal \N__42521\ : std_logic;
signal \N__42518\ : std_logic;
signal \N__42515\ : std_logic;
signal \N__42512\ : std_logic;
signal \N__42509\ : std_logic;
signal \N__42506\ : std_logic;
signal \N__42503\ : std_logic;
signal \N__42500\ : std_logic;
signal \N__42497\ : std_logic;
signal \N__42494\ : std_logic;
signal \N__42491\ : std_logic;
signal \N__42488\ : std_logic;
signal \N__42485\ : std_logic;
signal \N__42482\ : std_logic;
signal \N__42479\ : std_logic;
signal \N__42476\ : std_logic;
signal \N__42475\ : std_logic;
signal \N__42474\ : std_logic;
signal \N__42471\ : std_logic;
signal \N__42470\ : std_logic;
signal \N__42467\ : std_logic;
signal \N__42464\ : std_logic;
signal \N__42461\ : std_logic;
signal \N__42458\ : std_logic;
signal \N__42455\ : std_logic;
signal \N__42448\ : std_logic;
signal \N__42445\ : std_logic;
signal \N__42442\ : std_logic;
signal \N__42437\ : std_logic;
signal \N__42436\ : std_logic;
signal \N__42433\ : std_logic;
signal \N__42432\ : std_logic;
signal \N__42431\ : std_logic;
signal \N__42428\ : std_logic;
signal \N__42425\ : std_logic;
signal \N__42422\ : std_logic;
signal \N__42419\ : std_logic;
signal \N__42416\ : std_logic;
signal \N__42409\ : std_logic;
signal \N__42404\ : std_logic;
signal \N__42401\ : std_logic;
signal \N__42398\ : std_logic;
signal \N__42395\ : std_logic;
signal \N__42392\ : std_logic;
signal \N__42391\ : std_logic;
signal \N__42388\ : std_logic;
signal \N__42385\ : std_logic;
signal \N__42380\ : std_logic;
signal \N__42379\ : std_logic;
signal \N__42376\ : std_logic;
signal \N__42373\ : std_logic;
signal \N__42370\ : std_logic;
signal \N__42369\ : std_logic;
signal \N__42366\ : std_logic;
signal \N__42363\ : std_logic;
signal \N__42360\ : std_logic;
signal \N__42357\ : std_logic;
signal \N__42354\ : std_logic;
signal \N__42347\ : std_logic;
signal \N__42344\ : std_logic;
signal \N__42341\ : std_logic;
signal \N__42338\ : std_logic;
signal \N__42335\ : std_logic;
signal \N__42332\ : std_logic;
signal \N__42329\ : std_logic;
signal \N__42326\ : std_logic;
signal \N__42323\ : std_logic;
signal \N__42320\ : std_logic;
signal \N__42319\ : std_logic;
signal \N__42318\ : std_logic;
signal \N__42315\ : std_logic;
signal \N__42312\ : std_logic;
signal \N__42309\ : std_logic;
signal \N__42306\ : std_logic;
signal \N__42299\ : std_logic;
signal \N__42296\ : std_logic;
signal \N__42293\ : std_logic;
signal \N__42290\ : std_logic;
signal \N__42289\ : std_logic;
signal \N__42288\ : std_logic;
signal \N__42285\ : std_logic;
signal \N__42282\ : std_logic;
signal \N__42279\ : std_logic;
signal \N__42276\ : std_logic;
signal \N__42269\ : std_logic;
signal \N__42266\ : std_logic;
signal \N__42263\ : std_logic;
signal \N__42260\ : std_logic;
signal \N__42259\ : std_logic;
signal \N__42258\ : std_logic;
signal \N__42255\ : std_logic;
signal \N__42252\ : std_logic;
signal \N__42249\ : std_logic;
signal \N__42246\ : std_logic;
signal \N__42239\ : std_logic;
signal \N__42236\ : std_logic;
signal \N__42233\ : std_logic;
signal \N__42230\ : std_logic;
signal \N__42229\ : std_logic;
signal \N__42228\ : std_logic;
signal \N__42225\ : std_logic;
signal \N__42222\ : std_logic;
signal \N__42219\ : std_logic;
signal \N__42216\ : std_logic;
signal \N__42209\ : std_logic;
signal \N__42206\ : std_logic;
signal \N__42203\ : std_logic;
signal \N__42200\ : std_logic;
signal \N__42199\ : std_logic;
signal \N__42198\ : std_logic;
signal \N__42195\ : std_logic;
signal \N__42192\ : std_logic;
signal \N__42189\ : std_logic;
signal \N__42186\ : std_logic;
signal \N__42179\ : std_logic;
signal \N__42176\ : std_logic;
signal \N__42173\ : std_logic;
signal \N__42170\ : std_logic;
signal \N__42169\ : std_logic;
signal \N__42168\ : std_logic;
signal \N__42165\ : std_logic;
signal \N__42162\ : std_logic;
signal \N__42159\ : std_logic;
signal \N__42156\ : std_logic;
signal \N__42149\ : std_logic;
signal \N__42146\ : std_logic;
signal \N__42143\ : std_logic;
signal \N__42140\ : std_logic;
signal \N__42139\ : std_logic;
signal \N__42138\ : std_logic;
signal \N__42135\ : std_logic;
signal \N__42132\ : std_logic;
signal \N__42129\ : std_logic;
signal \N__42126\ : std_logic;
signal \N__42119\ : std_logic;
signal \N__42118\ : std_logic;
signal \N__42115\ : std_logic;
signal \N__42112\ : std_logic;
signal \N__42109\ : std_logic;
signal \N__42104\ : std_logic;
signal \N__42101\ : std_logic;
signal \N__42098\ : std_logic;
signal \N__42095\ : std_logic;
signal \N__42094\ : std_logic;
signal \N__42093\ : std_logic;
signal \N__42090\ : std_logic;
signal \N__42087\ : std_logic;
signal \N__42084\ : std_logic;
signal \N__42081\ : std_logic;
signal \N__42074\ : std_logic;
signal \N__42073\ : std_logic;
signal \N__42070\ : std_logic;
signal \N__42067\ : std_logic;
signal \N__42064\ : std_logic;
signal \N__42059\ : std_logic;
signal \N__42056\ : std_logic;
signal \N__42053\ : std_logic;
signal \N__42050\ : std_logic;
signal \N__42047\ : std_logic;
signal \N__42046\ : std_logic;
signal \N__42045\ : std_logic;
signal \N__42042\ : std_logic;
signal \N__42039\ : std_logic;
signal \N__42036\ : std_logic;
signal \N__42033\ : std_logic;
signal \N__42026\ : std_logic;
signal \N__42023\ : std_logic;
signal \N__42020\ : std_logic;
signal \N__42017\ : std_logic;
signal \N__42016\ : std_logic;
signal \N__42013\ : std_logic;
signal \N__42012\ : std_logic;
signal \N__42011\ : std_logic;
signal \N__42010\ : std_logic;
signal \N__42007\ : std_logic;
signal \N__42004\ : std_logic;
signal \N__42001\ : std_logic;
signal \N__41998\ : std_logic;
signal \N__41995\ : std_logic;
signal \N__41992\ : std_logic;
signal \N__41987\ : std_logic;
signal \N__41984\ : std_logic;
signal \N__41981\ : std_logic;
signal \N__41978\ : std_logic;
signal \N__41975\ : std_logic;
signal \N__41970\ : std_logic;
signal \N__41963\ : std_logic;
signal \N__41960\ : std_logic;
signal \N__41959\ : std_logic;
signal \N__41958\ : std_logic;
signal \N__41955\ : std_logic;
signal \N__41952\ : std_logic;
signal \N__41949\ : std_logic;
signal \N__41946\ : std_logic;
signal \N__41939\ : std_logic;
signal \N__41936\ : std_logic;
signal \N__41935\ : std_logic;
signal \N__41934\ : std_logic;
signal \N__41931\ : std_logic;
signal \N__41928\ : std_logic;
signal \N__41925\ : std_logic;
signal \N__41922\ : std_logic;
signal \N__41915\ : std_logic;
signal \N__41912\ : std_logic;
signal \N__41911\ : std_logic;
signal \N__41910\ : std_logic;
signal \N__41907\ : std_logic;
signal \N__41904\ : std_logic;
signal \N__41901\ : std_logic;
signal \N__41898\ : std_logic;
signal \N__41891\ : std_logic;
signal \N__41888\ : std_logic;
signal \N__41887\ : std_logic;
signal \N__41886\ : std_logic;
signal \N__41883\ : std_logic;
signal \N__41880\ : std_logic;
signal \N__41877\ : std_logic;
signal \N__41874\ : std_logic;
signal \N__41867\ : std_logic;
signal \N__41864\ : std_logic;
signal \N__41863\ : std_logic;
signal \N__41862\ : std_logic;
signal \N__41859\ : std_logic;
signal \N__41856\ : std_logic;
signal \N__41853\ : std_logic;
signal \N__41850\ : std_logic;
signal \N__41843\ : std_logic;
signal \N__41840\ : std_logic;
signal \N__41837\ : std_logic;
signal \N__41836\ : std_logic;
signal \N__41833\ : std_logic;
signal \N__41830\ : std_logic;
signal \N__41825\ : std_logic;
signal \N__41822\ : std_logic;
signal \N__41821\ : std_logic;
signal \N__41820\ : std_logic;
signal \N__41817\ : std_logic;
signal \N__41814\ : std_logic;
signal \N__41811\ : std_logic;
signal \N__41808\ : std_logic;
signal \N__41801\ : std_logic;
signal \N__41798\ : std_logic;
signal \N__41797\ : std_logic;
signal \N__41794\ : std_logic;
signal \N__41791\ : std_logic;
signal \N__41788\ : std_logic;
signal \N__41785\ : std_logic;
signal \N__41780\ : std_logic;
signal \N__41777\ : std_logic;
signal \N__41776\ : std_logic;
signal \N__41775\ : std_logic;
signal \N__41772\ : std_logic;
signal \N__41769\ : std_logic;
signal \N__41766\ : std_logic;
signal \N__41763\ : std_logic;
signal \N__41756\ : std_logic;
signal \N__41753\ : std_logic;
signal \N__41752\ : std_logic;
signal \N__41749\ : std_logic;
signal \N__41746\ : std_logic;
signal \N__41743\ : std_logic;
signal \N__41740\ : std_logic;
signal \N__41735\ : std_logic;
signal \N__41732\ : std_logic;
signal \N__41731\ : std_logic;
signal \N__41730\ : std_logic;
signal \N__41727\ : std_logic;
signal \N__41724\ : std_logic;
signal \N__41721\ : std_logic;
signal \N__41718\ : std_logic;
signal \N__41711\ : std_logic;
signal \N__41708\ : std_logic;
signal \N__41707\ : std_logic;
signal \N__41706\ : std_logic;
signal \N__41705\ : std_logic;
signal \N__41702\ : std_logic;
signal \N__41699\ : std_logic;
signal \N__41698\ : std_logic;
signal \N__41693\ : std_logic;
signal \N__41688\ : std_logic;
signal \N__41685\ : std_logic;
signal \N__41682\ : std_logic;
signal \N__41679\ : std_logic;
signal \N__41674\ : std_logic;
signal \N__41669\ : std_logic;
signal \N__41666\ : std_logic;
signal \N__41665\ : std_logic;
signal \N__41664\ : std_logic;
signal \N__41661\ : std_logic;
signal \N__41658\ : std_logic;
signal \N__41655\ : std_logic;
signal \N__41652\ : std_logic;
signal \N__41645\ : std_logic;
signal \N__41644\ : std_logic;
signal \N__41643\ : std_logic;
signal \N__41642\ : std_logic;
signal \N__41639\ : std_logic;
signal \N__41638\ : std_logic;
signal \N__41635\ : std_logic;
signal \N__41632\ : std_logic;
signal \N__41629\ : std_logic;
signal \N__41624\ : std_logic;
signal \N__41619\ : std_logic;
signal \N__41614\ : std_logic;
signal \N__41611\ : std_logic;
signal \N__41608\ : std_logic;
signal \N__41603\ : std_logic;
signal \N__41600\ : std_logic;
signal \N__41599\ : std_logic;
signal \N__41598\ : std_logic;
signal \N__41595\ : std_logic;
signal \N__41592\ : std_logic;
signal \N__41589\ : std_logic;
signal \N__41586\ : std_logic;
signal \N__41579\ : std_logic;
signal \N__41576\ : std_logic;
signal \N__41575\ : std_logic;
signal \N__41574\ : std_logic;
signal \N__41571\ : std_logic;
signal \N__41568\ : std_logic;
signal \N__41565\ : std_logic;
signal \N__41562\ : std_logic;
signal \N__41555\ : std_logic;
signal \N__41554\ : std_logic;
signal \N__41551\ : std_logic;
signal \N__41550\ : std_logic;
signal \N__41547\ : std_logic;
signal \N__41544\ : std_logic;
signal \N__41541\ : std_logic;
signal \N__41538\ : std_logic;
signal \N__41535\ : std_logic;
signal \N__41530\ : std_logic;
signal \N__41527\ : std_logic;
signal \N__41524\ : std_logic;
signal \N__41519\ : std_logic;
signal \N__41516\ : std_logic;
signal \N__41515\ : std_logic;
signal \N__41514\ : std_logic;
signal \N__41511\ : std_logic;
signal \N__41508\ : std_logic;
signal \N__41505\ : std_logic;
signal \N__41502\ : std_logic;
signal \N__41495\ : std_logic;
signal \N__41492\ : std_logic;
signal \N__41489\ : std_logic;
signal \N__41488\ : std_logic;
signal \N__41487\ : std_logic;
signal \N__41484\ : std_logic;
signal \N__41479\ : std_logic;
signal \N__41474\ : std_logic;
signal \N__41471\ : std_logic;
signal \N__41468\ : std_logic;
signal \N__41467\ : std_logic;
signal \N__41466\ : std_logic;
signal \N__41463\ : std_logic;
signal \N__41460\ : std_logic;
signal \N__41457\ : std_logic;
signal \N__41454\ : std_logic;
signal \N__41447\ : std_logic;
signal \N__41446\ : std_logic;
signal \N__41443\ : std_logic;
signal \N__41442\ : std_logic;
signal \N__41439\ : std_logic;
signal \N__41436\ : std_logic;
signal \N__41431\ : std_logic;
signal \N__41428\ : std_logic;
signal \N__41425\ : std_logic;
signal \N__41420\ : std_logic;
signal \N__41417\ : std_logic;
signal \N__41416\ : std_logic;
signal \N__41415\ : std_logic;
signal \N__41412\ : std_logic;
signal \N__41409\ : std_logic;
signal \N__41406\ : std_logic;
signal \N__41403\ : std_logic;
signal \N__41396\ : std_logic;
signal \N__41395\ : std_logic;
signal \N__41392\ : std_logic;
signal \N__41391\ : std_logic;
signal \N__41388\ : std_logic;
signal \N__41385\ : std_logic;
signal \N__41380\ : std_logic;
signal \N__41377\ : std_logic;
signal \N__41374\ : std_logic;
signal \N__41369\ : std_logic;
signal \N__41366\ : std_logic;
signal \N__41363\ : std_logic;
signal \N__41362\ : std_logic;
signal \N__41361\ : std_logic;
signal \N__41358\ : std_logic;
signal \N__41355\ : std_logic;
signal \N__41352\ : std_logic;
signal \N__41349\ : std_logic;
signal \N__41342\ : std_logic;
signal \N__41339\ : std_logic;
signal \N__41336\ : std_logic;
signal \N__41333\ : std_logic;
signal \N__41330\ : std_logic;
signal \N__41327\ : std_logic;
signal \N__41324\ : std_logic;
signal \N__41321\ : std_logic;
signal \N__41318\ : std_logic;
signal \N__41315\ : std_logic;
signal \N__41312\ : std_logic;
signal \N__41311\ : std_logic;
signal \N__41308\ : std_logic;
signal \N__41305\ : std_logic;
signal \N__41304\ : std_logic;
signal \N__41301\ : std_logic;
signal \N__41298\ : std_logic;
signal \N__41295\ : std_logic;
signal \N__41288\ : std_logic;
signal \N__41285\ : std_logic;
signal \N__41282\ : std_logic;
signal \N__41279\ : std_logic;
signal \N__41276\ : std_logic;
signal \N__41273\ : std_logic;
signal \N__41272\ : std_logic;
signal \N__41269\ : std_logic;
signal \N__41266\ : std_logic;
signal \N__41263\ : std_logic;
signal \N__41260\ : std_logic;
signal \N__41257\ : std_logic;
signal \N__41254\ : std_logic;
signal \N__41249\ : std_logic;
signal \N__41248\ : std_logic;
signal \N__41247\ : std_logic;
signal \N__41244\ : std_logic;
signal \N__41241\ : std_logic;
signal \N__41238\ : std_logic;
signal \N__41231\ : std_logic;
signal \N__41228\ : std_logic;
signal \N__41227\ : std_logic;
signal \N__41226\ : std_logic;
signal \N__41223\ : std_logic;
signal \N__41220\ : std_logic;
signal \N__41217\ : std_logic;
signal \N__41214\ : std_logic;
signal \N__41207\ : std_logic;
signal \N__41206\ : std_logic;
signal \N__41205\ : std_logic;
signal \N__41202\ : std_logic;
signal \N__41199\ : std_logic;
signal \N__41196\ : std_logic;
signal \N__41193\ : std_logic;
signal \N__41190\ : std_logic;
signal \N__41187\ : std_logic;
signal \N__41184\ : std_logic;
signal \N__41181\ : std_logic;
signal \N__41174\ : std_logic;
signal \N__41171\ : std_logic;
signal \N__41170\ : std_logic;
signal \N__41169\ : std_logic;
signal \N__41166\ : std_logic;
signal \N__41163\ : std_logic;
signal \N__41160\ : std_logic;
signal \N__41157\ : std_logic;
signal \N__41150\ : std_logic;
signal \N__41147\ : std_logic;
signal \N__41144\ : std_logic;
signal \N__41141\ : std_logic;
signal \N__41138\ : std_logic;
signal \N__41135\ : std_logic;
signal \N__41132\ : std_logic;
signal \N__41129\ : std_logic;
signal \N__41126\ : std_logic;
signal \N__41123\ : std_logic;
signal \N__41120\ : std_logic;
signal \N__41117\ : std_logic;
signal \N__41114\ : std_logic;
signal \N__41111\ : std_logic;
signal \N__41108\ : std_logic;
signal \N__41105\ : std_logic;
signal \N__41102\ : std_logic;
signal \N__41099\ : std_logic;
signal \N__41096\ : std_logic;
signal \N__41093\ : std_logic;
signal \N__41090\ : std_logic;
signal \N__41087\ : std_logic;
signal \N__41084\ : std_logic;
signal \N__41081\ : std_logic;
signal \N__41080\ : std_logic;
signal \N__41077\ : std_logic;
signal \N__41074\ : std_logic;
signal \N__41073\ : std_logic;
signal \N__41070\ : std_logic;
signal \N__41067\ : std_logic;
signal \N__41064\ : std_logic;
signal \N__41057\ : std_logic;
signal \N__41054\ : std_logic;
signal \N__41051\ : std_logic;
signal \N__41048\ : std_logic;
signal \N__41045\ : std_logic;
signal \N__41042\ : std_logic;
signal \N__41039\ : std_logic;
signal \N__41036\ : std_logic;
signal \N__41033\ : std_logic;
signal \N__41030\ : std_logic;
signal \N__41027\ : std_logic;
signal \N__41026\ : std_logic;
signal \N__41023\ : std_logic;
signal \N__41020\ : std_logic;
signal \N__41019\ : std_logic;
signal \N__41014\ : std_logic;
signal \N__41011\ : std_logic;
signal \N__41006\ : std_logic;
signal \N__41003\ : std_logic;
signal \N__41000\ : std_logic;
signal \N__40997\ : std_logic;
signal \N__40994\ : std_logic;
signal \N__40991\ : std_logic;
signal \N__40988\ : std_logic;
signal \N__40985\ : std_logic;
signal \N__40982\ : std_logic;
signal \N__40979\ : std_logic;
signal \N__40976\ : std_logic;
signal \N__40973\ : std_logic;
signal \N__40970\ : std_logic;
signal \N__40967\ : std_logic;
signal \N__40964\ : std_logic;
signal \N__40961\ : std_logic;
signal \N__40958\ : std_logic;
signal \N__40955\ : std_logic;
signal \N__40952\ : std_logic;
signal \N__40949\ : std_logic;
signal \N__40946\ : std_logic;
signal \N__40943\ : std_logic;
signal \N__40940\ : std_logic;
signal \N__40937\ : std_logic;
signal \N__40934\ : std_logic;
signal \N__40931\ : std_logic;
signal \N__40928\ : std_logic;
signal \N__40925\ : std_logic;
signal \N__40922\ : std_logic;
signal \N__40919\ : std_logic;
signal \N__40916\ : std_logic;
signal \N__40913\ : std_logic;
signal \N__40910\ : std_logic;
signal \N__40907\ : std_logic;
signal \N__40904\ : std_logic;
signal \N__40901\ : std_logic;
signal \N__40898\ : std_logic;
signal \N__40895\ : std_logic;
signal \N__40892\ : std_logic;
signal \N__40889\ : std_logic;
signal \N__40886\ : std_logic;
signal \N__40883\ : std_logic;
signal \N__40880\ : std_logic;
signal \N__40877\ : std_logic;
signal \N__40874\ : std_logic;
signal \N__40871\ : std_logic;
signal \N__40868\ : std_logic;
signal \N__40865\ : std_logic;
signal \N__40862\ : std_logic;
signal \N__40859\ : std_logic;
signal \N__40856\ : std_logic;
signal \N__40853\ : std_logic;
signal \N__40852\ : std_logic;
signal \N__40851\ : std_logic;
signal \N__40850\ : std_logic;
signal \N__40849\ : std_logic;
signal \N__40848\ : std_logic;
signal \N__40847\ : std_logic;
signal \N__40846\ : std_logic;
signal \N__40845\ : std_logic;
signal \N__40844\ : std_logic;
signal \N__40843\ : std_logic;
signal \N__40842\ : std_logic;
signal \N__40839\ : std_logic;
signal \N__40832\ : std_logic;
signal \N__40831\ : std_logic;
signal \N__40822\ : std_logic;
signal \N__40817\ : std_logic;
signal \N__40812\ : std_logic;
signal \N__40809\ : std_logic;
signal \N__40806\ : std_logic;
signal \N__40803\ : std_logic;
signal \N__40800\ : std_logic;
signal \N__40795\ : std_logic;
signal \N__40794\ : std_logic;
signal \N__40793\ : std_logic;
signal \N__40792\ : std_logic;
signal \N__40791\ : std_logic;
signal \N__40790\ : std_logic;
signal \N__40789\ : std_logic;
signal \N__40788\ : std_logic;
signal \N__40787\ : std_logic;
signal \N__40786\ : std_logic;
signal \N__40785\ : std_logic;
signal \N__40784\ : std_logic;
signal \N__40781\ : std_logic;
signal \N__40778\ : std_logic;
signal \N__40775\ : std_logic;
signal \N__40772\ : std_logic;
signal \N__40769\ : std_logic;
signal \N__40762\ : std_logic;
signal \N__40745\ : std_logic;
signal \N__40730\ : std_logic;
signal \N__40729\ : std_logic;
signal \N__40728\ : std_logic;
signal \N__40725\ : std_logic;
signal \N__40724\ : std_logic;
signal \N__40723\ : std_logic;
signal \N__40722\ : std_logic;
signal \N__40721\ : std_logic;
signal \N__40720\ : std_logic;
signal \N__40719\ : std_logic;
signal \N__40718\ : std_logic;
signal \N__40717\ : std_logic;
signal \N__40716\ : std_logic;
signal \N__40713\ : std_logic;
signal \N__40710\ : std_logic;
signal \N__40709\ : std_logic;
signal \N__40706\ : std_logic;
signal \N__40703\ : std_logic;
signal \N__40702\ : std_logic;
signal \N__40701\ : std_logic;
signal \N__40700\ : std_logic;
signal \N__40699\ : std_logic;
signal \N__40698\ : std_logic;
signal \N__40697\ : std_logic;
signal \N__40696\ : std_logic;
signal \N__40695\ : std_logic;
signal \N__40694\ : std_logic;
signal \N__40693\ : std_logic;
signal \N__40688\ : std_logic;
signal \N__40685\ : std_logic;
signal \N__40684\ : std_logic;
signal \N__40683\ : std_logic;
signal \N__40682\ : std_logic;
signal \N__40681\ : std_logic;
signal \N__40672\ : std_logic;
signal \N__40671\ : std_logic;
signal \N__40670\ : std_logic;
signal \N__40667\ : std_logic;
signal \N__40666\ : std_logic;
signal \N__40659\ : std_logic;
signal \N__40654\ : std_logic;
signal \N__40653\ : std_logic;
signal \N__40652\ : std_logic;
signal \N__40649\ : std_logic;
signal \N__40632\ : std_logic;
signal \N__40629\ : std_logic;
signal \N__40626\ : std_logic;
signal \N__40615\ : std_logic;
signal \N__40612\ : std_logic;
signal \N__40603\ : std_logic;
signal \N__40600\ : std_logic;
signal \N__40597\ : std_logic;
signal \N__40592\ : std_logic;
signal \N__40587\ : std_logic;
signal \N__40582\ : std_logic;
signal \N__40577\ : std_logic;
signal \N__40570\ : std_logic;
signal \N__40559\ : std_logic;
signal \N__40558\ : std_logic;
signal \N__40555\ : std_logic;
signal \N__40554\ : std_logic;
signal \N__40553\ : std_logic;
signal \N__40552\ : std_logic;
signal \N__40551\ : std_logic;
signal \N__40548\ : std_logic;
signal \N__40547\ : std_logic;
signal \N__40546\ : std_logic;
signal \N__40541\ : std_logic;
signal \N__40538\ : std_logic;
signal \N__40537\ : std_logic;
signal \N__40536\ : std_logic;
signal \N__40535\ : std_logic;
signal \N__40534\ : std_logic;
signal \N__40533\ : std_logic;
signal \N__40532\ : std_logic;
signal \N__40531\ : std_logic;
signal \N__40530\ : std_logic;
signal \N__40529\ : std_logic;
signal \N__40526\ : std_logic;
signal \N__40525\ : std_logic;
signal \N__40524\ : std_logic;
signal \N__40521\ : std_logic;
signal \N__40520\ : std_logic;
signal \N__40519\ : std_logic;
signal \N__40512\ : std_logic;
signal \N__40511\ : std_logic;
signal \N__40510\ : std_logic;
signal \N__40509\ : std_logic;
signal \N__40506\ : std_logic;
signal \N__40503\ : std_logic;
signal \N__40502\ : std_logic;
signal \N__40499\ : std_logic;
signal \N__40498\ : std_logic;
signal \N__40497\ : std_logic;
signal \N__40496\ : std_logic;
signal \N__40493\ : std_logic;
signal \N__40490\ : std_logic;
signal \N__40489\ : std_logic;
signal \N__40488\ : std_logic;
signal \N__40487\ : std_logic;
signal \N__40486\ : std_logic;
signal \N__40485\ : std_logic;
signal \N__40482\ : std_logic;
signal \N__40479\ : std_logic;
signal \N__40478\ : std_logic;
signal \N__40477\ : std_logic;
signal \N__40476\ : std_logic;
signal \N__40475\ : std_logic;
signal \N__40472\ : std_logic;
signal \N__40471\ : std_logic;
signal \N__40468\ : std_logic;
signal \N__40465\ : std_logic;
signal \N__40464\ : std_logic;
signal \N__40463\ : std_logic;
signal \N__40462\ : std_logic;
signal \N__40461\ : std_logic;
signal \N__40458\ : std_logic;
signal \N__40445\ : std_logic;
signal \N__40442\ : std_logic;
signal \N__40437\ : std_logic;
signal \N__40434\ : std_logic;
signal \N__40429\ : std_logic;
signal \N__40418\ : std_logic;
signal \N__40407\ : std_logic;
signal \N__40390\ : std_logic;
signal \N__40385\ : std_logic;
signal \N__40374\ : std_logic;
signal \N__40371\ : std_logic;
signal \N__40362\ : std_logic;
signal \N__40359\ : std_logic;
signal \N__40358\ : std_logic;
signal \N__40355\ : std_logic;
signal \N__40346\ : std_logic;
signal \N__40343\ : std_logic;
signal \N__40340\ : std_logic;
signal \N__40335\ : std_logic;
signal \N__40332\ : std_logic;
signal \N__40329\ : std_logic;
signal \N__40326\ : std_logic;
signal \N__40323\ : std_logic;
signal \N__40318\ : std_logic;
signal \N__40307\ : std_logic;
signal \N__40304\ : std_logic;
signal \N__40301\ : std_logic;
signal \N__40300\ : std_logic;
signal \N__40297\ : std_logic;
signal \N__40294\ : std_logic;
signal \N__40291\ : std_logic;
signal \N__40286\ : std_logic;
signal \N__40283\ : std_logic;
signal \N__40280\ : std_logic;
signal \N__40279\ : std_logic;
signal \N__40276\ : std_logic;
signal \N__40273\ : std_logic;
signal \N__40270\ : std_logic;
signal \N__40265\ : std_logic;
signal \N__40262\ : std_logic;
signal \N__40259\ : std_logic;
signal \N__40258\ : std_logic;
signal \N__40255\ : std_logic;
signal \N__40252\ : std_logic;
signal \N__40249\ : std_logic;
signal \N__40244\ : std_logic;
signal \N__40243\ : std_logic;
signal \N__40242\ : std_logic;
signal \N__40241\ : std_logic;
signal \N__40240\ : std_logic;
signal \N__40239\ : std_logic;
signal \N__40238\ : std_logic;
signal \N__40237\ : std_logic;
signal \N__40236\ : std_logic;
signal \N__40235\ : std_logic;
signal \N__40234\ : std_logic;
signal \N__40233\ : std_logic;
signal \N__40232\ : std_logic;
signal \N__40231\ : std_logic;
signal \N__40230\ : std_logic;
signal \N__40229\ : std_logic;
signal \N__40220\ : std_logic;
signal \N__40203\ : std_logic;
signal \N__40202\ : std_logic;
signal \N__40201\ : std_logic;
signal \N__40200\ : std_logic;
signal \N__40199\ : std_logic;
signal \N__40198\ : std_logic;
signal \N__40197\ : std_logic;
signal \N__40194\ : std_logic;
signal \N__40193\ : std_logic;
signal \N__40188\ : std_logic;
signal \N__40185\ : std_logic;
signal \N__40184\ : std_logic;
signal \N__40179\ : std_logic;
signal \N__40176\ : std_logic;
signal \N__40165\ : std_logic;
signal \N__40162\ : std_logic;
signal \N__40159\ : std_logic;
signal \N__40156\ : std_logic;
signal \N__40151\ : std_logic;
signal \N__40148\ : std_logic;
signal \N__40145\ : std_logic;
signal \N__40136\ : std_logic;
signal \N__40127\ : std_logic;
signal \N__40126\ : std_logic;
signal \N__40125\ : std_logic;
signal \N__40124\ : std_logic;
signal \N__40123\ : std_logic;
signal \N__40122\ : std_logic;
signal \N__40121\ : std_logic;
signal \N__40120\ : std_logic;
signal \N__40117\ : std_logic;
signal \N__40116\ : std_logic;
signal \N__40115\ : std_logic;
signal \N__40114\ : std_logic;
signal \N__40113\ : std_logic;
signal \N__40110\ : std_logic;
signal \N__40107\ : std_logic;
signal \N__40104\ : std_logic;
signal \N__40101\ : std_logic;
signal \N__40100\ : std_logic;
signal \N__40097\ : std_logic;
signal \N__40094\ : std_logic;
signal \N__40091\ : std_logic;
signal \N__40090\ : std_logic;
signal \N__40087\ : std_logic;
signal \N__40070\ : std_logic;
signal \N__40067\ : std_logic;
signal \N__40066\ : std_logic;
signal \N__40065\ : std_logic;
signal \N__40064\ : std_logic;
signal \N__40063\ : std_logic;
signal \N__40062\ : std_logic;
signal \N__40061\ : std_logic;
signal \N__40060\ : std_logic;
signal \N__40051\ : std_logic;
signal \N__40048\ : std_logic;
signal \N__40045\ : std_logic;
signal \N__40040\ : std_logic;
signal \N__40029\ : std_logic;
signal \N__40026\ : std_logic;
signal \N__40025\ : std_logic;
signal \N__40024\ : std_logic;
signal \N__40021\ : std_logic;
signal \N__40018\ : std_logic;
signal \N__40013\ : std_logic;
signal \N__40010\ : std_logic;
signal \N__40007\ : std_logic;
signal \N__40006\ : std_logic;
signal \N__40001\ : std_logic;
signal \N__39996\ : std_logic;
signal \N__39991\ : std_logic;
signal \N__39988\ : std_logic;
signal \N__39985\ : std_logic;
signal \N__39974\ : std_logic;
signal \N__39971\ : std_logic;
signal \N__39968\ : std_logic;
signal \N__39965\ : std_logic;
signal \N__39964\ : std_logic;
signal \N__39963\ : std_logic;
signal \N__39962\ : std_logic;
signal \N__39961\ : std_logic;
signal \N__39960\ : std_logic;
signal \N__39959\ : std_logic;
signal \N__39958\ : std_logic;
signal \N__39957\ : std_logic;
signal \N__39956\ : std_logic;
signal \N__39955\ : std_logic;
signal \N__39954\ : std_logic;
signal \N__39953\ : std_logic;
signal \N__39952\ : std_logic;
signal \N__39951\ : std_logic;
signal \N__39950\ : std_logic;
signal \N__39949\ : std_logic;
signal \N__39948\ : std_logic;
signal \N__39939\ : std_logic;
signal \N__39938\ : std_logic;
signal \N__39937\ : std_logic;
signal \N__39936\ : std_logic;
signal \N__39933\ : std_logic;
signal \N__39930\ : std_logic;
signal \N__39927\ : std_logic;
signal \N__39924\ : std_logic;
signal \N__39923\ : std_logic;
signal \N__39920\ : std_logic;
signal \N__39917\ : std_logic;
signal \N__39916\ : std_logic;
signal \N__39915\ : std_logic;
signal \N__39898\ : std_logic;
signal \N__39895\ : std_logic;
signal \N__39892\ : std_logic;
signal \N__39881\ : std_logic;
signal \N__39878\ : std_logic;
signal \N__39875\ : std_logic;
signal \N__39870\ : std_logic;
signal \N__39865\ : std_logic;
signal \N__39862\ : std_logic;
signal \N__39859\ : std_logic;
signal \N__39856\ : std_logic;
signal \N__39847\ : std_logic;
signal \N__39836\ : std_logic;
signal \N__39833\ : std_logic;
signal \N__39832\ : std_logic;
signal \N__39829\ : std_logic;
signal \N__39826\ : std_logic;
signal \N__39823\ : std_logic;
signal \N__39818\ : std_logic;
signal \N__39817\ : std_logic;
signal \N__39814\ : std_logic;
signal \N__39811\ : std_logic;
signal \N__39808\ : std_logic;
signal \N__39805\ : std_logic;
signal \N__39802\ : std_logic;
signal \N__39801\ : std_logic;
signal \N__39798\ : std_logic;
signal \N__39795\ : std_logic;
signal \N__39792\ : std_logic;
signal \N__39789\ : std_logic;
signal \N__39784\ : std_logic;
signal \N__39779\ : std_logic;
signal \N__39776\ : std_logic;
signal \N__39773\ : std_logic;
signal \N__39770\ : std_logic;
signal \N__39767\ : std_logic;
signal \N__39766\ : std_logic;
signal \N__39763\ : std_logic;
signal \N__39760\ : std_logic;
signal \N__39759\ : std_logic;
signal \N__39758\ : std_logic;
signal \N__39755\ : std_logic;
signal \N__39752\ : std_logic;
signal \N__39749\ : std_logic;
signal \N__39746\ : std_logic;
signal \N__39743\ : std_logic;
signal \N__39740\ : std_logic;
signal \N__39737\ : std_logic;
signal \N__39728\ : std_logic;
signal \N__39725\ : std_logic;
signal \N__39724\ : std_logic;
signal \N__39723\ : std_logic;
signal \N__39722\ : std_logic;
signal \N__39719\ : std_logic;
signal \N__39716\ : std_logic;
signal \N__39713\ : std_logic;
signal \N__39712\ : std_logic;
signal \N__39709\ : std_logic;
signal \N__39704\ : std_logic;
signal \N__39701\ : std_logic;
signal \N__39698\ : std_logic;
signal \N__39695\ : std_logic;
signal \N__39690\ : std_logic;
signal \N__39687\ : std_logic;
signal \N__39682\ : std_logic;
signal \N__39677\ : std_logic;
signal \N__39674\ : std_logic;
signal \N__39673\ : std_logic;
signal \N__39670\ : std_logic;
signal \N__39667\ : std_logic;
signal \N__39664\ : std_logic;
signal \N__39659\ : std_logic;
signal \N__39656\ : std_logic;
signal \N__39655\ : std_logic;
signal \N__39652\ : std_logic;
signal \N__39649\ : std_logic;
signal \N__39646\ : std_logic;
signal \N__39641\ : std_logic;
signal \N__39638\ : std_logic;
signal \N__39635\ : std_logic;
signal \N__39634\ : std_logic;
signal \N__39631\ : std_logic;
signal \N__39628\ : std_logic;
signal \N__39625\ : std_logic;
signal \N__39620\ : std_logic;
signal \N__39619\ : std_logic;
signal \N__39616\ : std_logic;
signal \N__39613\ : std_logic;
signal \N__39608\ : std_logic;
signal \N__39607\ : std_logic;
signal \N__39604\ : std_logic;
signal \N__39601\ : std_logic;
signal \N__39596\ : std_logic;
signal \N__39593\ : std_logic;
signal \N__39592\ : std_logic;
signal \N__39591\ : std_logic;
signal \N__39588\ : std_logic;
signal \N__39585\ : std_logic;
signal \N__39582\ : std_logic;
signal \N__39581\ : std_logic;
signal \N__39578\ : std_logic;
signal \N__39575\ : std_logic;
signal \N__39572\ : std_logic;
signal \N__39569\ : std_logic;
signal \N__39566\ : std_logic;
signal \N__39563\ : std_logic;
signal \N__39560\ : std_logic;
signal \N__39551\ : std_logic;
signal \N__39550\ : std_logic;
signal \N__39549\ : std_logic;
signal \N__39548\ : std_logic;
signal \N__39547\ : std_logic;
signal \N__39546\ : std_logic;
signal \N__39545\ : std_logic;
signal \N__39544\ : std_logic;
signal \N__39543\ : std_logic;
signal \N__39542\ : std_logic;
signal \N__39541\ : std_logic;
signal \N__39540\ : std_logic;
signal \N__39539\ : std_logic;
signal \N__39538\ : std_logic;
signal \N__39537\ : std_logic;
signal \N__39536\ : std_logic;
signal \N__39527\ : std_logic;
signal \N__39518\ : std_logic;
signal \N__39517\ : std_logic;
signal \N__39516\ : std_logic;
signal \N__39515\ : std_logic;
signal \N__39514\ : std_logic;
signal \N__39513\ : std_logic;
signal \N__39512\ : std_logic;
signal \N__39511\ : std_logic;
signal \N__39510\ : std_logic;
signal \N__39509\ : std_logic;
signal \N__39508\ : std_logic;
signal \N__39507\ : std_logic;
signal \N__39506\ : std_logic;
signal \N__39505\ : std_logic;
signal \N__39504\ : std_logic;
signal \N__39495\ : std_logic;
signal \N__39486\ : std_logic;
signal \N__39481\ : std_logic;
signal \N__39472\ : std_logic;
signal \N__39467\ : std_logic;
signal \N__39458\ : std_logic;
signal \N__39449\ : std_logic;
signal \N__39444\ : std_logic;
signal \N__39435\ : std_logic;
signal \N__39428\ : std_logic;
signal \N__39425\ : std_logic;
signal \N__39424\ : std_logic;
signal \N__39423\ : std_logic;
signal \N__39420\ : std_logic;
signal \N__39417\ : std_logic;
signal \N__39414\ : std_logic;
signal \N__39411\ : std_logic;
signal \N__39406\ : std_logic;
signal \N__39405\ : std_logic;
signal \N__39402\ : std_logic;
signal \N__39399\ : std_logic;
signal \N__39396\ : std_logic;
signal \N__39389\ : std_logic;
signal \N__39386\ : std_logic;
signal \N__39383\ : std_logic;
signal \N__39380\ : std_logic;
signal \N__39377\ : std_logic;
signal \N__39374\ : std_logic;
signal \N__39371\ : std_logic;
signal \N__39368\ : std_logic;
signal \N__39365\ : std_logic;
signal \N__39364\ : std_logic;
signal \N__39361\ : std_logic;
signal \N__39358\ : std_logic;
signal \N__39353\ : std_logic;
signal \N__39352\ : std_logic;
signal \N__39349\ : std_logic;
signal \N__39346\ : std_logic;
signal \N__39343\ : std_logic;
signal \N__39340\ : std_logic;
signal \N__39337\ : std_logic;
signal \N__39332\ : std_logic;
signal \N__39329\ : std_logic;
signal \N__39326\ : std_logic;
signal \N__39323\ : std_logic;
signal \N__39320\ : std_logic;
signal \N__39317\ : std_logic;
signal \N__39314\ : std_logic;
signal \N__39311\ : std_logic;
signal \N__39308\ : std_logic;
signal \N__39305\ : std_logic;
signal \N__39302\ : std_logic;
signal \N__39299\ : std_logic;
signal \N__39296\ : std_logic;
signal \N__39293\ : std_logic;
signal \N__39290\ : std_logic;
signal \N__39287\ : std_logic;
signal \N__39284\ : std_logic;
signal \N__39281\ : std_logic;
signal \N__39278\ : std_logic;
signal \N__39275\ : std_logic;
signal \N__39272\ : std_logic;
signal \N__39269\ : std_logic;
signal \N__39266\ : std_logic;
signal \N__39263\ : std_logic;
signal \N__39260\ : std_logic;
signal \N__39257\ : std_logic;
signal \N__39254\ : std_logic;
signal \N__39251\ : std_logic;
signal \N__39248\ : std_logic;
signal \N__39245\ : std_logic;
signal \N__39242\ : std_logic;
signal \N__39241\ : std_logic;
signal \N__39238\ : std_logic;
signal \N__39235\ : std_logic;
signal \N__39230\ : std_logic;
signal \N__39227\ : std_logic;
signal \N__39224\ : std_logic;
signal \N__39221\ : std_logic;
signal \N__39220\ : std_logic;
signal \N__39219\ : std_logic;
signal \N__39216\ : std_logic;
signal \N__39213\ : std_logic;
signal \N__39210\ : std_logic;
signal \N__39207\ : std_logic;
signal \N__39206\ : std_logic;
signal \N__39205\ : std_logic;
signal \N__39202\ : std_logic;
signal \N__39201\ : std_logic;
signal \N__39198\ : std_logic;
signal \N__39195\ : std_logic;
signal \N__39190\ : std_logic;
signal \N__39187\ : std_logic;
signal \N__39184\ : std_logic;
signal \N__39179\ : std_logic;
signal \N__39176\ : std_logic;
signal \N__39167\ : std_logic;
signal \N__39164\ : std_logic;
signal \N__39161\ : std_logic;
signal \N__39158\ : std_logic;
signal \N__39155\ : std_logic;
signal \N__39152\ : std_logic;
signal \N__39149\ : std_logic;
signal \N__39146\ : std_logic;
signal \N__39143\ : std_logic;
signal \N__39140\ : std_logic;
signal \N__39139\ : std_logic;
signal \N__39136\ : std_logic;
signal \N__39133\ : std_logic;
signal \N__39128\ : std_logic;
signal \N__39127\ : std_logic;
signal \N__39126\ : std_logic;
signal \N__39123\ : std_logic;
signal \N__39120\ : std_logic;
signal \N__39117\ : std_logic;
signal \N__39114\ : std_logic;
signal \N__39111\ : std_logic;
signal \N__39104\ : std_logic;
signal \N__39103\ : std_logic;
signal \N__39102\ : std_logic;
signal \N__39101\ : std_logic;
signal \N__39098\ : std_logic;
signal \N__39095\ : std_logic;
signal \N__39090\ : std_logic;
signal \N__39087\ : std_logic;
signal \N__39080\ : std_logic;
signal \N__39077\ : std_logic;
signal \N__39074\ : std_logic;
signal \N__39073\ : std_logic;
signal \N__39070\ : std_logic;
signal \N__39067\ : std_logic;
signal \N__39062\ : std_logic;
signal \N__39059\ : std_logic;
signal \N__39056\ : std_logic;
signal \N__39055\ : std_logic;
signal \N__39052\ : std_logic;
signal \N__39049\ : std_logic;
signal \N__39044\ : std_logic;
signal \N__39041\ : std_logic;
signal \N__39038\ : std_logic;
signal \N__39037\ : std_logic;
signal \N__39034\ : std_logic;
signal \N__39031\ : std_logic;
signal \N__39026\ : std_logic;
signal \N__39023\ : std_logic;
signal \N__39020\ : std_logic;
signal \N__39019\ : std_logic;
signal \N__39016\ : std_logic;
signal \N__39013\ : std_logic;
signal \N__39008\ : std_logic;
signal \N__39005\ : std_logic;
signal \N__39002\ : std_logic;
signal \N__39001\ : std_logic;
signal \N__38998\ : std_logic;
signal \N__38995\ : std_logic;
signal \N__38990\ : std_logic;
signal \N__38987\ : std_logic;
signal \N__38984\ : std_logic;
signal \N__38981\ : std_logic;
signal \N__38978\ : std_logic;
signal \N__38975\ : std_logic;
signal \N__38972\ : std_logic;
signal \N__38969\ : std_logic;
signal \N__38968\ : std_logic;
signal \N__38965\ : std_logic;
signal \N__38962\ : std_logic;
signal \N__38959\ : std_logic;
signal \N__38954\ : std_logic;
signal \N__38951\ : std_logic;
signal \N__38948\ : std_logic;
signal \N__38945\ : std_logic;
signal \N__38944\ : std_logic;
signal \N__38941\ : std_logic;
signal \N__38938\ : std_logic;
signal \N__38933\ : std_logic;
signal \N__38930\ : std_logic;
signal \N__38927\ : std_logic;
signal \N__38926\ : std_logic;
signal \N__38923\ : std_logic;
signal \N__38920\ : std_logic;
signal \N__38915\ : std_logic;
signal \N__38912\ : std_logic;
signal \N__38909\ : std_logic;
signal \N__38908\ : std_logic;
signal \N__38905\ : std_logic;
signal \N__38902\ : std_logic;
signal \N__38897\ : std_logic;
signal \N__38894\ : std_logic;
signal \N__38891\ : std_logic;
signal \N__38890\ : std_logic;
signal \N__38887\ : std_logic;
signal \N__38884\ : std_logic;
signal \N__38879\ : std_logic;
signal \N__38876\ : std_logic;
signal \N__38873\ : std_logic;
signal \N__38872\ : std_logic;
signal \N__38869\ : std_logic;
signal \N__38866\ : std_logic;
signal \N__38861\ : std_logic;
signal \N__38858\ : std_logic;
signal \N__38855\ : std_logic;
signal \N__38852\ : std_logic;
signal \N__38851\ : std_logic;
signal \N__38848\ : std_logic;
signal \N__38845\ : std_logic;
signal \N__38840\ : std_logic;
signal \N__38837\ : std_logic;
signal \N__38834\ : std_logic;
signal \N__38833\ : std_logic;
signal \N__38830\ : std_logic;
signal \N__38827\ : std_logic;
signal \N__38822\ : std_logic;
signal \N__38819\ : std_logic;
signal \N__38816\ : std_logic;
signal \N__38813\ : std_logic;
signal \N__38812\ : std_logic;
signal \N__38809\ : std_logic;
signal \N__38806\ : std_logic;
signal \N__38803\ : std_logic;
signal \N__38800\ : std_logic;
signal \N__38795\ : std_logic;
signal \N__38792\ : std_logic;
signal \N__38789\ : std_logic;
signal \N__38788\ : std_logic;
signal \N__38785\ : std_logic;
signal \N__38782\ : std_logic;
signal \N__38777\ : std_logic;
signal \N__38774\ : std_logic;
signal \N__38771\ : std_logic;
signal \N__38768\ : std_logic;
signal \N__38767\ : std_logic;
signal \N__38764\ : std_logic;
signal \N__38761\ : std_logic;
signal \N__38758\ : std_logic;
signal \N__38753\ : std_logic;
signal \N__38750\ : std_logic;
signal \N__38747\ : std_logic;
signal \N__38744\ : std_logic;
signal \N__38743\ : std_logic;
signal \N__38740\ : std_logic;
signal \N__38737\ : std_logic;
signal \N__38734\ : std_logic;
signal \N__38729\ : std_logic;
signal \N__38726\ : std_logic;
signal \N__38723\ : std_logic;
signal \N__38722\ : std_logic;
signal \N__38719\ : std_logic;
signal \N__38716\ : std_logic;
signal \N__38713\ : std_logic;
signal \N__38708\ : std_logic;
signal \N__38705\ : std_logic;
signal \N__38702\ : std_logic;
signal \N__38699\ : std_logic;
signal \N__38698\ : std_logic;
signal \N__38697\ : std_logic;
signal \N__38692\ : std_logic;
signal \N__38689\ : std_logic;
signal \N__38686\ : std_logic;
signal \N__38683\ : std_logic;
signal \N__38682\ : std_logic;
signal \N__38681\ : std_logic;
signal \N__38680\ : std_logic;
signal \N__38677\ : std_logic;
signal \N__38674\ : std_logic;
signal \N__38671\ : std_logic;
signal \N__38668\ : std_logic;
signal \N__38665\ : std_logic;
signal \N__38662\ : std_logic;
signal \N__38659\ : std_logic;
signal \N__38656\ : std_logic;
signal \N__38651\ : std_logic;
signal \N__38642\ : std_logic;
signal \N__38639\ : std_logic;
signal \N__38636\ : std_logic;
signal \N__38633\ : std_logic;
signal \N__38630\ : std_logic;
signal \N__38627\ : std_logic;
signal \N__38624\ : std_logic;
signal \N__38621\ : std_logic;
signal \N__38620\ : std_logic;
signal \N__38617\ : std_logic;
signal \N__38614\ : std_logic;
signal \N__38613\ : std_logic;
signal \N__38610\ : std_logic;
signal \N__38607\ : std_logic;
signal \N__38604\ : std_logic;
signal \N__38597\ : std_logic;
signal \N__38594\ : std_logic;
signal \N__38591\ : std_logic;
signal \N__38590\ : std_logic;
signal \N__38587\ : std_logic;
signal \N__38584\ : std_logic;
signal \N__38579\ : std_logic;
signal \N__38576\ : std_logic;
signal \N__38573\ : std_logic;
signal \N__38570\ : std_logic;
signal \N__38567\ : std_logic;
signal \N__38566\ : std_logic;
signal \N__38563\ : std_logic;
signal \N__38560\ : std_logic;
signal \N__38555\ : std_logic;
signal \N__38552\ : std_logic;
signal \N__38549\ : std_logic;
signal \N__38548\ : std_logic;
signal \N__38545\ : std_logic;
signal \N__38542\ : std_logic;
signal \N__38539\ : std_logic;
signal \N__38534\ : std_logic;
signal \N__38531\ : std_logic;
signal \N__38528\ : std_logic;
signal \N__38527\ : std_logic;
signal \N__38524\ : std_logic;
signal \N__38521\ : std_logic;
signal \N__38518\ : std_logic;
signal \N__38513\ : std_logic;
signal \N__38510\ : std_logic;
signal \N__38507\ : std_logic;
signal \N__38506\ : std_logic;
signal \N__38503\ : std_logic;
signal \N__38500\ : std_logic;
signal \N__38497\ : std_logic;
signal \N__38492\ : std_logic;
signal \N__38489\ : std_logic;
signal \N__38486\ : std_logic;
signal \N__38485\ : std_logic;
signal \N__38482\ : std_logic;
signal \N__38479\ : std_logic;
signal \N__38476\ : std_logic;
signal \N__38471\ : std_logic;
signal \N__38468\ : std_logic;
signal \N__38465\ : std_logic;
signal \N__38464\ : std_logic;
signal \N__38461\ : std_logic;
signal \N__38458\ : std_logic;
signal \N__38455\ : std_logic;
signal \N__38450\ : std_logic;
signal \N__38447\ : std_logic;
signal \N__38444\ : std_logic;
signal \N__38443\ : std_logic;
signal \N__38440\ : std_logic;
signal \N__38437\ : std_logic;
signal \N__38434\ : std_logic;
signal \N__38429\ : std_logic;
signal \N__38426\ : std_logic;
signal \N__38423\ : std_logic;
signal \N__38420\ : std_logic;
signal \N__38417\ : std_logic;
signal \N__38414\ : std_logic;
signal \N__38411\ : std_logic;
signal \N__38408\ : std_logic;
signal \N__38407\ : std_logic;
signal \N__38404\ : std_logic;
signal \N__38401\ : std_logic;
signal \N__38398\ : std_logic;
signal \N__38395\ : std_logic;
signal \N__38392\ : std_logic;
signal \N__38387\ : std_logic;
signal \N__38384\ : std_logic;
signal \N__38381\ : std_logic;
signal \N__38378\ : std_logic;
signal \N__38377\ : std_logic;
signal \N__38374\ : std_logic;
signal \N__38371\ : std_logic;
signal \N__38366\ : std_logic;
signal \N__38363\ : std_logic;
signal \N__38360\ : std_logic;
signal \N__38357\ : std_logic;
signal \N__38354\ : std_logic;
signal \N__38353\ : std_logic;
signal \N__38350\ : std_logic;
signal \N__38347\ : std_logic;
signal \N__38342\ : std_logic;
signal \N__38339\ : std_logic;
signal \N__38336\ : std_logic;
signal \N__38333\ : std_logic;
signal \N__38332\ : std_logic;
signal \N__38329\ : std_logic;
signal \N__38326\ : std_logic;
signal \N__38321\ : std_logic;
signal \N__38318\ : std_logic;
signal \N__38315\ : std_logic;
signal \N__38312\ : std_logic;
signal \N__38311\ : std_logic;
signal \N__38308\ : std_logic;
signal \N__38305\ : std_logic;
signal \N__38300\ : std_logic;
signal \N__38297\ : std_logic;
signal \N__38294\ : std_logic;
signal \N__38291\ : std_logic;
signal \N__38288\ : std_logic;
signal \N__38287\ : std_logic;
signal \N__38284\ : std_logic;
signal \N__38281\ : std_logic;
signal \N__38276\ : std_logic;
signal \N__38273\ : std_logic;
signal \N__38270\ : std_logic;
signal \N__38269\ : std_logic;
signal \N__38266\ : std_logic;
signal \N__38263\ : std_logic;
signal \N__38260\ : std_logic;
signal \N__38255\ : std_logic;
signal \N__38252\ : std_logic;
signal \N__38249\ : std_logic;
signal \N__38246\ : std_logic;
signal \N__38243\ : std_logic;
signal \N__38240\ : std_logic;
signal \N__38239\ : std_logic;
signal \N__38236\ : std_logic;
signal \N__38233\ : std_logic;
signal \N__38230\ : std_logic;
signal \N__38225\ : std_logic;
signal \N__38222\ : std_logic;
signal \N__38219\ : std_logic;
signal \N__38218\ : std_logic;
signal \N__38215\ : std_logic;
signal \N__38212\ : std_logic;
signal \N__38209\ : std_logic;
signal \N__38204\ : std_logic;
signal \N__38201\ : std_logic;
signal \N__38198\ : std_logic;
signal \N__38195\ : std_logic;
signal \N__38192\ : std_logic;
signal \N__38191\ : std_logic;
signal \N__38190\ : std_logic;
signal \N__38189\ : std_logic;
signal \N__38186\ : std_logic;
signal \N__38183\ : std_logic;
signal \N__38180\ : std_logic;
signal \N__38177\ : std_logic;
signal \N__38170\ : std_logic;
signal \N__38167\ : std_logic;
signal \N__38164\ : std_logic;
signal \N__38159\ : std_logic;
signal \N__38156\ : std_logic;
signal \N__38153\ : std_logic;
signal \N__38150\ : std_logic;
signal \N__38147\ : std_logic;
signal \N__38144\ : std_logic;
signal \N__38141\ : std_logic;
signal \N__38138\ : std_logic;
signal \N__38135\ : std_logic;
signal \N__38132\ : std_logic;
signal \N__38131\ : std_logic;
signal \N__38130\ : std_logic;
signal \N__38129\ : std_logic;
signal \N__38126\ : std_logic;
signal \N__38125\ : std_logic;
signal \N__38124\ : std_logic;
signal \N__38123\ : std_logic;
signal \N__38122\ : std_logic;
signal \N__38121\ : std_logic;
signal \N__38120\ : std_logic;
signal \N__38119\ : std_logic;
signal \N__38118\ : std_logic;
signal \N__38117\ : std_logic;
signal \N__38116\ : std_logic;
signal \N__38115\ : std_logic;
signal \N__38114\ : std_logic;
signal \N__38113\ : std_logic;
signal \N__38110\ : std_logic;
signal \N__38107\ : std_logic;
signal \N__38106\ : std_logic;
signal \N__38105\ : std_logic;
signal \N__38104\ : std_logic;
signal \N__38089\ : std_logic;
signal \N__38072\ : std_logic;
signal \N__38063\ : std_logic;
signal \N__38062\ : std_logic;
signal \N__38059\ : std_logic;
signal \N__38058\ : std_logic;
signal \N__38055\ : std_logic;
signal \N__38052\ : std_logic;
signal \N__38049\ : std_logic;
signal \N__38048\ : std_logic;
signal \N__38047\ : std_logic;
signal \N__38042\ : std_logic;
signal \N__38039\ : std_logic;
signal \N__38034\ : std_logic;
signal \N__38031\ : std_logic;
signal \N__38026\ : std_logic;
signal \N__38015\ : std_logic;
signal \N__38014\ : std_logic;
signal \N__38013\ : std_logic;
signal \N__38012\ : std_logic;
signal \N__38011\ : std_logic;
signal \N__38010\ : std_logic;
signal \N__38009\ : std_logic;
signal \N__38008\ : std_logic;
signal \N__38007\ : std_logic;
signal \N__38004\ : std_logic;
signal \N__38001\ : std_logic;
signal \N__37998\ : std_logic;
signal \N__37995\ : std_logic;
signal \N__37994\ : std_logic;
signal \N__37993\ : std_logic;
signal \N__37992\ : std_logic;
signal \N__37991\ : std_logic;
signal \N__37988\ : std_logic;
signal \N__37985\ : std_logic;
signal \N__37982\ : std_logic;
signal \N__37981\ : std_logic;
signal \N__37980\ : std_logic;
signal \N__37979\ : std_logic;
signal \N__37978\ : std_logic;
signal \N__37975\ : std_logic;
signal \N__37974\ : std_logic;
signal \N__37973\ : std_logic;
signal \N__37972\ : std_logic;
signal \N__37969\ : std_logic;
signal \N__37952\ : std_logic;
signal \N__37939\ : std_logic;
signal \N__37938\ : std_logic;
signal \N__37935\ : std_logic;
signal \N__37934\ : std_logic;
signal \N__37933\ : std_logic;
signal \N__37928\ : std_logic;
signal \N__37925\ : std_logic;
signal \N__37922\ : std_logic;
signal \N__37921\ : std_logic;
signal \N__37914\ : std_logic;
signal \N__37905\ : std_logic;
signal \N__37900\ : std_logic;
signal \N__37897\ : std_logic;
signal \N__37894\ : std_logic;
signal \N__37891\ : std_logic;
signal \N__37888\ : std_logic;
signal \N__37885\ : std_logic;
signal \N__37874\ : std_logic;
signal \N__37873\ : std_logic;
signal \N__37872\ : std_logic;
signal \N__37871\ : std_logic;
signal \N__37870\ : std_logic;
signal \N__37869\ : std_logic;
signal \N__37866\ : std_logic;
signal \N__37863\ : std_logic;
signal \N__37862\ : std_logic;
signal \N__37861\ : std_logic;
signal \N__37860\ : std_logic;
signal \N__37859\ : std_logic;
signal \N__37858\ : std_logic;
signal \N__37855\ : std_logic;
signal \N__37852\ : std_logic;
signal \N__37849\ : std_logic;
signal \N__37846\ : std_logic;
signal \N__37845\ : std_logic;
signal \N__37844\ : std_logic;
signal \N__37843\ : std_logic;
signal \N__37842\ : std_logic;
signal \N__37841\ : std_logic;
signal \N__37840\ : std_logic;
signal \N__37839\ : std_logic;
signal \N__37838\ : std_logic;
signal \N__37833\ : std_logic;
signal \N__37822\ : std_logic;
signal \N__37813\ : std_logic;
signal \N__37804\ : std_logic;
signal \N__37799\ : std_logic;
signal \N__37794\ : std_logic;
signal \N__37793\ : std_logic;
signal \N__37792\ : std_logic;
signal \N__37791\ : std_logic;
signal \N__37786\ : std_logic;
signal \N__37781\ : std_logic;
signal \N__37780\ : std_logic;
signal \N__37775\ : std_logic;
signal \N__37774\ : std_logic;
signal \N__37769\ : std_logic;
signal \N__37766\ : std_logic;
signal \N__37761\ : std_logic;
signal \N__37758\ : std_logic;
signal \N__37755\ : std_logic;
signal \N__37752\ : std_logic;
signal \N__37739\ : std_logic;
signal \N__37736\ : std_logic;
signal \N__37733\ : std_logic;
signal \N__37730\ : std_logic;
signal \N__37729\ : std_logic;
signal \N__37726\ : std_logic;
signal \N__37725\ : std_logic;
signal \N__37722\ : std_logic;
signal \N__37719\ : std_logic;
signal \N__37716\ : std_logic;
signal \N__37709\ : std_logic;
signal \N__37706\ : std_logic;
signal \N__37703\ : std_logic;
signal \N__37700\ : std_logic;
signal \N__37697\ : std_logic;
signal \N__37694\ : std_logic;
signal \N__37691\ : std_logic;
signal \N__37688\ : std_logic;
signal \N__37685\ : std_logic;
signal \N__37682\ : std_logic;
signal \N__37679\ : std_logic;
signal \N__37676\ : std_logic;
signal \N__37673\ : std_logic;
signal \N__37670\ : std_logic;
signal \N__37667\ : std_logic;
signal \N__37664\ : std_logic;
signal \N__37661\ : std_logic;
signal \N__37658\ : std_logic;
signal \N__37655\ : std_logic;
signal \N__37652\ : std_logic;
signal \N__37649\ : std_logic;
signal \N__37646\ : std_logic;
signal \N__37643\ : std_logic;
signal \N__37640\ : std_logic;
signal \N__37637\ : std_logic;
signal \N__37634\ : std_logic;
signal \N__37631\ : std_logic;
signal \N__37628\ : std_logic;
signal \N__37625\ : std_logic;
signal \N__37622\ : std_logic;
signal \N__37619\ : std_logic;
signal \N__37616\ : std_logic;
signal \N__37613\ : std_logic;
signal \N__37610\ : std_logic;
signal \N__37607\ : std_logic;
signal \N__37604\ : std_logic;
signal \N__37601\ : std_logic;
signal \N__37598\ : std_logic;
signal \N__37595\ : std_logic;
signal \N__37592\ : std_logic;
signal \N__37589\ : std_logic;
signal \N__37586\ : std_logic;
signal \N__37583\ : std_logic;
signal \N__37580\ : std_logic;
signal \N__37577\ : std_logic;
signal \N__37574\ : std_logic;
signal \N__37571\ : std_logic;
signal \N__37568\ : std_logic;
signal \N__37565\ : std_logic;
signal \N__37562\ : std_logic;
signal \N__37559\ : std_logic;
signal \N__37556\ : std_logic;
signal \N__37553\ : std_logic;
signal \N__37550\ : std_logic;
signal \N__37547\ : std_logic;
signal \N__37544\ : std_logic;
signal \N__37541\ : std_logic;
signal \N__37538\ : std_logic;
signal \N__37535\ : std_logic;
signal \N__37532\ : std_logic;
signal \N__37529\ : std_logic;
signal \N__37526\ : std_logic;
signal \N__37523\ : std_logic;
signal \N__37520\ : std_logic;
signal \N__37517\ : std_logic;
signal \N__37514\ : std_logic;
signal \N__37511\ : std_logic;
signal \N__37508\ : std_logic;
signal \N__37505\ : std_logic;
signal \N__37502\ : std_logic;
signal \N__37499\ : std_logic;
signal \N__37496\ : std_logic;
signal \N__37493\ : std_logic;
signal \N__37490\ : std_logic;
signal \N__37487\ : std_logic;
signal \N__37484\ : std_logic;
signal \N__37481\ : std_logic;
signal \N__37478\ : std_logic;
signal \N__37475\ : std_logic;
signal \N__37472\ : std_logic;
signal \N__37469\ : std_logic;
signal \N__37466\ : std_logic;
signal \N__37463\ : std_logic;
signal \N__37460\ : std_logic;
signal \N__37457\ : std_logic;
signal \N__37454\ : std_logic;
signal \N__37451\ : std_logic;
signal \N__37448\ : std_logic;
signal \N__37445\ : std_logic;
signal \N__37442\ : std_logic;
signal \N__37439\ : std_logic;
signal \N__37436\ : std_logic;
signal \N__37433\ : std_logic;
signal \N__37430\ : std_logic;
signal \N__37427\ : std_logic;
signal \N__37424\ : std_logic;
signal \N__37421\ : std_logic;
signal \N__37418\ : std_logic;
signal \N__37415\ : std_logic;
signal \N__37412\ : std_logic;
signal \N__37409\ : std_logic;
signal \N__37406\ : std_logic;
signal \N__37403\ : std_logic;
signal \N__37400\ : std_logic;
signal \N__37397\ : std_logic;
signal \N__37394\ : std_logic;
signal \N__37391\ : std_logic;
signal \N__37388\ : std_logic;
signal \N__37385\ : std_logic;
signal \N__37382\ : std_logic;
signal \N__37379\ : std_logic;
signal \N__37376\ : std_logic;
signal \N__37373\ : std_logic;
signal \N__37372\ : std_logic;
signal \N__37369\ : std_logic;
signal \N__37366\ : std_logic;
signal \N__37363\ : std_logic;
signal \N__37358\ : std_logic;
signal \N__37355\ : std_logic;
signal \N__37352\ : std_logic;
signal \N__37349\ : std_logic;
signal \N__37346\ : std_logic;
signal \N__37345\ : std_logic;
signal \N__37342\ : std_logic;
signal \N__37339\ : std_logic;
signal \N__37336\ : std_logic;
signal \N__37331\ : std_logic;
signal \N__37328\ : std_logic;
signal \N__37325\ : std_logic;
signal \N__37322\ : std_logic;
signal \N__37321\ : std_logic;
signal \N__37318\ : std_logic;
signal \N__37315\ : std_logic;
signal \N__37310\ : std_logic;
signal \N__37307\ : std_logic;
signal \N__37304\ : std_logic;
signal \N__37301\ : std_logic;
signal \N__37298\ : std_logic;
signal \N__37295\ : std_logic;
signal \N__37292\ : std_logic;
signal \N__37289\ : std_logic;
signal \N__37286\ : std_logic;
signal \N__37283\ : std_logic;
signal \N__37280\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37274\ : std_logic;
signal \N__37271\ : std_logic;
signal \N__37268\ : std_logic;
signal \N__37265\ : std_logic;
signal \N__37262\ : std_logic;
signal \N__37259\ : std_logic;
signal \N__37256\ : std_logic;
signal \N__37253\ : std_logic;
signal \N__37250\ : std_logic;
signal \N__37247\ : std_logic;
signal \N__37244\ : std_logic;
signal \N__37241\ : std_logic;
signal \N__37238\ : std_logic;
signal \N__37235\ : std_logic;
signal \N__37232\ : std_logic;
signal \N__37231\ : std_logic;
signal \N__37228\ : std_logic;
signal \N__37225\ : std_logic;
signal \N__37220\ : std_logic;
signal \N__37217\ : std_logic;
signal \N__37214\ : std_logic;
signal \N__37211\ : std_logic;
signal \N__37208\ : std_logic;
signal \N__37205\ : std_logic;
signal \N__37204\ : std_logic;
signal \N__37201\ : std_logic;
signal \N__37198\ : std_logic;
signal \N__37193\ : std_logic;
signal \N__37190\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37184\ : std_logic;
signal \N__37181\ : std_logic;
signal \N__37178\ : std_logic;
signal \N__37177\ : std_logic;
signal \N__37174\ : std_logic;
signal \N__37171\ : std_logic;
signal \N__37166\ : std_logic;
signal \N__37163\ : std_logic;
signal \N__37160\ : std_logic;
signal \N__37157\ : std_logic;
signal \N__37154\ : std_logic;
signal \N__37151\ : std_logic;
signal \N__37148\ : std_logic;
signal \N__37147\ : std_logic;
signal \N__37144\ : std_logic;
signal \N__37141\ : std_logic;
signal \N__37136\ : std_logic;
signal \N__37133\ : std_logic;
signal \N__37130\ : std_logic;
signal \N__37127\ : std_logic;
signal \N__37124\ : std_logic;
signal \N__37121\ : std_logic;
signal \N__37120\ : std_logic;
signal \N__37117\ : std_logic;
signal \N__37114\ : std_logic;
signal \N__37109\ : std_logic;
signal \N__37106\ : std_logic;
signal \N__37103\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37097\ : std_logic;
signal \N__37096\ : std_logic;
signal \N__37093\ : std_logic;
signal \N__37090\ : std_logic;
signal \N__37085\ : std_logic;
signal \N__37082\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37076\ : std_logic;
signal \N__37075\ : std_logic;
signal \N__37072\ : std_logic;
signal \N__37069\ : std_logic;
signal \N__37064\ : std_logic;
signal \N__37061\ : std_logic;
signal \N__37058\ : std_logic;
signal \N__37057\ : std_logic;
signal \N__37054\ : std_logic;
signal \N__37051\ : std_logic;
signal \N__37048\ : std_logic;
signal \N__37043\ : std_logic;
signal \N__37040\ : std_logic;
signal \N__37037\ : std_logic;
signal \N__37034\ : std_logic;
signal \N__37031\ : std_logic;
signal \N__37030\ : std_logic;
signal \N__37027\ : std_logic;
signal \N__37026\ : std_logic;
signal \N__37023\ : std_logic;
signal \N__37020\ : std_logic;
signal \N__37017\ : std_logic;
signal \N__37010\ : std_logic;
signal \N__37009\ : std_logic;
signal \N__37006\ : std_logic;
signal \N__37003\ : std_logic;
signal \N__36998\ : std_logic;
signal \N__36995\ : std_logic;
signal \N__36992\ : std_logic;
signal \N__36989\ : std_logic;
signal \N__36986\ : std_logic;
signal \N__36983\ : std_logic;
signal \N__36980\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36974\ : std_logic;
signal \N__36971\ : std_logic;
signal \N__36968\ : std_logic;
signal \N__36965\ : std_logic;
signal \N__36964\ : std_logic;
signal \N__36961\ : std_logic;
signal \N__36958\ : std_logic;
signal \N__36953\ : std_logic;
signal \N__36950\ : std_logic;
signal \N__36947\ : std_logic;
signal \N__36944\ : std_logic;
signal \N__36941\ : std_logic;
signal \N__36938\ : std_logic;
signal \N__36937\ : std_logic;
signal \N__36934\ : std_logic;
signal \N__36931\ : std_logic;
signal \N__36926\ : std_logic;
signal \N__36923\ : std_logic;
signal \N__36920\ : std_logic;
signal \N__36917\ : std_logic;
signal \N__36914\ : std_logic;
signal \N__36911\ : std_logic;
signal \N__36908\ : std_logic;
signal \N__36905\ : std_logic;
signal \N__36902\ : std_logic;
signal \N__36901\ : std_logic;
signal \N__36898\ : std_logic;
signal \N__36895\ : std_logic;
signal \N__36890\ : std_logic;
signal \N__36887\ : std_logic;
signal \N__36884\ : std_logic;
signal \N__36881\ : std_logic;
signal \N__36878\ : std_logic;
signal \N__36875\ : std_logic;
signal \N__36874\ : std_logic;
signal \N__36871\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36863\ : std_logic;
signal \N__36860\ : std_logic;
signal \N__36857\ : std_logic;
signal \N__36854\ : std_logic;
signal \N__36851\ : std_logic;
signal \N__36848\ : std_logic;
signal \N__36845\ : std_logic;
signal \N__36842\ : std_logic;
signal \N__36839\ : std_logic;
signal \N__36836\ : std_logic;
signal \N__36833\ : std_logic;
signal \N__36830\ : std_logic;
signal \N__36827\ : std_logic;
signal \N__36824\ : std_logic;
signal \N__36823\ : std_logic;
signal \N__36820\ : std_logic;
signal \N__36819\ : std_logic;
signal \N__36816\ : std_logic;
signal \N__36813\ : std_logic;
signal \N__36810\ : std_logic;
signal \N__36805\ : std_logic;
signal \N__36800\ : std_logic;
signal \N__36799\ : std_logic;
signal \N__36796\ : std_logic;
signal \N__36793\ : std_logic;
signal \N__36792\ : std_logic;
signal \N__36789\ : std_logic;
signal \N__36786\ : std_logic;
signal \N__36783\ : std_logic;
signal \N__36780\ : std_logic;
signal \N__36777\ : std_logic;
signal \N__36774\ : std_logic;
signal \N__36767\ : std_logic;
signal \N__36764\ : std_logic;
signal \N__36763\ : std_logic;
signal \N__36762\ : std_logic;
signal \N__36759\ : std_logic;
signal \N__36754\ : std_logic;
signal \N__36751\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36743\ : std_logic;
signal \N__36742\ : std_logic;
signal \N__36741\ : std_logic;
signal \N__36738\ : std_logic;
signal \N__36733\ : std_logic;
signal \N__36728\ : std_logic;
signal \N__36725\ : std_logic;
signal \N__36724\ : std_logic;
signal \N__36723\ : std_logic;
signal \N__36720\ : std_logic;
signal \N__36717\ : std_logic;
signal \N__36714\ : std_logic;
signal \N__36709\ : std_logic;
signal \N__36704\ : std_logic;
signal \N__36701\ : std_logic;
signal \N__36700\ : std_logic;
signal \N__36699\ : std_logic;
signal \N__36698\ : std_logic;
signal \N__36697\ : std_logic;
signal \N__36696\ : std_logic;
signal \N__36693\ : std_logic;
signal \N__36686\ : std_logic;
signal \N__36681\ : std_logic;
signal \N__36676\ : std_logic;
signal \N__36673\ : std_logic;
signal \N__36670\ : std_logic;
signal \N__36667\ : std_logic;
signal \N__36664\ : std_logic;
signal \N__36661\ : std_logic;
signal \N__36658\ : std_logic;
signal \N__36655\ : std_logic;
signal \N__36650\ : std_logic;
signal \N__36647\ : std_logic;
signal \N__36646\ : std_logic;
signal \N__36645\ : std_logic;
signal \N__36642\ : std_logic;
signal \N__36637\ : std_logic;
signal \N__36634\ : std_logic;
signal \N__36629\ : std_logic;
signal \N__36626\ : std_logic;
signal \N__36623\ : std_logic;
signal \N__36620\ : std_logic;
signal \N__36617\ : std_logic;
signal \N__36614\ : std_logic;
signal \N__36611\ : std_logic;
signal \N__36608\ : std_logic;
signal \N__36605\ : std_logic;
signal \N__36602\ : std_logic;
signal \N__36599\ : std_logic;
signal \N__36598\ : std_logic;
signal \N__36597\ : std_logic;
signal \N__36596\ : std_logic;
signal \N__36593\ : std_logic;
signal \N__36590\ : std_logic;
signal \N__36585\ : std_logic;
signal \N__36582\ : std_logic;
signal \N__36575\ : std_logic;
signal \N__36574\ : std_logic;
signal \N__36573\ : std_logic;
signal \N__36570\ : std_logic;
signal \N__36567\ : std_logic;
signal \N__36564\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36554\ : std_logic;
signal \N__36553\ : std_logic;
signal \N__36552\ : std_logic;
signal \N__36549\ : std_logic;
signal \N__36546\ : std_logic;
signal \N__36543\ : std_logic;
signal \N__36536\ : std_logic;
signal \N__36535\ : std_logic;
signal \N__36534\ : std_logic;
signal \N__36531\ : std_logic;
signal \N__36526\ : std_logic;
signal \N__36525\ : std_logic;
signal \N__36520\ : std_logic;
signal \N__36517\ : std_logic;
signal \N__36512\ : std_logic;
signal \N__36509\ : std_logic;
signal \N__36508\ : std_logic;
signal \N__36507\ : std_logic;
signal \N__36504\ : std_logic;
signal \N__36501\ : std_logic;
signal \N__36498\ : std_logic;
signal \N__36491\ : std_logic;
signal \N__36490\ : std_logic;
signal \N__36489\ : std_logic;
signal \N__36486\ : std_logic;
signal \N__36483\ : std_logic;
signal \N__36480\ : std_logic;
signal \N__36473\ : std_logic;
signal \N__36470\ : std_logic;
signal \N__36467\ : std_logic;
signal \N__36464\ : std_logic;
signal \N__36461\ : std_logic;
signal \N__36458\ : std_logic;
signal \N__36455\ : std_logic;
signal \N__36452\ : std_logic;
signal \N__36451\ : std_logic;
signal \N__36448\ : std_logic;
signal \N__36445\ : std_logic;
signal \N__36442\ : std_logic;
signal \N__36441\ : std_logic;
signal \N__36440\ : std_logic;
signal \N__36437\ : std_logic;
signal \N__36434\ : std_logic;
signal \N__36431\ : std_logic;
signal \N__36428\ : std_logic;
signal \N__36419\ : std_logic;
signal \N__36418\ : std_logic;
signal \N__36417\ : std_logic;
signal \N__36414\ : std_logic;
signal \N__36413\ : std_logic;
signal \N__36410\ : std_logic;
signal \N__36407\ : std_logic;
signal \N__36404\ : std_logic;
signal \N__36403\ : std_logic;
signal \N__36400\ : std_logic;
signal \N__36397\ : std_logic;
signal \N__36394\ : std_logic;
signal \N__36391\ : std_logic;
signal \N__36388\ : std_logic;
signal \N__36385\ : std_logic;
signal \N__36382\ : std_logic;
signal \N__36379\ : std_logic;
signal \N__36374\ : std_logic;
signal \N__36365\ : std_logic;
signal \N__36364\ : std_logic;
signal \N__36361\ : std_logic;
signal \N__36358\ : std_logic;
signal \N__36353\ : std_logic;
signal \N__36350\ : std_logic;
signal \N__36347\ : std_logic;
signal \N__36344\ : std_logic;
signal \N__36341\ : std_logic;
signal \N__36338\ : std_logic;
signal \N__36335\ : std_logic;
signal \N__36332\ : std_logic;
signal \N__36329\ : std_logic;
signal \N__36326\ : std_logic;
signal \N__36325\ : std_logic;
signal \N__36324\ : std_logic;
signal \N__36323\ : std_logic;
signal \N__36322\ : std_logic;
signal \N__36321\ : std_logic;
signal \N__36320\ : std_logic;
signal \N__36319\ : std_logic;
signal \N__36318\ : std_logic;
signal \N__36317\ : std_logic;
signal \N__36316\ : std_logic;
signal \N__36315\ : std_logic;
signal \N__36312\ : std_logic;
signal \N__36295\ : std_logic;
signal \N__36294\ : std_logic;
signal \N__36293\ : std_logic;
signal \N__36292\ : std_logic;
signal \N__36291\ : std_logic;
signal \N__36290\ : std_logic;
signal \N__36289\ : std_logic;
signal \N__36288\ : std_logic;
signal \N__36287\ : std_logic;
signal \N__36280\ : std_logic;
signal \N__36279\ : std_logic;
signal \N__36278\ : std_logic;
signal \N__36273\ : std_logic;
signal \N__36256\ : std_logic;
signal \N__36255\ : std_logic;
signal \N__36252\ : std_logic;
signal \N__36249\ : std_logic;
signal \N__36246\ : std_logic;
signal \N__36245\ : std_logic;
signal \N__36240\ : std_logic;
signal \N__36237\ : std_logic;
signal \N__36232\ : std_logic;
signal \N__36229\ : std_logic;
signal \N__36226\ : std_logic;
signal \N__36223\ : std_logic;
signal \N__36216\ : std_logic;
signal \N__36209\ : std_logic;
signal \N__36208\ : std_logic;
signal \N__36207\ : std_logic;
signal \N__36206\ : std_logic;
signal \N__36205\ : std_logic;
signal \N__36204\ : std_logic;
signal \N__36201\ : std_logic;
signal \N__36198\ : std_logic;
signal \N__36197\ : std_logic;
signal \N__36194\ : std_logic;
signal \N__36193\ : std_logic;
signal \N__36192\ : std_logic;
signal \N__36191\ : std_logic;
signal \N__36188\ : std_logic;
signal \N__36185\ : std_logic;
signal \N__36184\ : std_logic;
signal \N__36183\ : std_logic;
signal \N__36182\ : std_logic;
signal \N__36181\ : std_logic;
signal \N__36180\ : std_logic;
signal \N__36177\ : std_logic;
signal \N__36176\ : std_logic;
signal \N__36173\ : std_logic;
signal \N__36156\ : std_logic;
signal \N__36155\ : std_logic;
signal \N__36152\ : std_logic;
signal \N__36149\ : std_logic;
signal \N__36148\ : std_logic;
signal \N__36145\ : std_logic;
signal \N__36144\ : std_logic;
signal \N__36143\ : std_logic;
signal \N__36140\ : std_logic;
signal \N__36137\ : std_logic;
signal \N__36134\ : std_logic;
signal \N__36131\ : std_logic;
signal \N__36126\ : std_logic;
signal \N__36109\ : std_logic;
signal \N__36106\ : std_logic;
signal \N__36105\ : std_logic;
signal \N__36104\ : std_logic;
signal \N__36103\ : std_logic;
signal \N__36102\ : std_logic;
signal \N__36099\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36091\ : std_logic;
signal \N__36088\ : std_logic;
signal \N__36081\ : std_logic;
signal \N__36078\ : std_logic;
signal \N__36065\ : std_logic;
signal \N__36064\ : std_logic;
signal \N__36063\ : std_logic;
signal \N__36062\ : std_logic;
signal \N__36061\ : std_logic;
signal \N__36060\ : std_logic;
signal \N__36057\ : std_logic;
signal \N__36056\ : std_logic;
signal \N__36055\ : std_logic;
signal \N__36054\ : std_logic;
signal \N__36053\ : std_logic;
signal \N__36052\ : std_logic;
signal \N__36051\ : std_logic;
signal \N__36050\ : std_logic;
signal \N__36047\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36038\ : std_logic;
signal \N__36037\ : std_logic;
signal \N__36036\ : std_logic;
signal \N__36035\ : std_logic;
signal \N__36034\ : std_logic;
signal \N__36031\ : std_logic;
signal \N__36028\ : std_logic;
signal \N__36025\ : std_logic;
signal \N__36022\ : std_logic;
signal \N__36021\ : std_logic;
signal \N__36018\ : std_logic;
signal \N__36017\ : std_logic;
signal \N__36016\ : std_logic;
signal \N__36013\ : std_logic;
signal \N__36010\ : std_logic;
signal \N__36007\ : std_logic;
signal \N__36004\ : std_logic;
signal \N__36003\ : std_logic;
signal \N__36002\ : std_logic;
signal \N__36001\ : std_logic;
signal \N__36000\ : std_logic;
signal \N__35991\ : std_logic;
signal \N__35982\ : std_logic;
signal \N__35979\ : std_logic;
signal \N__35976\ : std_logic;
signal \N__35969\ : std_logic;
signal \N__35966\ : std_logic;
signal \N__35963\ : std_logic;
signal \N__35960\ : std_logic;
signal \N__35951\ : std_logic;
signal \N__35942\ : std_logic;
signal \N__35933\ : std_logic;
signal \N__35930\ : std_logic;
signal \N__35925\ : std_logic;
signal \N__35912\ : std_logic;
signal \N__35909\ : std_logic;
signal \N__35906\ : std_logic;
signal \N__35903\ : std_logic;
signal \N__35900\ : std_logic;
signal \N__35897\ : std_logic;
signal \N__35894\ : std_logic;
signal \N__35891\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35887\ : std_logic;
signal \N__35884\ : std_logic;
signal \N__35881\ : std_logic;
signal \N__35880\ : std_logic;
signal \N__35879\ : std_logic;
signal \N__35874\ : std_logic;
signal \N__35871\ : std_logic;
signal \N__35868\ : std_logic;
signal \N__35865\ : std_logic;
signal \N__35862\ : std_logic;
signal \N__35861\ : std_logic;
signal \N__35858\ : std_logic;
signal \N__35855\ : std_logic;
signal \N__35852\ : std_logic;
signal \N__35849\ : std_logic;
signal \N__35846\ : std_logic;
signal \N__35841\ : std_logic;
signal \N__35838\ : std_logic;
signal \N__35837\ : std_logic;
signal \N__35836\ : std_logic;
signal \N__35833\ : std_logic;
signal \N__35828\ : std_logic;
signal \N__35825\ : std_logic;
signal \N__35822\ : std_logic;
signal \N__35813\ : std_logic;
signal \N__35810\ : std_logic;
signal \N__35807\ : std_logic;
signal \N__35804\ : std_logic;
signal \N__35801\ : std_logic;
signal \N__35798\ : std_logic;
signal \N__35795\ : std_logic;
signal \N__35792\ : std_logic;
signal \N__35789\ : std_logic;
signal \N__35786\ : std_logic;
signal \N__35783\ : std_logic;
signal \N__35780\ : std_logic;
signal \N__35777\ : std_logic;
signal \N__35774\ : std_logic;
signal \N__35771\ : std_logic;
signal \N__35768\ : std_logic;
signal \N__35765\ : std_logic;
signal \N__35762\ : std_logic;
signal \N__35759\ : std_logic;
signal \N__35756\ : std_logic;
signal \N__35753\ : std_logic;
signal \N__35750\ : std_logic;
signal \N__35747\ : std_logic;
signal \N__35744\ : std_logic;
signal \N__35741\ : std_logic;
signal \N__35738\ : std_logic;
signal \N__35735\ : std_logic;
signal \N__35732\ : std_logic;
signal \N__35729\ : std_logic;
signal \N__35726\ : std_logic;
signal \N__35723\ : std_logic;
signal \N__35720\ : std_logic;
signal \N__35717\ : std_logic;
signal \N__35714\ : std_logic;
signal \N__35711\ : std_logic;
signal \N__35708\ : std_logic;
signal \N__35705\ : std_logic;
signal \N__35702\ : std_logic;
signal \N__35699\ : std_logic;
signal \N__35696\ : std_logic;
signal \N__35693\ : std_logic;
signal \N__35690\ : std_logic;
signal \N__35687\ : std_logic;
signal \N__35684\ : std_logic;
signal \N__35681\ : std_logic;
signal \N__35678\ : std_logic;
signal \N__35675\ : std_logic;
signal \N__35672\ : std_logic;
signal \N__35669\ : std_logic;
signal \N__35666\ : std_logic;
signal \N__35663\ : std_logic;
signal \N__35660\ : std_logic;
signal \N__35657\ : std_logic;
signal \N__35654\ : std_logic;
signal \N__35651\ : std_logic;
signal \N__35648\ : std_logic;
signal \N__35645\ : std_logic;
signal \N__35642\ : std_logic;
signal \N__35639\ : std_logic;
signal \N__35636\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35630\ : std_logic;
signal \N__35627\ : std_logic;
signal \N__35624\ : std_logic;
signal \N__35621\ : std_logic;
signal \N__35618\ : std_logic;
signal \N__35617\ : std_logic;
signal \N__35616\ : std_logic;
signal \N__35615\ : std_logic;
signal \N__35612\ : std_logic;
signal \N__35611\ : std_logic;
signal \N__35610\ : std_logic;
signal \N__35605\ : std_logic;
signal \N__35604\ : std_logic;
signal \N__35601\ : std_logic;
signal \N__35600\ : std_logic;
signal \N__35599\ : std_logic;
signal \N__35598\ : std_logic;
signal \N__35597\ : std_logic;
signal \N__35596\ : std_logic;
signal \N__35595\ : std_logic;
signal \N__35594\ : std_logic;
signal \N__35587\ : std_logic;
signal \N__35586\ : std_logic;
signal \N__35585\ : std_logic;
signal \N__35584\ : std_logic;
signal \N__35583\ : std_logic;
signal \N__35580\ : std_logic;
signal \N__35577\ : std_logic;
signal \N__35568\ : std_logic;
signal \N__35559\ : std_logic;
signal \N__35556\ : std_logic;
signal \N__35547\ : std_logic;
signal \N__35544\ : std_logic;
signal \N__35543\ : std_logic;
signal \N__35542\ : std_logic;
signal \N__35541\ : std_logic;
signal \N__35540\ : std_logic;
signal \N__35537\ : std_logic;
signal \N__35528\ : std_logic;
signal \N__35525\ : std_logic;
signal \N__35516\ : std_logic;
signal \N__35513\ : std_logic;
signal \N__35508\ : std_logic;
signal \N__35501\ : std_logic;
signal \N__35500\ : std_logic;
signal \N__35499\ : std_logic;
signal \N__35496\ : std_logic;
signal \N__35493\ : std_logic;
signal \N__35490\ : std_logic;
signal \N__35489\ : std_logic;
signal \N__35488\ : std_logic;
signal \N__35485\ : std_logic;
signal \N__35482\ : std_logic;
signal \N__35479\ : std_logic;
signal \N__35476\ : std_logic;
signal \N__35473\ : std_logic;
signal \N__35470\ : std_logic;
signal \N__35467\ : std_logic;
signal \N__35462\ : std_logic;
signal \N__35453\ : std_logic;
signal \N__35452\ : std_logic;
signal \N__35451\ : std_logic;
signal \N__35450\ : std_logic;
signal \N__35449\ : std_logic;
signal \N__35448\ : std_logic;
signal \N__35447\ : std_logic;
signal \N__35440\ : std_logic;
signal \N__35439\ : std_logic;
signal \N__35438\ : std_logic;
signal \N__35437\ : std_logic;
signal \N__35436\ : std_logic;
signal \N__35427\ : std_logic;
signal \N__35424\ : std_logic;
signal \N__35415\ : std_logic;
signal \N__35414\ : std_logic;
signal \N__35413\ : std_logic;
signal \N__35412\ : std_logic;
signal \N__35409\ : std_logic;
signal \N__35404\ : std_logic;
signal \N__35397\ : std_logic;
signal \N__35390\ : std_logic;
signal \N__35387\ : std_logic;
signal \N__35384\ : std_logic;
signal \N__35381\ : std_logic;
signal \N__35378\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35372\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35368\ : std_logic;
signal \N__35365\ : std_logic;
signal \N__35364\ : std_logic;
signal \N__35361\ : std_logic;
signal \N__35360\ : std_logic;
signal \N__35357\ : std_logic;
signal \N__35354\ : std_logic;
signal \N__35351\ : std_logic;
signal \N__35350\ : std_logic;
signal \N__35347\ : std_logic;
signal \N__35342\ : std_logic;
signal \N__35339\ : std_logic;
signal \N__35336\ : std_logic;
signal \N__35333\ : std_logic;
signal \N__35330\ : std_logic;
signal \N__35327\ : std_logic;
signal \N__35324\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35312\ : std_logic;
signal \N__35311\ : std_logic;
signal \N__35308\ : std_logic;
signal \N__35305\ : std_logic;
signal \N__35304\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35298\ : std_logic;
signal \N__35295\ : std_logic;
signal \N__35292\ : std_logic;
signal \N__35289\ : std_logic;
signal \N__35286\ : std_logic;
signal \N__35279\ : std_logic;
signal \N__35278\ : std_logic;
signal \N__35275\ : std_logic;
signal \N__35274\ : std_logic;
signal \N__35271\ : std_logic;
signal \N__35268\ : std_logic;
signal \N__35267\ : std_logic;
signal \N__35264\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35258\ : std_logic;
signal \N__35253\ : std_logic;
signal \N__35252\ : std_logic;
signal \N__35249\ : std_logic;
signal \N__35244\ : std_logic;
signal \N__35241\ : std_logic;
signal \N__35238\ : std_logic;
signal \N__35235\ : std_logic;
signal \N__35228\ : std_logic;
signal \N__35225\ : std_logic;
signal \N__35222\ : std_logic;
signal \N__35221\ : std_logic;
signal \N__35218\ : std_logic;
signal \N__35215\ : std_logic;
signal \N__35214\ : std_logic;
signal \N__35213\ : std_logic;
signal \N__35210\ : std_logic;
signal \N__35207\ : std_logic;
signal \N__35202\ : std_logic;
signal \N__35195\ : std_logic;
signal \N__35194\ : std_logic;
signal \N__35191\ : std_logic;
signal \N__35188\ : std_logic;
signal \N__35187\ : std_logic;
signal \N__35184\ : std_logic;
signal \N__35181\ : std_logic;
signal \N__35180\ : std_logic;
signal \N__35177\ : std_logic;
signal \N__35176\ : std_logic;
signal \N__35173\ : std_logic;
signal \N__35170\ : std_logic;
signal \N__35167\ : std_logic;
signal \N__35164\ : std_logic;
signal \N__35161\ : std_logic;
signal \N__35158\ : std_logic;
signal \N__35151\ : std_logic;
signal \N__35144\ : std_logic;
signal \N__35143\ : std_logic;
signal \N__35140\ : std_logic;
signal \N__35137\ : std_logic;
signal \N__35136\ : std_logic;
signal \N__35133\ : std_logic;
signal \N__35132\ : std_logic;
signal \N__35131\ : std_logic;
signal \N__35128\ : std_logic;
signal \N__35125\ : std_logic;
signal \N__35122\ : std_logic;
signal \N__35119\ : std_logic;
signal \N__35116\ : std_logic;
signal \N__35113\ : std_logic;
signal \N__35110\ : std_logic;
signal \N__35105\ : std_logic;
signal \N__35096\ : std_logic;
signal \N__35095\ : std_logic;
signal \N__35092\ : std_logic;
signal \N__35091\ : std_logic;
signal \N__35090\ : std_logic;
signal \N__35089\ : std_logic;
signal \N__35086\ : std_logic;
signal \N__35083\ : std_logic;
signal \N__35080\ : std_logic;
signal \N__35075\ : std_logic;
signal \N__35072\ : std_logic;
signal \N__35067\ : std_logic;
signal \N__35064\ : std_logic;
signal \N__35057\ : std_logic;
signal \N__35056\ : std_logic;
signal \N__35053\ : std_logic;
signal \N__35050\ : std_logic;
signal \N__35047\ : std_logic;
signal \N__35046\ : std_logic;
signal \N__35045\ : std_logic;
signal \N__35040\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35036\ : std_logic;
signal \N__35033\ : std_logic;
signal \N__35030\ : std_logic;
signal \N__35027\ : std_logic;
signal \N__35024\ : std_logic;
signal \N__35015\ : std_logic;
signal \N__35014\ : std_logic;
signal \N__35013\ : std_logic;
signal \N__35012\ : std_logic;
signal \N__35011\ : std_logic;
signal \N__35010\ : std_logic;
signal \N__35009\ : std_logic;
signal \N__35002\ : std_logic;
signal \N__34993\ : std_logic;
signal \N__34992\ : std_logic;
signal \N__34991\ : std_logic;
signal \N__34990\ : std_logic;
signal \N__34989\ : std_logic;
signal \N__34988\ : std_logic;
signal \N__34987\ : std_logic;
signal \N__34986\ : std_logic;
signal \N__34985\ : std_logic;
signal \N__34982\ : std_logic;
signal \N__34979\ : std_logic;
signal \N__34976\ : std_logic;
signal \N__34969\ : std_logic;
signal \N__34964\ : std_logic;
signal \N__34963\ : std_logic;
signal \N__34958\ : std_logic;
signal \N__34955\ : std_logic;
signal \N__34950\ : std_logic;
signal \N__34949\ : std_logic;
signal \N__34948\ : std_logic;
signal \N__34945\ : std_logic;
signal \N__34942\ : std_logic;
signal \N__34939\ : std_logic;
signal \N__34936\ : std_logic;
signal \N__34933\ : std_logic;
signal \N__34930\ : std_logic;
signal \N__34925\ : std_logic;
signal \N__34922\ : std_logic;
signal \N__34915\ : std_logic;
signal \N__34904\ : std_logic;
signal \N__34903\ : std_logic;
signal \N__34900\ : std_logic;
signal \N__34897\ : std_logic;
signal \N__34894\ : std_logic;
signal \N__34893\ : std_logic;
signal \N__34888\ : std_logic;
signal \N__34885\ : std_logic;
signal \N__34880\ : std_logic;
signal \N__34877\ : std_logic;
signal \N__34874\ : std_logic;
signal \N__34873\ : std_logic;
signal \N__34870\ : std_logic;
signal \N__34867\ : std_logic;
signal \N__34864\ : std_logic;
signal \N__34861\ : std_logic;
signal \N__34856\ : std_logic;
signal \N__34853\ : std_logic;
signal \N__34850\ : std_logic;
signal \N__34847\ : std_logic;
signal \N__34844\ : std_logic;
signal \N__34843\ : std_logic;
signal \N__34840\ : std_logic;
signal \N__34837\ : std_logic;
signal \N__34834\ : std_logic;
signal \N__34831\ : std_logic;
signal \N__34828\ : std_logic;
signal \N__34823\ : std_logic;
signal \N__34820\ : std_logic;
signal \N__34817\ : std_logic;
signal \N__34816\ : std_logic;
signal \N__34813\ : std_logic;
signal \N__34810\ : std_logic;
signal \N__34809\ : std_logic;
signal \N__34808\ : std_logic;
signal \N__34807\ : std_logic;
signal \N__34804\ : std_logic;
signal \N__34801\ : std_logic;
signal \N__34796\ : std_logic;
signal \N__34793\ : std_logic;
signal \N__34786\ : std_logic;
signal \N__34783\ : std_logic;
signal \N__34780\ : std_logic;
signal \N__34775\ : std_logic;
signal \N__34772\ : std_logic;
signal \N__34771\ : std_logic;
signal \N__34770\ : std_logic;
signal \N__34769\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34765\ : std_logic;
signal \N__34758\ : std_logic;
signal \N__34755\ : std_logic;
signal \N__34752\ : std_logic;
signal \N__34749\ : std_logic;
signal \N__34742\ : std_logic;
signal \N__34741\ : std_logic;
signal \N__34738\ : std_logic;
signal \N__34737\ : std_logic;
signal \N__34736\ : std_logic;
signal \N__34733\ : std_logic;
signal \N__34732\ : std_logic;
signal \N__34729\ : std_logic;
signal \N__34726\ : std_logic;
signal \N__34721\ : std_logic;
signal \N__34718\ : std_logic;
signal \N__34715\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34709\ : std_logic;
signal \N__34706\ : std_logic;
signal \N__34703\ : std_logic;
signal \N__34698\ : std_logic;
signal \N__34691\ : std_logic;
signal \N__34688\ : std_logic;
signal \N__34685\ : std_logic;
signal \N__34682\ : std_logic;
signal \N__34681\ : std_logic;
signal \N__34680\ : std_logic;
signal \N__34677\ : std_logic;
signal \N__34674\ : std_logic;
signal \N__34673\ : std_logic;
signal \N__34672\ : std_logic;
signal \N__34669\ : std_logic;
signal \N__34664\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34658\ : std_logic;
signal \N__34649\ : std_logic;
signal \N__34648\ : std_logic;
signal \N__34645\ : std_logic;
signal \N__34642\ : std_logic;
signal \N__34641\ : std_logic;
signal \N__34640\ : std_logic;
signal \N__34637\ : std_logic;
signal \N__34636\ : std_logic;
signal \N__34633\ : std_logic;
signal \N__34630\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34624\ : std_logic;
signal \N__34621\ : std_logic;
signal \N__34616\ : std_logic;
signal \N__34607\ : std_logic;
signal \N__34606\ : std_logic;
signal \N__34603\ : std_logic;
signal \N__34600\ : std_logic;
signal \N__34597\ : std_logic;
signal \N__34596\ : std_logic;
signal \N__34595\ : std_logic;
signal \N__34592\ : std_logic;
signal \N__34589\ : std_logic;
signal \N__34586\ : std_logic;
signal \N__34583\ : std_logic;
signal \N__34578\ : std_logic;
signal \N__34575\ : std_logic;
signal \N__34572\ : std_logic;
signal \N__34565\ : std_logic;
signal \N__34562\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34557\ : std_logic;
signal \N__34556\ : std_logic;
signal \N__34553\ : std_logic;
signal \N__34550\ : std_logic;
signal \N__34547\ : std_logic;
signal \N__34544\ : std_logic;
signal \N__34543\ : std_logic;
signal \N__34540\ : std_logic;
signal \N__34533\ : std_logic;
signal \N__34530\ : std_logic;
signal \N__34527\ : std_logic;
signal \N__34524\ : std_logic;
signal \N__34517\ : std_logic;
signal \N__34514\ : std_logic;
signal \N__34513\ : std_logic;
signal \N__34512\ : std_logic;
signal \N__34511\ : std_logic;
signal \N__34508\ : std_logic;
signal \N__34505\ : std_logic;
signal \N__34502\ : std_logic;
signal \N__34499\ : std_logic;
signal \N__34492\ : std_logic;
signal \N__34487\ : std_logic;
signal \N__34486\ : std_logic;
signal \N__34483\ : std_logic;
signal \N__34480\ : std_logic;
signal \N__34477\ : std_logic;
signal \N__34472\ : std_logic;
signal \N__34469\ : std_logic;
signal \N__34466\ : std_logic;
signal \N__34463\ : std_logic;
signal \N__34460\ : std_logic;
signal \N__34457\ : std_logic;
signal \N__34454\ : std_logic;
signal \N__34453\ : std_logic;
signal \N__34452\ : std_logic;
signal \N__34451\ : std_logic;
signal \N__34450\ : std_logic;
signal \N__34447\ : std_logic;
signal \N__34444\ : std_logic;
signal \N__34439\ : std_logic;
signal \N__34436\ : std_logic;
signal \N__34431\ : std_logic;
signal \N__34428\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34422\ : std_logic;
signal \N__34419\ : std_logic;
signal \N__34412\ : std_logic;
signal \N__34411\ : std_logic;
signal \N__34410\ : std_logic;
signal \N__34407\ : std_logic;
signal \N__34404\ : std_logic;
signal \N__34401\ : std_logic;
signal \N__34396\ : std_logic;
signal \N__34393\ : std_logic;
signal \N__34390\ : std_logic;
signal \N__34387\ : std_logic;
signal \N__34384\ : std_logic;
signal \N__34379\ : std_logic;
signal \N__34378\ : std_logic;
signal \N__34375\ : std_logic;
signal \N__34372\ : std_logic;
signal \N__34371\ : std_logic;
signal \N__34368\ : std_logic;
signal \N__34363\ : std_logic;
signal \N__34358\ : std_logic;
signal \N__34355\ : std_logic;
signal \N__34352\ : std_logic;
signal \N__34349\ : std_logic;
signal \N__34346\ : std_logic;
signal \N__34345\ : std_logic;
signal \N__34342\ : std_logic;
signal \N__34341\ : std_logic;
signal \N__34340\ : std_logic;
signal \N__34337\ : std_logic;
signal \N__34334\ : std_logic;
signal \N__34329\ : std_logic;
signal \N__34322\ : std_logic;
signal \N__34321\ : std_logic;
signal \N__34318\ : std_logic;
signal \N__34315\ : std_logic;
signal \N__34314\ : std_logic;
signal \N__34309\ : std_logic;
signal \N__34306\ : std_logic;
signal \N__34303\ : std_logic;
signal \N__34298\ : std_logic;
signal \N__34295\ : std_logic;
signal \N__34294\ : std_logic;
signal \N__34293\ : std_logic;
signal \N__34292\ : std_logic;
signal \N__34287\ : std_logic;
signal \N__34286\ : std_logic;
signal \N__34285\ : std_logic;
signal \N__34280\ : std_logic;
signal \N__34277\ : std_logic;
signal \N__34274\ : std_logic;
signal \N__34271\ : std_logic;
signal \N__34268\ : std_logic;
signal \N__34259\ : std_logic;
signal \N__34256\ : std_logic;
signal \N__34253\ : std_logic;
signal \N__34252\ : std_logic;
signal \N__34249\ : std_logic;
signal \N__34248\ : std_logic;
signal \N__34245\ : std_logic;
signal \N__34242\ : std_logic;
signal \N__34239\ : std_logic;
signal \N__34238\ : std_logic;
signal \N__34235\ : std_logic;
signal \N__34232\ : std_logic;
signal \N__34227\ : std_logic;
signal \N__34220\ : std_logic;
signal \N__34219\ : std_logic;
signal \N__34216\ : std_logic;
signal \N__34213\ : std_logic;
signal \N__34208\ : std_logic;
signal \N__34205\ : std_logic;
signal \N__34202\ : std_logic;
signal \N__34201\ : std_logic;
signal \N__34196\ : std_logic;
signal \N__34193\ : std_logic;
signal \N__34190\ : std_logic;
signal \N__34187\ : std_logic;
signal \N__34184\ : std_logic;
signal \N__34181\ : std_logic;
signal \N__34178\ : std_logic;
signal \N__34177\ : std_logic;
signal \N__34176\ : std_logic;
signal \N__34173\ : std_logic;
signal \N__34170\ : std_logic;
signal \N__34167\ : std_logic;
signal \N__34162\ : std_logic;
signal \N__34159\ : std_logic;
signal \N__34156\ : std_logic;
signal \N__34153\ : std_logic;
signal \N__34150\ : std_logic;
signal \N__34145\ : std_logic;
signal \N__34142\ : std_logic;
signal \N__34141\ : std_logic;
signal \N__34140\ : std_logic;
signal \N__34137\ : std_logic;
signal \N__34136\ : std_logic;
signal \N__34133\ : std_logic;
signal \N__34130\ : std_logic;
signal \N__34127\ : std_logic;
signal \N__34124\ : std_logic;
signal \N__34123\ : std_logic;
signal \N__34120\ : std_logic;
signal \N__34113\ : std_logic;
signal \N__34110\ : std_logic;
signal \N__34105\ : std_logic;
signal \N__34102\ : std_logic;
signal \N__34099\ : std_logic;
signal \N__34094\ : std_logic;
signal \N__34091\ : std_logic;
signal \N__34088\ : std_logic;
signal \N__34085\ : std_logic;
signal \N__34082\ : std_logic;
signal \N__34079\ : std_logic;
signal \N__34076\ : std_logic;
signal \N__34073\ : std_logic;
signal \N__34070\ : std_logic;
signal \N__34067\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34061\ : std_logic;
signal \N__34058\ : std_logic;
signal \N__34055\ : std_logic;
signal \N__34052\ : std_logic;
signal \N__34049\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34043\ : std_logic;
signal \N__34040\ : std_logic;
signal \N__34037\ : std_logic;
signal \N__34034\ : std_logic;
signal \N__34031\ : std_logic;
signal \N__34028\ : std_logic;
signal \N__34025\ : std_logic;
signal \N__34022\ : std_logic;
signal \N__34019\ : std_logic;
signal \N__34016\ : std_logic;
signal \N__34013\ : std_logic;
signal \N__34010\ : std_logic;
signal \N__34007\ : std_logic;
signal \N__34004\ : std_logic;
signal \N__34001\ : std_logic;
signal \N__33998\ : std_logic;
signal \N__33995\ : std_logic;
signal \N__33994\ : std_logic;
signal \N__33991\ : std_logic;
signal \N__33988\ : std_logic;
signal \N__33987\ : std_logic;
signal \N__33984\ : std_logic;
signal \N__33981\ : std_logic;
signal \N__33978\ : std_logic;
signal \N__33975\ : std_logic;
signal \N__33972\ : std_logic;
signal \N__33969\ : std_logic;
signal \N__33966\ : std_logic;
signal \N__33961\ : std_logic;
signal \N__33958\ : std_logic;
signal \N__33955\ : std_logic;
signal \N__33950\ : std_logic;
signal \N__33949\ : std_logic;
signal \N__33946\ : std_logic;
signal \N__33945\ : std_logic;
signal \N__33942\ : std_logic;
signal \N__33941\ : std_logic;
signal \N__33938\ : std_logic;
signal \N__33935\ : std_logic;
signal \N__33930\ : std_logic;
signal \N__33927\ : std_logic;
signal \N__33920\ : std_logic;
signal \N__33917\ : std_logic;
signal \N__33914\ : std_logic;
signal \N__33911\ : std_logic;
signal \N__33908\ : std_logic;
signal \N__33905\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33899\ : std_logic;
signal \N__33896\ : std_logic;
signal \N__33895\ : std_logic;
signal \N__33892\ : std_logic;
signal \N__33889\ : std_logic;
signal \N__33884\ : std_logic;
signal \N__33883\ : std_logic;
signal \N__33880\ : std_logic;
signal \N__33877\ : std_logic;
signal \N__33872\ : std_logic;
signal \N__33871\ : std_logic;
signal \N__33868\ : std_logic;
signal \N__33865\ : std_logic;
signal \N__33864\ : std_logic;
signal \N__33861\ : std_logic;
signal \N__33856\ : std_logic;
signal \N__33851\ : std_logic;
signal \N__33848\ : std_logic;
signal \N__33845\ : std_logic;
signal \N__33844\ : std_logic;
signal \N__33841\ : std_logic;
signal \N__33838\ : std_logic;
signal \N__33833\ : std_logic;
signal \N__33830\ : std_logic;
signal \N__33827\ : std_logic;
signal \N__33824\ : std_logic;
signal \N__33821\ : std_logic;
signal \N__33818\ : std_logic;
signal \N__33817\ : std_logic;
signal \N__33814\ : std_logic;
signal \N__33813\ : std_logic;
signal \N__33806\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33802\ : std_logic;
signal \N__33797\ : std_logic;
signal \N__33794\ : std_logic;
signal \N__33791\ : std_logic;
signal \N__33788\ : std_logic;
signal \N__33785\ : std_logic;
signal \N__33782\ : std_logic;
signal \N__33779\ : std_logic;
signal \N__33778\ : std_logic;
signal \N__33775\ : std_logic;
signal \N__33774\ : std_logic;
signal \N__33771\ : std_logic;
signal \N__33766\ : std_logic;
signal \N__33761\ : std_logic;
signal \N__33760\ : std_logic;
signal \N__33755\ : std_logic;
signal \N__33752\ : std_logic;
signal \N__33749\ : std_logic;
signal \N__33746\ : std_logic;
signal \N__33743\ : std_logic;
signal \N__33742\ : std_logic;
signal \N__33739\ : std_logic;
signal \N__33736\ : std_logic;
signal \N__33731\ : std_logic;
signal \N__33730\ : std_logic;
signal \N__33729\ : std_logic;
signal \N__33726\ : std_logic;
signal \N__33723\ : std_logic;
signal \N__33722\ : std_logic;
signal \N__33719\ : std_logic;
signal \N__33718\ : std_logic;
signal \N__33715\ : std_logic;
signal \N__33712\ : std_logic;
signal \N__33709\ : std_logic;
signal \N__33706\ : std_logic;
signal \N__33703\ : std_logic;
signal \N__33700\ : std_logic;
signal \N__33697\ : std_logic;
signal \N__33694\ : std_logic;
signal \N__33693\ : std_logic;
signal \N__33688\ : std_logic;
signal \N__33683\ : std_logic;
signal \N__33680\ : std_logic;
signal \N__33677\ : std_logic;
signal \N__33674\ : std_logic;
signal \N__33671\ : std_logic;
signal \N__33668\ : std_logic;
signal \N__33665\ : std_logic;
signal \N__33662\ : std_logic;
signal \N__33655\ : std_logic;
signal \N__33652\ : std_logic;
signal \N__33649\ : std_logic;
signal \N__33644\ : std_logic;
signal \N__33641\ : std_logic;
signal \N__33638\ : std_logic;
signal \N__33635\ : std_logic;
signal \N__33632\ : std_logic;
signal \N__33629\ : std_logic;
signal \N__33626\ : std_logic;
signal \N__33625\ : std_logic;
signal \N__33622\ : std_logic;
signal \N__33619\ : std_logic;
signal \N__33614\ : std_logic;
signal \N__33611\ : std_logic;
signal \N__33608\ : std_logic;
signal \N__33605\ : std_logic;
signal \N__33602\ : std_logic;
signal \N__33599\ : std_logic;
signal \N__33596\ : std_logic;
signal \N__33593\ : std_logic;
signal \N__33590\ : std_logic;
signal \N__33587\ : std_logic;
signal \N__33584\ : std_logic;
signal \N__33581\ : std_logic;
signal \N__33578\ : std_logic;
signal \N__33575\ : std_logic;
signal \N__33572\ : std_logic;
signal \N__33569\ : std_logic;
signal \N__33566\ : std_logic;
signal \N__33565\ : std_logic;
signal \N__33562\ : std_logic;
signal \N__33561\ : std_logic;
signal \N__33558\ : std_logic;
signal \N__33557\ : std_logic;
signal \N__33556\ : std_logic;
signal \N__33553\ : std_logic;
signal \N__33550\ : std_logic;
signal \N__33547\ : std_logic;
signal \N__33544\ : std_logic;
signal \N__33541\ : std_logic;
signal \N__33540\ : std_logic;
signal \N__33537\ : std_logic;
signal \N__33534\ : std_logic;
signal \N__33529\ : std_logic;
signal \N__33526\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33518\ : std_logic;
signal \N__33515\ : std_logic;
signal \N__33512\ : std_logic;
signal \N__33509\ : std_logic;
signal \N__33504\ : std_logic;
signal \N__33499\ : std_logic;
signal \N__33494\ : std_logic;
signal \N__33491\ : std_logic;
signal \N__33488\ : std_logic;
signal \N__33485\ : std_logic;
signal \N__33482\ : std_logic;
signal \N__33479\ : std_logic;
signal \N__33476\ : std_logic;
signal \N__33473\ : std_logic;
signal \N__33470\ : std_logic;
signal \N__33467\ : std_logic;
signal \N__33464\ : std_logic;
signal \N__33461\ : std_logic;
signal \N__33458\ : std_logic;
signal \N__33455\ : std_logic;
signal \N__33452\ : std_logic;
signal \N__33449\ : std_logic;
signal \N__33446\ : std_logic;
signal \N__33443\ : std_logic;
signal \N__33440\ : std_logic;
signal \N__33437\ : std_logic;
signal \N__33434\ : std_logic;
signal \N__33431\ : std_logic;
signal \N__33428\ : std_logic;
signal \N__33425\ : std_logic;
signal \N__33422\ : std_logic;
signal \N__33419\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33413\ : std_logic;
signal \N__33410\ : std_logic;
signal \N__33407\ : std_logic;
signal \N__33404\ : std_logic;
signal \N__33401\ : std_logic;
signal \N__33398\ : std_logic;
signal \N__33395\ : std_logic;
signal \N__33392\ : std_logic;
signal \N__33389\ : std_logic;
signal \N__33386\ : std_logic;
signal \N__33383\ : std_logic;
signal \N__33380\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33374\ : std_logic;
signal \N__33371\ : std_logic;
signal \N__33368\ : std_logic;
signal \N__33365\ : std_logic;
signal \N__33362\ : std_logic;
signal \N__33359\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33353\ : std_logic;
signal \N__33350\ : std_logic;
signal \N__33347\ : std_logic;
signal \N__33344\ : std_logic;
signal \N__33341\ : std_logic;
signal \N__33338\ : std_logic;
signal \N__33335\ : std_logic;
signal \N__33332\ : std_logic;
signal \N__33329\ : std_logic;
signal \N__33326\ : std_logic;
signal \N__33323\ : std_logic;
signal \N__33320\ : std_logic;
signal \N__33317\ : std_logic;
signal \N__33314\ : std_logic;
signal \N__33311\ : std_logic;
signal \N__33308\ : std_logic;
signal \N__33305\ : std_logic;
signal \N__33302\ : std_logic;
signal \N__33299\ : std_logic;
signal \N__33296\ : std_logic;
signal \N__33293\ : std_logic;
signal \N__33290\ : std_logic;
signal \N__33287\ : std_logic;
signal \N__33284\ : std_logic;
signal \N__33281\ : std_logic;
signal \N__33278\ : std_logic;
signal \N__33275\ : std_logic;
signal \N__33272\ : std_logic;
signal \N__33269\ : std_logic;
signal \N__33266\ : std_logic;
signal \N__33263\ : std_logic;
signal \N__33260\ : std_logic;
signal \N__33257\ : std_logic;
signal \N__33254\ : std_logic;
signal \N__33251\ : std_logic;
signal \N__33248\ : std_logic;
signal \N__33245\ : std_logic;
signal \N__33242\ : std_logic;
signal \N__33239\ : std_logic;
signal \N__33236\ : std_logic;
signal \N__33233\ : std_logic;
signal \N__33230\ : std_logic;
signal \N__33227\ : std_logic;
signal \N__33224\ : std_logic;
signal \N__33221\ : std_logic;
signal \N__33218\ : std_logic;
signal \N__33215\ : std_logic;
signal \N__33212\ : std_logic;
signal \N__33209\ : std_logic;
signal \N__33206\ : std_logic;
signal \N__33203\ : std_logic;
signal \N__33200\ : std_logic;
signal \N__33197\ : std_logic;
signal \N__33194\ : std_logic;
signal \N__33191\ : std_logic;
signal \N__33188\ : std_logic;
signal \N__33185\ : std_logic;
signal \N__33182\ : std_logic;
signal \N__33179\ : std_logic;
signal \N__33176\ : std_logic;
signal \N__33173\ : std_logic;
signal \N__33170\ : std_logic;
signal \N__33167\ : std_logic;
signal \N__33164\ : std_logic;
signal \N__33161\ : std_logic;
signal \N__33158\ : std_logic;
signal \N__33155\ : std_logic;
signal \N__33152\ : std_logic;
signal \N__33149\ : std_logic;
signal \N__33146\ : std_logic;
signal \N__33143\ : std_logic;
signal \N__33142\ : std_logic;
signal \N__33139\ : std_logic;
signal \N__33136\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33119\ : std_logic;
signal \N__33116\ : std_logic;
signal \N__33113\ : std_logic;
signal \N__33110\ : std_logic;
signal \N__33107\ : std_logic;
signal \N__33104\ : std_logic;
signal \N__33101\ : std_logic;
signal \N__33098\ : std_logic;
signal \N__33095\ : std_logic;
signal \N__33092\ : std_logic;
signal \N__33089\ : std_logic;
signal \N__33086\ : std_logic;
signal \N__33083\ : std_logic;
signal \N__33082\ : std_logic;
signal \N__33081\ : std_logic;
signal \N__33080\ : std_logic;
signal \N__33079\ : std_logic;
signal \N__33078\ : std_logic;
signal \N__33077\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33075\ : std_logic;
signal \N__33074\ : std_logic;
signal \N__33073\ : std_logic;
signal \N__33070\ : std_logic;
signal \N__33069\ : std_logic;
signal \N__33068\ : std_logic;
signal \N__33067\ : std_logic;
signal \N__33066\ : std_logic;
signal \N__33065\ : std_logic;
signal \N__33064\ : std_logic;
signal \N__33063\ : std_logic;
signal \N__33062\ : std_logic;
signal \N__33045\ : std_logic;
signal \N__33042\ : std_logic;
signal \N__33041\ : std_logic;
signal \N__33038\ : std_logic;
signal \N__33037\ : std_logic;
signal \N__33036\ : std_logic;
signal \N__33035\ : std_logic;
signal \N__33034\ : std_logic;
signal \N__33031\ : std_logic;
signal \N__33028\ : std_logic;
signal \N__33015\ : std_logic;
signal \N__33012\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33010\ : std_logic;
signal \N__33009\ : std_logic;
signal \N__33008\ : std_logic;
signal \N__33007\ : std_logic;
signal \N__33006\ : std_logic;
signal \N__33005\ : std_logic;
signal \N__33004\ : std_logic;
signal \N__33003\ : std_logic;
signal \N__33000\ : std_logic;
signal \N__32997\ : std_logic;
signal \N__32994\ : std_logic;
signal \N__32991\ : std_logic;
signal \N__32982\ : std_logic;
signal \N__32979\ : std_logic;
signal \N__32976\ : std_logic;
signal \N__32971\ : std_logic;
signal \N__32968\ : std_logic;
signal \N__32963\ : std_logic;
signal \N__32958\ : std_logic;
signal \N__32955\ : std_logic;
signal \N__32950\ : std_logic;
signal \N__32947\ : std_logic;
signal \N__32944\ : std_logic;
signal \N__32939\ : std_logic;
signal \N__32926\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32908\ : std_logic;
signal \N__32907\ : std_logic;
signal \N__32904\ : std_logic;
signal \N__32901\ : std_logic;
signal \N__32900\ : std_logic;
signal \N__32899\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32897\ : std_logic;
signal \N__32896\ : std_logic;
signal \N__32895\ : std_logic;
signal \N__32892\ : std_logic;
signal \N__32891\ : std_logic;
signal \N__32888\ : std_logic;
signal \N__32885\ : std_logic;
signal \N__32882\ : std_logic;
signal \N__32881\ : std_logic;
signal \N__32870\ : std_logic;
signal \N__32865\ : std_logic;
signal \N__32864\ : std_logic;
signal \N__32863\ : std_logic;
signal \N__32862\ : std_logic;
signal \N__32861\ : std_logic;
signal \N__32860\ : std_logic;
signal \N__32859\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32846\ : std_logic;
signal \N__32843\ : std_logic;
signal \N__32842\ : std_logic;
signal \N__32841\ : std_logic;
signal \N__32840\ : std_logic;
signal \N__32839\ : std_logic;
signal \N__32838\ : std_logic;
signal \N__32837\ : std_logic;
signal \N__32836\ : std_logic;
signal \N__32835\ : std_logic;
signal \N__32834\ : std_logic;
signal \N__32831\ : std_logic;
signal \N__32830\ : std_logic;
signal \N__32827\ : std_logic;
signal \N__32826\ : std_logic;
signal \N__32825\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32819\ : std_logic;
signal \N__32816\ : std_logic;
signal \N__32815\ : std_logic;
signal \N__32812\ : std_logic;
signal \N__32811\ : std_logic;
signal \N__32810\ : std_logic;
signal \N__32807\ : std_logic;
signal \N__32804\ : std_logic;
signal \N__32799\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32783\ : std_logic;
signal \N__32770\ : std_logic;
signal \N__32753\ : std_logic;
signal \N__32738\ : std_logic;
signal \N__32735\ : std_logic;
signal \N__32732\ : std_logic;
signal \N__32729\ : std_logic;
signal \N__32726\ : std_logic;
signal \N__32723\ : std_logic;
signal \N__32722\ : std_logic;
signal \N__32721\ : std_logic;
signal \N__32720\ : std_logic;
signal \N__32717\ : std_logic;
signal \N__32716\ : std_logic;
signal \N__32715\ : std_logic;
signal \N__32714\ : std_logic;
signal \N__32713\ : std_logic;
signal \N__32712\ : std_logic;
signal \N__32711\ : std_logic;
signal \N__32710\ : std_logic;
signal \N__32709\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32707\ : std_logic;
signal \N__32706\ : std_logic;
signal \N__32705\ : std_logic;
signal \N__32704\ : std_logic;
signal \N__32703\ : std_logic;
signal \N__32698\ : std_logic;
signal \N__32695\ : std_logic;
signal \N__32694\ : std_logic;
signal \N__32693\ : std_logic;
signal \N__32692\ : std_logic;
signal \N__32691\ : std_logic;
signal \N__32688\ : std_logic;
signal \N__32671\ : std_logic;
signal \N__32658\ : std_logic;
signal \N__32657\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32655\ : std_logic;
signal \N__32654\ : std_logic;
signal \N__32653\ : std_logic;
signal \N__32648\ : std_logic;
signal \N__32639\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32629\ : std_logic;
signal \N__32618\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32597\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32593\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32589\ : std_logic;
signal \N__32588\ : std_logic;
signal \N__32585\ : std_logic;
signal \N__32582\ : std_logic;
signal \N__32579\ : std_logic;
signal \N__32576\ : std_logic;
signal \N__32573\ : std_logic;
signal \N__32566\ : std_logic;
signal \N__32561\ : std_logic;
signal \N__32560\ : std_logic;
signal \N__32559\ : std_logic;
signal \N__32556\ : std_logic;
signal \N__32555\ : std_logic;
signal \N__32554\ : std_logic;
signal \N__32553\ : std_logic;
signal \N__32552\ : std_logic;
signal \N__32551\ : std_logic;
signal \N__32550\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32548\ : std_logic;
signal \N__32547\ : std_logic;
signal \N__32544\ : std_logic;
signal \N__32541\ : std_logic;
signal \N__32540\ : std_logic;
signal \N__32537\ : std_logic;
signal \N__32534\ : std_logic;
signal \N__32531\ : std_logic;
signal \N__32530\ : std_logic;
signal \N__32527\ : std_logic;
signal \N__32524\ : std_logic;
signal \N__32521\ : std_logic;
signal \N__32518\ : std_logic;
signal \N__32515\ : std_logic;
signal \N__32514\ : std_logic;
signal \N__32513\ : std_logic;
signal \N__32510\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32504\ : std_logic;
signal \N__32501\ : std_logic;
signal \N__32498\ : std_logic;
signal \N__32497\ : std_logic;
signal \N__32492\ : std_logic;
signal \N__32491\ : std_logic;
signal \N__32490\ : std_logic;
signal \N__32489\ : std_logic;
signal \N__32486\ : std_logic;
signal \N__32485\ : std_logic;
signal \N__32484\ : std_logic;
signal \N__32481\ : std_logic;
signal \N__32480\ : std_logic;
signal \N__32477\ : std_logic;
signal \N__32470\ : std_logic;
signal \N__32467\ : std_logic;
signal \N__32464\ : std_logic;
signal \N__32461\ : std_logic;
signal \N__32456\ : std_logic;
signal \N__32453\ : std_logic;
signal \N__32448\ : std_logic;
signal \N__32445\ : std_logic;
signal \N__32442\ : std_logic;
signal \N__32439\ : std_logic;
signal \N__32436\ : std_logic;
signal \N__32433\ : std_logic;
signal \N__32432\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32426\ : std_logic;
signal \N__32423\ : std_logic;
signal \N__32420\ : std_logic;
signal \N__32417\ : std_logic;
signal \N__32414\ : std_logic;
signal \N__32411\ : std_logic;
signal \N__32404\ : std_logic;
signal \N__32401\ : std_logic;
signal \N__32396\ : std_logic;
signal \N__32393\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32381\ : std_logic;
signal \N__32376\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32370\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32358\ : std_logic;
signal \N__32349\ : std_logic;
signal \N__32344\ : std_logic;
signal \N__32333\ : std_logic;
signal \N__32330\ : std_logic;
signal \N__32327\ : std_logic;
signal \N__32324\ : std_logic;
signal \N__32321\ : std_logic;
signal \N__32318\ : std_logic;
signal \N__32317\ : std_logic;
signal \N__32314\ : std_logic;
signal \N__32311\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32305\ : std_logic;
signal \N__32302\ : std_logic;
signal \N__32299\ : std_logic;
signal \N__32296\ : std_logic;
signal \N__32293\ : std_logic;
signal \N__32292\ : std_logic;
signal \N__32289\ : std_logic;
signal \N__32286\ : std_logic;
signal \N__32283\ : std_logic;
signal \N__32280\ : std_logic;
signal \N__32277\ : std_logic;
signal \N__32274\ : std_logic;
signal \N__32267\ : std_logic;
signal \N__32264\ : std_logic;
signal \N__32261\ : std_logic;
signal \N__32258\ : std_logic;
signal \N__32255\ : std_logic;
signal \N__32254\ : std_logic;
signal \N__32249\ : std_logic;
signal \N__32246\ : std_logic;
signal \N__32245\ : std_logic;
signal \N__32240\ : std_logic;
signal \N__32239\ : std_logic;
signal \N__32236\ : std_logic;
signal \N__32233\ : std_logic;
signal \N__32230\ : std_logic;
signal \N__32225\ : std_logic;
signal \N__32222\ : std_logic;
signal \N__32219\ : std_logic;
signal \N__32216\ : std_logic;
signal \N__32215\ : std_logic;
signal \N__32212\ : std_logic;
signal \N__32209\ : std_logic;
signal \N__32204\ : std_logic;
signal \N__32203\ : std_logic;
signal \N__32200\ : std_logic;
signal \N__32197\ : std_logic;
signal \N__32194\ : std_logic;
signal \N__32189\ : std_logic;
signal \N__32186\ : std_logic;
signal \N__32183\ : std_logic;
signal \N__32180\ : std_logic;
signal \N__32179\ : std_logic;
signal \N__32176\ : std_logic;
signal \N__32173\ : std_logic;
signal \N__32168\ : std_logic;
signal \N__32167\ : std_logic;
signal \N__32164\ : std_logic;
signal \N__32161\ : std_logic;
signal \N__32158\ : std_logic;
signal \N__32153\ : std_logic;
signal \N__32150\ : std_logic;
signal \N__32147\ : std_logic;
signal \N__32144\ : std_logic;
signal \N__32143\ : std_logic;
signal \N__32140\ : std_logic;
signal \N__32137\ : std_logic;
signal \N__32136\ : std_logic;
signal \N__32133\ : std_logic;
signal \N__32130\ : std_logic;
signal \N__32127\ : std_logic;
signal \N__32124\ : std_logic;
signal \N__32121\ : std_logic;
signal \N__32114\ : std_logic;
signal \N__32111\ : std_logic;
signal \N__32108\ : std_logic;
signal \N__32105\ : std_logic;
signal \N__32104\ : std_logic;
signal \N__32101\ : std_logic;
signal \N__32098\ : std_logic;
signal \N__32097\ : std_logic;
signal \N__32094\ : std_logic;
signal \N__32091\ : std_logic;
signal \N__32088\ : std_logic;
signal \N__32085\ : std_logic;
signal \N__32082\ : std_logic;
signal \N__32075\ : std_logic;
signal \N__32072\ : std_logic;
signal \N__32069\ : std_logic;
signal \N__32066\ : std_logic;
signal \N__32063\ : std_logic;
signal \N__32062\ : std_logic;
signal \N__32059\ : std_logic;
signal \N__32056\ : std_logic;
signal \N__32053\ : std_logic;
signal \N__32048\ : std_logic;
signal \N__32047\ : std_logic;
signal \N__32044\ : std_logic;
signal \N__32041\ : std_logic;
signal \N__32040\ : std_logic;
signal \N__32035\ : std_logic;
signal \N__32032\ : std_logic;
signal \N__32029\ : std_logic;
signal \N__32024\ : std_logic;
signal \N__32021\ : std_logic;
signal \N__32018\ : std_logic;
signal \N__32015\ : std_logic;
signal \N__32012\ : std_logic;
signal \N__32009\ : std_logic;
signal \N__32008\ : std_logic;
signal \N__32005\ : std_logic;
signal \N__32002\ : std_logic;
signal \N__31999\ : std_logic;
signal \N__31994\ : std_logic;
signal \N__31993\ : std_logic;
signal \N__31990\ : std_logic;
signal \N__31987\ : std_logic;
signal \N__31986\ : std_logic;
signal \N__31981\ : std_logic;
signal \N__31978\ : std_logic;
signal \N__31975\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31961\ : std_logic;
signal \N__31958\ : std_logic;
signal \N__31957\ : std_logic;
signal \N__31956\ : std_logic;
signal \N__31955\ : std_logic;
signal \N__31954\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31940\ : std_logic;
signal \N__31937\ : std_logic;
signal \N__31934\ : std_logic;
signal \N__31931\ : std_logic;
signal \N__31928\ : std_logic;
signal \N__31927\ : std_logic;
signal \N__31924\ : std_logic;
signal \N__31921\ : std_logic;
signal \N__31918\ : std_logic;
signal \N__31915\ : std_logic;
signal \N__31910\ : std_logic;
signal \N__31907\ : std_logic;
signal \N__31906\ : std_logic;
signal \N__31901\ : std_logic;
signal \N__31900\ : std_logic;
signal \N__31897\ : std_logic;
signal \N__31894\ : std_logic;
signal \N__31891\ : std_logic;
signal \N__31886\ : std_logic;
signal \N__31883\ : std_logic;
signal \N__31880\ : std_logic;
signal \N__31877\ : std_logic;
signal \N__31876\ : std_logic;
signal \N__31873\ : std_logic;
signal \N__31870\ : std_logic;
signal \N__31865\ : std_logic;
signal \N__31864\ : std_logic;
signal \N__31861\ : std_logic;
signal \N__31858\ : std_logic;
signal \N__31855\ : std_logic;
signal \N__31850\ : std_logic;
signal \N__31847\ : std_logic;
signal \N__31844\ : std_logic;
signal \N__31841\ : std_logic;
signal \N__31840\ : std_logic;
signal \N__31837\ : std_logic;
signal \N__31834\ : std_logic;
signal \N__31829\ : std_logic;
signal \N__31828\ : std_logic;
signal \N__31825\ : std_logic;
signal \N__31822\ : std_logic;
signal \N__31819\ : std_logic;
signal \N__31814\ : std_logic;
signal \N__31811\ : std_logic;
signal \N__31808\ : std_logic;
signal \N__31805\ : std_logic;
signal \N__31804\ : std_logic;
signal \N__31801\ : std_logic;
signal \N__31798\ : std_logic;
signal \N__31797\ : std_logic;
signal \N__31794\ : std_logic;
signal \N__31791\ : std_logic;
signal \N__31788\ : std_logic;
signal \N__31785\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31775\ : std_logic;
signal \N__31772\ : std_logic;
signal \N__31769\ : std_logic;
signal \N__31766\ : std_logic;
signal \N__31765\ : std_logic;
signal \N__31762\ : std_logic;
signal \N__31759\ : std_logic;
signal \N__31758\ : std_logic;
signal \N__31755\ : std_logic;
signal \N__31752\ : std_logic;
signal \N__31749\ : std_logic;
signal \N__31746\ : std_logic;
signal \N__31743\ : std_logic;
signal \N__31736\ : std_logic;
signal \N__31733\ : std_logic;
signal \N__31730\ : std_logic;
signal \N__31727\ : std_logic;
signal \N__31726\ : std_logic;
signal \N__31723\ : std_logic;
signal \N__31720\ : std_logic;
signal \N__31719\ : std_logic;
signal \N__31714\ : std_logic;
signal \N__31711\ : std_logic;
signal \N__31708\ : std_logic;
signal \N__31703\ : std_logic;
signal \N__31700\ : std_logic;
signal \N__31697\ : std_logic;
signal \N__31694\ : std_logic;
signal \N__31691\ : std_logic;
signal \N__31690\ : std_logic;
signal \N__31687\ : std_logic;
signal \N__31684\ : std_logic;
signal \N__31683\ : std_logic;
signal \N__31678\ : std_logic;
signal \N__31675\ : std_logic;
signal \N__31672\ : std_logic;
signal \N__31667\ : std_logic;
signal \N__31664\ : std_logic;
signal \N__31661\ : std_logic;
signal \N__31658\ : std_logic;
signal \N__31655\ : std_logic;
signal \N__31654\ : std_logic;
signal \N__31649\ : std_logic;
signal \N__31648\ : std_logic;
signal \N__31645\ : std_logic;
signal \N__31642\ : std_logic;
signal \N__31639\ : std_logic;
signal \N__31634\ : std_logic;
signal \N__31631\ : std_logic;
signal \N__31628\ : std_logic;
signal \N__31625\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31621\ : std_logic;
signal \N__31616\ : std_logic;
signal \N__31615\ : std_logic;
signal \N__31612\ : std_logic;
signal \N__31609\ : std_logic;
signal \N__31606\ : std_logic;
signal \N__31601\ : std_logic;
signal \N__31598\ : std_logic;
signal \N__31595\ : std_logic;
signal \N__31592\ : std_logic;
signal \N__31591\ : std_logic;
signal \N__31586\ : std_logic;
signal \N__31585\ : std_logic;
signal \N__31582\ : std_logic;
signal \N__31579\ : std_logic;
signal \N__31576\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31568\ : std_logic;
signal \N__31565\ : std_logic;
signal \N__31562\ : std_logic;
signal \N__31561\ : std_logic;
signal \N__31558\ : std_logic;
signal \N__31555\ : std_logic;
signal \N__31552\ : std_logic;
signal \N__31551\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31545\ : std_logic;
signal \N__31542\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31536\ : std_logic;
signal \N__31529\ : std_logic;
signal \N__31526\ : std_logic;
signal \N__31523\ : std_logic;
signal \N__31520\ : std_logic;
signal \N__31519\ : std_logic;
signal \N__31516\ : std_logic;
signal \N__31513\ : std_logic;
signal \N__31510\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31503\ : std_logic;
signal \N__31500\ : std_logic;
signal \N__31497\ : std_logic;
signal \N__31494\ : std_logic;
signal \N__31487\ : std_logic;
signal \N__31484\ : std_logic;
signal \N__31481\ : std_logic;
signal \N__31478\ : std_logic;
signal \N__31477\ : std_logic;
signal \N__31474\ : std_logic;
signal \N__31471\ : std_logic;
signal \N__31470\ : std_logic;
signal \N__31465\ : std_logic;
signal \N__31462\ : std_logic;
signal \N__31459\ : std_logic;
signal \N__31454\ : std_logic;
signal \N__31451\ : std_logic;
signal \N__31448\ : std_logic;
signal \N__31445\ : std_logic;
signal \N__31442\ : std_logic;
signal \N__31441\ : std_logic;
signal \N__31438\ : std_logic;
signal \N__31435\ : std_logic;
signal \N__31434\ : std_logic;
signal \N__31429\ : std_logic;
signal \N__31426\ : std_logic;
signal \N__31423\ : std_logic;
signal \N__31418\ : std_logic;
signal \N__31415\ : std_logic;
signal \N__31412\ : std_logic;
signal \N__31409\ : std_logic;
signal \N__31406\ : std_logic;
signal \N__31403\ : std_logic;
signal \N__31402\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31396\ : std_logic;
signal \N__31393\ : std_logic;
signal \N__31390\ : std_logic;
signal \N__31387\ : std_logic;
signal \N__31382\ : std_logic;
signal \N__31379\ : std_logic;
signal \N__31376\ : std_logic;
signal \N__31373\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31367\ : std_logic;
signal \N__31366\ : std_logic;
signal \N__31363\ : std_logic;
signal \N__31360\ : std_logic;
signal \N__31357\ : std_logic;
signal \N__31354\ : std_logic;
signal \N__31353\ : std_logic;
signal \N__31350\ : std_logic;
signal \N__31347\ : std_logic;
signal \N__31344\ : std_logic;
signal \N__31337\ : std_logic;
signal \N__31336\ : std_logic;
signal \N__31333\ : std_logic;
signal \N__31332\ : std_logic;
signal \N__31329\ : std_logic;
signal \N__31324\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31320\ : std_logic;
signal \N__31317\ : std_logic;
signal \N__31314\ : std_logic;
signal \N__31311\ : std_logic;
signal \N__31308\ : std_logic;
signal \N__31305\ : std_logic;
signal \N__31298\ : std_logic;
signal \N__31295\ : std_logic;
signal \N__31292\ : std_logic;
signal \N__31289\ : std_logic;
signal \N__31286\ : std_logic;
signal \N__31283\ : std_logic;
signal \N__31282\ : std_logic;
signal \N__31279\ : std_logic;
signal \N__31276\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31271\ : std_logic;
signal \N__31268\ : std_logic;
signal \N__31265\ : std_logic;
signal \N__31262\ : std_logic;
signal \N__31259\ : std_logic;
signal \N__31256\ : std_logic;
signal \N__31253\ : std_logic;
signal \N__31250\ : std_logic;
signal \N__31247\ : std_logic;
signal \N__31242\ : std_logic;
signal \N__31235\ : std_logic;
signal \N__31232\ : std_logic;
signal \N__31231\ : std_logic;
signal \N__31230\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31224\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31220\ : std_logic;
signal \N__31215\ : std_logic;
signal \N__31212\ : std_logic;
signal \N__31209\ : std_logic;
signal \N__31206\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31200\ : std_logic;
signal \N__31193\ : std_logic;
signal \N__31190\ : std_logic;
signal \N__31189\ : std_logic;
signal \N__31188\ : std_logic;
signal \N__31185\ : std_logic;
signal \N__31182\ : std_logic;
signal \N__31179\ : std_logic;
signal \N__31178\ : std_logic;
signal \N__31175\ : std_logic;
signal \N__31172\ : std_logic;
signal \N__31169\ : std_logic;
signal \N__31166\ : std_logic;
signal \N__31163\ : std_logic;
signal \N__31160\ : std_logic;
signal \N__31157\ : std_logic;
signal \N__31154\ : std_logic;
signal \N__31145\ : std_logic;
signal \N__31142\ : std_logic;
signal \N__31141\ : std_logic;
signal \N__31140\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31132\ : std_logic;
signal \N__31129\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31125\ : std_logic;
signal \N__31122\ : std_logic;
signal \N__31119\ : std_logic;
signal \N__31112\ : std_logic;
signal \N__31109\ : std_logic;
signal \N__31106\ : std_logic;
signal \N__31103\ : std_logic;
signal \N__31100\ : std_logic;
signal \N__31099\ : std_logic;
signal \N__31096\ : std_logic;
signal \N__31093\ : std_logic;
signal \N__31090\ : std_logic;
signal \N__31087\ : std_logic;
signal \N__31086\ : std_logic;
signal \N__31083\ : std_logic;
signal \N__31080\ : std_logic;
signal \N__31077\ : std_logic;
signal \N__31074\ : std_logic;
signal \N__31067\ : std_logic;
signal \N__31064\ : std_logic;
signal \N__31061\ : std_logic;
signal \N__31060\ : std_logic;
signal \N__31057\ : std_logic;
signal \N__31054\ : std_logic;
signal \N__31051\ : std_logic;
signal \N__31048\ : std_logic;
signal \N__31047\ : std_logic;
signal \N__31044\ : std_logic;
signal \N__31041\ : std_logic;
signal \N__31038\ : std_logic;
signal \N__31035\ : std_logic;
signal \N__31028\ : std_logic;
signal \N__31025\ : std_logic;
signal \N__31022\ : std_logic;
signal \N__31019\ : std_logic;
signal \N__31018\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31012\ : std_logic;
signal \N__31009\ : std_logic;
signal \N__31006\ : std_logic;
signal \N__31001\ : std_logic;
signal \N__30998\ : std_logic;
signal \N__30995\ : std_logic;
signal \N__30992\ : std_logic;
signal \N__30989\ : std_logic;
signal \N__30988\ : std_logic;
signal \N__30987\ : std_logic;
signal \N__30982\ : std_logic;
signal \N__30979\ : std_logic;
signal \N__30976\ : std_logic;
signal \N__30971\ : std_logic;
signal \N__30968\ : std_logic;
signal \N__30965\ : std_logic;
signal \N__30962\ : std_logic;
signal \N__30959\ : std_logic;
signal \N__30958\ : std_logic;
signal \N__30955\ : std_logic;
signal \N__30952\ : std_logic;
signal \N__30947\ : std_logic;
signal \N__30946\ : std_logic;
signal \N__30943\ : std_logic;
signal \N__30940\ : std_logic;
signal \N__30937\ : std_logic;
signal \N__30932\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30926\ : std_logic;
signal \N__30923\ : std_logic;
signal \N__30922\ : std_logic;
signal \N__30919\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30911\ : std_logic;
signal \N__30910\ : std_logic;
signal \N__30907\ : std_logic;
signal \N__30904\ : std_logic;
signal \N__30901\ : std_logic;
signal \N__30896\ : std_logic;
signal \N__30893\ : std_logic;
signal \N__30890\ : std_logic;
signal \N__30887\ : std_logic;
signal \N__30886\ : std_logic;
signal \N__30885\ : std_logic;
signal \N__30882\ : std_logic;
signal \N__30879\ : std_logic;
signal \N__30876\ : std_logic;
signal \N__30871\ : std_logic;
signal \N__30868\ : std_logic;
signal \N__30867\ : std_logic;
signal \N__30864\ : std_logic;
signal \N__30861\ : std_logic;
signal \N__30858\ : std_logic;
signal \N__30855\ : std_logic;
signal \N__30850\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30844\ : std_logic;
signal \N__30843\ : std_logic;
signal \N__30840\ : std_logic;
signal \N__30837\ : std_logic;
signal \N__30834\ : std_logic;
signal \N__30831\ : std_logic;
signal \N__30828\ : std_logic;
signal \N__30827\ : std_logic;
signal \N__30824\ : std_logic;
signal \N__30819\ : std_logic;
signal \N__30816\ : std_logic;
signal \N__30809\ : std_logic;
signal \N__30806\ : std_logic;
signal \N__30805\ : std_logic;
signal \N__30802\ : std_logic;
signal \N__30801\ : std_logic;
signal \N__30798\ : std_logic;
signal \N__30797\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30788\ : std_logic;
signal \N__30785\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30776\ : std_logic;
signal \N__30773\ : std_logic;
signal \N__30764\ : std_logic;
signal \N__30763\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30759\ : std_logic;
signal \N__30756\ : std_logic;
signal \N__30753\ : std_logic;
signal \N__30750\ : std_logic;
signal \N__30747\ : std_logic;
signal \N__30746\ : std_logic;
signal \N__30741\ : std_logic;
signal \N__30738\ : std_logic;
signal \N__30735\ : std_logic;
signal \N__30728\ : std_logic;
signal \N__30725\ : std_logic;
signal \N__30722\ : std_logic;
signal \N__30719\ : std_logic;
signal \N__30716\ : std_logic;
signal \N__30713\ : std_logic;
signal \N__30710\ : std_logic;
signal \N__30707\ : std_logic;
signal \N__30704\ : std_logic;
signal \N__30701\ : std_logic;
signal \N__30698\ : std_logic;
signal \N__30697\ : std_logic;
signal \N__30696\ : std_logic;
signal \N__30693\ : std_logic;
signal \N__30690\ : std_logic;
signal \N__30687\ : std_logic;
signal \N__30684\ : std_logic;
signal \N__30683\ : std_logic;
signal \N__30680\ : std_logic;
signal \N__30677\ : std_logic;
signal \N__30674\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30661\ : std_logic;
signal \N__30656\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30654\ : std_logic;
signal \N__30651\ : std_logic;
signal \N__30648\ : std_logic;
signal \N__30645\ : std_logic;
signal \N__30644\ : std_logic;
signal \N__30641\ : std_logic;
signal \N__30638\ : std_logic;
signal \N__30635\ : std_logic;
signal \N__30632\ : std_logic;
signal \N__30629\ : std_logic;
signal \N__30624\ : std_logic;
signal \N__30621\ : std_logic;
signal \N__30614\ : std_logic;
signal \N__30611\ : std_logic;
signal \N__30608\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30598\ : std_logic;
signal \N__30597\ : std_logic;
signal \N__30596\ : std_logic;
signal \N__30593\ : std_logic;
signal \N__30590\ : std_logic;
signal \N__30585\ : std_logic;
signal \N__30582\ : std_logic;
signal \N__30579\ : std_logic;
signal \N__30576\ : std_logic;
signal \N__30571\ : std_logic;
signal \N__30566\ : std_logic;
signal \N__30563\ : std_logic;
signal \N__30562\ : std_logic;
signal \N__30561\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30553\ : std_logic;
signal \N__30552\ : std_logic;
signal \N__30549\ : std_logic;
signal \N__30546\ : std_logic;
signal \N__30543\ : std_logic;
signal \N__30540\ : std_logic;
signal \N__30537\ : std_logic;
signal \N__30534\ : std_logic;
signal \N__30527\ : std_logic;
signal \N__30524\ : std_logic;
signal \N__30521\ : std_logic;
signal \N__30518\ : std_logic;
signal \N__30515\ : std_logic;
signal \N__30512\ : std_logic;
signal \N__30509\ : std_logic;
signal \N__30508\ : std_logic;
signal \N__30507\ : std_logic;
signal \N__30506\ : std_logic;
signal \N__30503\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30495\ : std_logic;
signal \N__30492\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30486\ : std_logic;
signal \N__30483\ : std_logic;
signal \N__30480\ : std_logic;
signal \N__30477\ : std_logic;
signal \N__30470\ : std_logic;
signal \N__30467\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30465\ : std_logic;
signal \N__30460\ : std_logic;
signal \N__30459\ : std_logic;
signal \N__30456\ : std_logic;
signal \N__30453\ : std_logic;
signal \N__30450\ : std_logic;
signal \N__30447\ : std_logic;
signal \N__30444\ : std_logic;
signal \N__30441\ : std_logic;
signal \N__30434\ : std_logic;
signal \N__30431\ : std_logic;
signal \N__30428\ : std_logic;
signal \N__30425\ : std_logic;
signal \N__30422\ : std_logic;
signal \N__30419\ : std_logic;
signal \N__30416\ : std_logic;
signal \N__30413\ : std_logic;
signal \N__30410\ : std_logic;
signal \N__30407\ : std_logic;
signal \N__30404\ : std_logic;
signal \N__30403\ : std_logic;
signal \N__30402\ : std_logic;
signal \N__30399\ : std_logic;
signal \N__30396\ : std_logic;
signal \N__30393\ : std_logic;
signal \N__30392\ : std_logic;
signal \N__30389\ : std_logic;
signal \N__30386\ : std_logic;
signal \N__30381\ : std_logic;
signal \N__30378\ : std_logic;
signal \N__30375\ : std_logic;
signal \N__30372\ : std_logic;
signal \N__30365\ : std_logic;
signal \N__30362\ : std_logic;
signal \N__30359\ : std_logic;
signal \N__30356\ : std_logic;
signal \N__30353\ : std_logic;
signal \N__30350\ : std_logic;
signal \N__30349\ : std_logic;
signal \N__30348\ : std_logic;
signal \N__30347\ : std_logic;
signal \N__30344\ : std_logic;
signal \N__30341\ : std_logic;
signal \N__30336\ : std_logic;
signal \N__30333\ : std_logic;
signal \N__30330\ : std_logic;
signal \N__30327\ : std_logic;
signal \N__30320\ : std_logic;
signal \N__30317\ : std_logic;
signal \N__30314\ : std_logic;
signal \N__30311\ : std_logic;
signal \N__30308\ : std_logic;
signal \N__30305\ : std_logic;
signal \N__30302\ : std_logic;
signal \N__30301\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30293\ : std_logic;
signal \N__30290\ : std_logic;
signal \N__30289\ : std_logic;
signal \N__30286\ : std_logic;
signal \N__30285\ : std_logic;
signal \N__30282\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30280\ : std_logic;
signal \N__30279\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30272\ : std_logic;
signal \N__30265\ : std_logic;
signal \N__30262\ : std_logic;
signal \N__30259\ : std_logic;
signal \N__30248\ : std_logic;
signal \N__30247\ : std_logic;
signal \N__30246\ : std_logic;
signal \N__30245\ : std_logic;
signal \N__30244\ : std_logic;
signal \N__30237\ : std_logic;
signal \N__30234\ : std_logic;
signal \N__30233\ : std_logic;
signal \N__30232\ : std_logic;
signal \N__30229\ : std_logic;
signal \N__30226\ : std_logic;
signal \N__30223\ : std_logic;
signal \N__30220\ : std_logic;
signal \N__30217\ : std_logic;
signal \N__30210\ : std_logic;
signal \N__30203\ : std_logic;
signal \N__30202\ : std_logic;
signal \N__30199\ : std_logic;
signal \N__30198\ : std_logic;
signal \N__30195\ : std_logic;
signal \N__30194\ : std_logic;
signal \N__30191\ : std_logic;
signal \N__30188\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30184\ : std_logic;
signal \N__30181\ : std_logic;
signal \N__30178\ : std_logic;
signal \N__30175\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30169\ : std_logic;
signal \N__30164\ : std_logic;
signal \N__30161\ : std_logic;
signal \N__30152\ : std_logic;
signal \N__30149\ : std_logic;
signal \N__30146\ : std_logic;
signal \N__30143\ : std_logic;
signal \N__30140\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30134\ : std_logic;
signal \N__30131\ : std_logic;
signal \N__30128\ : std_logic;
signal \N__30125\ : std_logic;
signal \N__30124\ : std_logic;
signal \N__30121\ : std_logic;
signal \N__30118\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30116\ : std_logic;
signal \N__30113\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30105\ : std_logic;
signal \N__30104\ : std_logic;
signal \N__30101\ : std_logic;
signal \N__30096\ : std_logic;
signal \N__30093\ : std_logic;
signal \N__30086\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30082\ : std_logic;
signal \N__30079\ : std_logic;
signal \N__30076\ : std_logic;
signal \N__30075\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30068\ : std_logic;
signal \N__30065\ : std_logic;
signal \N__30060\ : std_logic;
signal \N__30057\ : std_logic;
signal \N__30054\ : std_logic;
signal \N__30047\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30041\ : std_logic;
signal \N__30040\ : std_logic;
signal \N__30037\ : std_logic;
signal \N__30034\ : std_logic;
signal \N__30031\ : std_logic;
signal \N__30028\ : std_logic;
signal \N__30025\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30015\ : std_logic;
signal \N__30008\ : std_logic;
signal \N__30005\ : std_logic;
signal \N__30002\ : std_logic;
signal \N__29999\ : std_logic;
signal \N__29996\ : std_logic;
signal \N__29993\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29987\ : std_logic;
signal \N__29984\ : std_logic;
signal \N__29981\ : std_logic;
signal \N__29978\ : std_logic;
signal \N__29975\ : std_logic;
signal \N__29972\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29968\ : std_logic;
signal \N__29965\ : std_logic;
signal \N__29962\ : std_logic;
signal \N__29959\ : std_logic;
signal \N__29956\ : std_logic;
signal \N__29953\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29947\ : std_logic;
signal \N__29944\ : std_logic;
signal \N__29941\ : std_logic;
signal \N__29938\ : std_logic;
signal \N__29933\ : std_logic;
signal \N__29930\ : std_logic;
signal \N__29927\ : std_logic;
signal \N__29924\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29918\ : std_logic;
signal \N__29915\ : std_logic;
signal \N__29912\ : std_logic;
signal \N__29909\ : std_logic;
signal \N__29906\ : std_logic;
signal \N__29903\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29897\ : std_logic;
signal \N__29894\ : std_logic;
signal \N__29891\ : std_logic;
signal \N__29888\ : std_logic;
signal \N__29885\ : std_logic;
signal \N__29882\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29876\ : std_logic;
signal \N__29873\ : std_logic;
signal \N__29870\ : std_logic;
signal \N__29867\ : std_logic;
signal \N__29864\ : std_logic;
signal \N__29861\ : std_logic;
signal \N__29858\ : std_logic;
signal \N__29855\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29849\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29843\ : std_logic;
signal \N__29840\ : std_logic;
signal \N__29837\ : std_logic;
signal \N__29834\ : std_logic;
signal \N__29831\ : std_logic;
signal \N__29828\ : std_logic;
signal \N__29825\ : std_logic;
signal \N__29822\ : std_logic;
signal \N__29819\ : std_logic;
signal \N__29816\ : std_logic;
signal \N__29813\ : std_logic;
signal \N__29810\ : std_logic;
signal \N__29807\ : std_logic;
signal \N__29804\ : std_logic;
signal \N__29801\ : std_logic;
signal \N__29798\ : std_logic;
signal \N__29795\ : std_logic;
signal \N__29792\ : std_logic;
signal \N__29789\ : std_logic;
signal \N__29786\ : std_logic;
signal \N__29783\ : std_logic;
signal \N__29780\ : std_logic;
signal \N__29777\ : std_logic;
signal \N__29774\ : std_logic;
signal \N__29771\ : std_logic;
signal \N__29768\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29764\ : std_logic;
signal \N__29763\ : std_logic;
signal \N__29760\ : std_logic;
signal \N__29757\ : std_logic;
signal \N__29754\ : std_logic;
signal \N__29751\ : std_logic;
signal \N__29748\ : std_logic;
signal \N__29741\ : std_logic;
signal \N__29738\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29729\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29723\ : std_logic;
signal \N__29720\ : std_logic;
signal \N__29717\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29708\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29704\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29695\ : std_logic;
signal \N__29694\ : std_logic;
signal \N__29693\ : std_logic;
signal \N__29690\ : std_logic;
signal \N__29687\ : std_logic;
signal \N__29684\ : std_logic;
signal \N__29681\ : std_logic;
signal \N__29678\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29672\ : std_logic;
signal \N__29669\ : std_logic;
signal \N__29666\ : std_logic;
signal \N__29659\ : std_logic;
signal \N__29654\ : std_logic;
signal \N__29651\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29645\ : std_logic;
signal \N__29642\ : std_logic;
signal \N__29639\ : std_logic;
signal \N__29636\ : std_logic;
signal \N__29633\ : std_logic;
signal \N__29632\ : std_logic;
signal \N__29631\ : std_logic;
signal \N__29628\ : std_logic;
signal \N__29625\ : std_logic;
signal \N__29622\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29616\ : std_logic;
signal \N__29615\ : std_logic;
signal \N__29612\ : std_logic;
signal \N__29607\ : std_logic;
signal \N__29604\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29588\ : std_logic;
signal \N__29585\ : std_logic;
signal \N__29582\ : std_logic;
signal \N__29579\ : std_logic;
signal \N__29576\ : std_logic;
signal \N__29575\ : std_logic;
signal \N__29572\ : std_logic;
signal \N__29569\ : std_logic;
signal \N__29568\ : std_logic;
signal \N__29565\ : std_logic;
signal \N__29562\ : std_logic;
signal \N__29561\ : std_logic;
signal \N__29558\ : std_logic;
signal \N__29555\ : std_logic;
signal \N__29552\ : std_logic;
signal \N__29549\ : std_logic;
signal \N__29546\ : std_logic;
signal \N__29543\ : std_logic;
signal \N__29538\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29528\ : std_logic;
signal \N__29525\ : std_logic;
signal \N__29522\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29516\ : std_logic;
signal \N__29513\ : std_logic;
signal \N__29510\ : std_logic;
signal \N__29509\ : std_logic;
signal \N__29508\ : std_logic;
signal \N__29507\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29503\ : std_logic;
signal \N__29500\ : std_logic;
signal \N__29499\ : std_logic;
signal \N__29496\ : std_logic;
signal \N__29495\ : std_logic;
signal \N__29492\ : std_logic;
signal \N__29491\ : std_logic;
signal \N__29488\ : std_logic;
signal \N__29485\ : std_logic;
signal \N__29470\ : std_logic;
signal \N__29467\ : std_logic;
signal \N__29464\ : std_logic;
signal \N__29461\ : std_logic;
signal \N__29458\ : std_logic;
signal \N__29453\ : std_logic;
signal \N__29450\ : std_logic;
signal \N__29447\ : std_logic;
signal \N__29446\ : std_logic;
signal \N__29443\ : std_logic;
signal \N__29440\ : std_logic;
signal \N__29437\ : std_logic;
signal \N__29434\ : std_logic;
signal \N__29431\ : std_logic;
signal \N__29428\ : std_logic;
signal \N__29423\ : std_logic;
signal \N__29422\ : std_logic;
signal \N__29419\ : std_logic;
signal \N__29418\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29414\ : std_logic;
signal \N__29411\ : std_logic;
signal \N__29408\ : std_logic;
signal \N__29405\ : std_logic;
signal \N__29402\ : std_logic;
signal \N__29395\ : std_logic;
signal \N__29392\ : std_logic;
signal \N__29389\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29378\ : std_logic;
signal \N__29375\ : std_logic;
signal \N__29372\ : std_logic;
signal \N__29369\ : std_logic;
signal \N__29366\ : std_logic;
signal \N__29363\ : std_logic;
signal \N__29360\ : std_logic;
signal \N__29357\ : std_logic;
signal \N__29356\ : std_logic;
signal \N__29355\ : std_logic;
signal \N__29354\ : std_logic;
signal \N__29351\ : std_logic;
signal \N__29348\ : std_logic;
signal \N__29343\ : std_logic;
signal \N__29336\ : std_logic;
signal \N__29335\ : std_logic;
signal \N__29332\ : std_logic;
signal \N__29329\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29323\ : std_logic;
signal \N__29320\ : std_logic;
signal \N__29317\ : std_logic;
signal \N__29314\ : std_logic;
signal \N__29309\ : std_logic;
signal \N__29306\ : std_logic;
signal \N__29303\ : std_logic;
signal \N__29300\ : std_logic;
signal \N__29297\ : std_logic;
signal \N__29296\ : std_logic;
signal \N__29293\ : std_logic;
signal \N__29292\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29282\ : std_logic;
signal \N__29279\ : std_logic;
signal \N__29274\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29265\ : std_logic;
signal \N__29258\ : std_logic;
signal \N__29257\ : std_logic;
signal \N__29254\ : std_logic;
signal \N__29251\ : std_logic;
signal \N__29248\ : std_logic;
signal \N__29245\ : std_logic;
signal \N__29242\ : std_logic;
signal \N__29237\ : std_logic;
signal \N__29234\ : std_logic;
signal \N__29231\ : std_logic;
signal \N__29228\ : std_logic;
signal \N__29225\ : std_logic;
signal \N__29222\ : std_logic;
signal \N__29219\ : std_logic;
signal \N__29218\ : std_logic;
signal \N__29217\ : std_logic;
signal \N__29216\ : std_logic;
signal \N__29213\ : std_logic;
signal \N__29210\ : std_logic;
signal \N__29207\ : std_logic;
signal \N__29204\ : std_logic;
signal \N__29201\ : std_logic;
signal \N__29198\ : std_logic;
signal \N__29193\ : std_logic;
signal \N__29186\ : std_logic;
signal \N__29185\ : std_logic;
signal \N__29182\ : std_logic;
signal \N__29179\ : std_logic;
signal \N__29176\ : std_logic;
signal \N__29173\ : std_logic;
signal \N__29170\ : std_logic;
signal \N__29165\ : std_logic;
signal \N__29162\ : std_logic;
signal \N__29159\ : std_logic;
signal \N__29156\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29150\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29146\ : std_logic;
signal \N__29143\ : std_logic;
signal \N__29140\ : std_logic;
signal \N__29137\ : std_logic;
signal \N__29134\ : std_logic;
signal \N__29131\ : std_logic;
signal \N__29128\ : std_logic;
signal \N__29125\ : std_logic;
signal \N__29120\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29111\ : std_logic;
signal \N__29108\ : std_logic;
signal \N__29107\ : std_logic;
signal \N__29104\ : std_logic;
signal \N__29101\ : std_logic;
signal \N__29100\ : std_logic;
signal \N__29097\ : std_logic;
signal \N__29094\ : std_logic;
signal \N__29093\ : std_logic;
signal \N__29090\ : std_logic;
signal \N__29087\ : std_logic;
signal \N__29084\ : std_logic;
signal \N__29079\ : std_logic;
signal \N__29072\ : std_logic;
signal \N__29069\ : std_logic;
signal \N__29066\ : std_logic;
signal \N__29063\ : std_logic;
signal \N__29060\ : std_logic;
signal \N__29057\ : std_logic;
signal \N__29056\ : std_logic;
signal \N__29053\ : std_logic;
signal \N__29050\ : std_logic;
signal \N__29047\ : std_logic;
signal \N__29046\ : std_logic;
signal \N__29045\ : std_logic;
signal \N__29042\ : std_logic;
signal \N__29039\ : std_logic;
signal \N__29036\ : std_logic;
signal \N__29033\ : std_logic;
signal \N__29024\ : std_logic;
signal \N__29023\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__29017\ : std_logic;
signal \N__29014\ : std_logic;
signal \N__29011\ : std_logic;
signal \N__29008\ : std_logic;
signal \N__29005\ : std_logic;
signal \N__29002\ : std_logic;
signal \N__28997\ : std_logic;
signal \N__28994\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28988\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28984\ : std_logic;
signal \N__28981\ : std_logic;
signal \N__28980\ : std_logic;
signal \N__28979\ : std_logic;
signal \N__28976\ : std_logic;
signal \N__28973\ : std_logic;
signal \N__28970\ : std_logic;
signal \N__28967\ : std_logic;
signal \N__28964\ : std_logic;
signal \N__28955\ : std_logic;
signal \N__28952\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28948\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28939\ : std_logic;
signal \N__28936\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28925\ : std_logic;
signal \N__28922\ : std_logic;
signal \N__28919\ : std_logic;
signal \N__28916\ : std_logic;
signal \N__28913\ : std_logic;
signal \N__28910\ : std_logic;
signal \N__28907\ : std_logic;
signal \N__28906\ : std_logic;
signal \N__28903\ : std_logic;
signal \N__28902\ : std_logic;
signal \N__28901\ : std_logic;
signal \N__28898\ : std_logic;
signal \N__28895\ : std_logic;
signal \N__28892\ : std_logic;
signal \N__28889\ : std_logic;
signal \N__28886\ : std_logic;
signal \N__28877\ : std_logic;
signal \N__28876\ : std_logic;
signal \N__28873\ : std_logic;
signal \N__28870\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28864\ : std_logic;
signal \N__28861\ : std_logic;
signal \N__28856\ : std_logic;
signal \N__28853\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28847\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28837\ : std_logic;
signal \N__28834\ : std_logic;
signal \N__28833\ : std_logic;
signal \N__28830\ : std_logic;
signal \N__28827\ : std_logic;
signal \N__28826\ : std_logic;
signal \N__28823\ : std_logic;
signal \N__28820\ : std_logic;
signal \N__28817\ : std_logic;
signal \N__28814\ : std_logic;
signal \N__28809\ : std_logic;
signal \N__28806\ : std_logic;
signal \N__28803\ : std_logic;
signal \N__28800\ : std_logic;
signal \N__28793\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28786\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28780\ : std_logic;
signal \N__28777\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28771\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28763\ : std_logic;
signal \N__28760\ : std_logic;
signal \N__28757\ : std_logic;
signal \N__28754\ : std_logic;
signal \N__28751\ : std_logic;
signal \N__28748\ : std_logic;
signal \N__28747\ : std_logic;
signal \N__28744\ : std_logic;
signal \N__28743\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28737\ : std_logic;
signal \N__28736\ : std_logic;
signal \N__28733\ : std_logic;
signal \N__28730\ : std_logic;
signal \N__28727\ : std_logic;
signal \N__28724\ : std_logic;
signal \N__28719\ : std_logic;
signal \N__28712\ : std_logic;
signal \N__28709\ : std_logic;
signal \N__28708\ : std_logic;
signal \N__28705\ : std_logic;
signal \N__28702\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28696\ : std_logic;
signal \N__28693\ : std_logic;
signal \N__28688\ : std_logic;
signal \N__28685\ : std_logic;
signal \N__28682\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28676\ : std_logic;
signal \N__28673\ : std_logic;
signal \N__28670\ : std_logic;
signal \N__28667\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28660\ : std_logic;
signal \N__28659\ : std_logic;
signal \N__28656\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28652\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28643\ : std_logic;
signal \N__28634\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28630\ : std_logic;
signal \N__28627\ : std_logic;
signal \N__28624\ : std_logic;
signal \N__28621\ : std_logic;
signal \N__28618\ : std_logic;
signal \N__28615\ : std_logic;
signal \N__28612\ : std_logic;
signal \N__28607\ : std_logic;
signal \N__28604\ : std_logic;
signal \N__28601\ : std_logic;
signal \N__28598\ : std_logic;
signal \N__28595\ : std_logic;
signal \N__28592\ : std_logic;
signal \N__28591\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28587\ : std_logic;
signal \N__28584\ : std_logic;
signal \N__28583\ : std_logic;
signal \N__28580\ : std_logic;
signal \N__28577\ : std_logic;
signal \N__28574\ : std_logic;
signal \N__28571\ : std_logic;
signal \N__28568\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28556\ : std_logic;
signal \N__28555\ : std_logic;
signal \N__28552\ : std_logic;
signal \N__28549\ : std_logic;
signal \N__28546\ : std_logic;
signal \N__28543\ : std_logic;
signal \N__28540\ : std_logic;
signal \N__28537\ : std_logic;
signal \N__28534\ : std_logic;
signal \N__28529\ : std_logic;
signal \N__28526\ : std_logic;
signal \N__28523\ : std_logic;
signal \N__28520\ : std_logic;
signal \N__28517\ : std_logic;
signal \N__28514\ : std_logic;
signal \N__28511\ : std_logic;
signal \N__28510\ : std_logic;
signal \N__28509\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28505\ : std_logic;
signal \N__28500\ : std_logic;
signal \N__28497\ : std_logic;
signal \N__28494\ : std_logic;
signal \N__28491\ : std_logic;
signal \N__28484\ : std_logic;
signal \N__28483\ : std_logic;
signal \N__28480\ : std_logic;
signal \N__28477\ : std_logic;
signal \N__28474\ : std_logic;
signal \N__28471\ : std_logic;
signal \N__28468\ : std_logic;
signal \N__28465\ : std_logic;
signal \N__28462\ : std_logic;
signal \N__28457\ : std_logic;
signal \N__28454\ : std_logic;
signal \N__28451\ : std_logic;
signal \N__28448\ : std_logic;
signal \N__28445\ : std_logic;
signal \N__28442\ : std_logic;
signal \N__28441\ : std_logic;
signal \N__28440\ : std_logic;
signal \N__28437\ : std_logic;
signal \N__28434\ : std_logic;
signal \N__28431\ : std_logic;
signal \N__28424\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28420\ : std_logic;
signal \N__28417\ : std_logic;
signal \N__28412\ : std_logic;
signal \N__28411\ : std_logic;
signal \N__28408\ : std_logic;
signal \N__28405\ : std_logic;
signal \N__28402\ : std_logic;
signal \N__28399\ : std_logic;
signal \N__28396\ : std_logic;
signal \N__28393\ : std_logic;
signal \N__28388\ : std_logic;
signal \N__28385\ : std_logic;
signal \N__28382\ : std_logic;
signal \N__28379\ : std_logic;
signal \N__28376\ : std_logic;
signal \N__28373\ : std_logic;
signal \N__28370\ : std_logic;
signal \N__28367\ : std_logic;
signal \N__28366\ : std_logic;
signal \N__28365\ : std_logic;
signal \N__28362\ : std_logic;
signal \N__28361\ : std_logic;
signal \N__28356\ : std_logic;
signal \N__28353\ : std_logic;
signal \N__28350\ : std_logic;
signal \N__28347\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28339\ : std_logic;
signal \N__28336\ : std_logic;
signal \N__28333\ : std_logic;
signal \N__28330\ : std_logic;
signal \N__28327\ : std_logic;
signal \N__28324\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28316\ : std_logic;
signal \N__28313\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28307\ : std_logic;
signal \N__28304\ : std_logic;
signal \N__28303\ : std_logic;
signal \N__28300\ : std_logic;
signal \N__28297\ : std_logic;
signal \N__28296\ : std_logic;
signal \N__28293\ : std_logic;
signal \N__28290\ : std_logic;
signal \N__28287\ : std_logic;
signal \N__28286\ : std_logic;
signal \N__28281\ : std_logic;
signal \N__28278\ : std_logic;
signal \N__28275\ : std_logic;
signal \N__28270\ : std_logic;
signal \N__28265\ : std_logic;
signal \N__28262\ : std_logic;
signal \N__28261\ : std_logic;
signal \N__28258\ : std_logic;
signal \N__28255\ : std_logic;
signal \N__28252\ : std_logic;
signal \N__28249\ : std_logic;
signal \N__28246\ : std_logic;
signal \N__28243\ : std_logic;
signal \N__28240\ : std_logic;
signal \N__28237\ : std_logic;
signal \N__28232\ : std_logic;
signal \N__28229\ : std_logic;
signal \N__28226\ : std_logic;
signal \N__28223\ : std_logic;
signal \N__28220\ : std_logic;
signal \N__28219\ : std_logic;
signal \N__28216\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28212\ : std_logic;
signal \N__28209\ : std_logic;
signal \N__28206\ : std_logic;
signal \N__28203\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28195\ : std_logic;
signal \N__28192\ : std_logic;
signal \N__28189\ : std_logic;
signal \N__28184\ : std_logic;
signal \N__28183\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28177\ : std_logic;
signal \N__28174\ : std_logic;
signal \N__28171\ : std_logic;
signal \N__28168\ : std_logic;
signal \N__28165\ : std_logic;
signal \N__28160\ : std_logic;
signal \N__28157\ : std_logic;
signal \N__28154\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28144\ : std_logic;
signal \N__28141\ : std_logic;
signal \N__28138\ : std_logic;
signal \N__28135\ : std_logic;
signal \N__28134\ : std_logic;
signal \N__28133\ : std_logic;
signal \N__28130\ : std_logic;
signal \N__28127\ : std_logic;
signal \N__28124\ : std_logic;
signal \N__28121\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28109\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28099\ : std_logic;
signal \N__28096\ : std_logic;
signal \N__28093\ : std_logic;
signal \N__28090\ : std_logic;
signal \N__28087\ : std_logic;
signal \N__28082\ : std_logic;
signal \N__28079\ : std_logic;
signal \N__28076\ : std_logic;
signal \N__28073\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28069\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28063\ : std_logic;
signal \N__28060\ : std_logic;
signal \N__28057\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28051\ : std_logic;
signal \N__28050\ : std_logic;
signal \N__28047\ : std_logic;
signal \N__28044\ : std_logic;
signal \N__28041\ : std_logic;
signal \N__28034\ : std_logic;
signal \N__28031\ : std_logic;
signal \N__28030\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28024\ : std_logic;
signal \N__28021\ : std_logic;
signal \N__28018\ : std_logic;
signal \N__28015\ : std_logic;
signal \N__28012\ : std_logic;
signal \N__28009\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__27998\ : std_logic;
signal \N__27995\ : std_logic;
signal \N__27992\ : std_logic;
signal \N__27991\ : std_logic;
signal \N__27988\ : std_logic;
signal \N__27985\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27978\ : std_logic;
signal \N__27975\ : std_logic;
signal \N__27972\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27964\ : std_logic;
signal \N__27961\ : std_logic;
signal \N__27958\ : std_logic;
signal \N__27955\ : std_logic;
signal \N__27952\ : std_logic;
signal \N__27949\ : std_logic;
signal \N__27946\ : std_logic;
signal \N__27941\ : std_logic;
signal \N__27938\ : std_logic;
signal \N__27935\ : std_logic;
signal \N__27932\ : std_logic;
signal \N__27929\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27922\ : std_logic;
signal \N__27919\ : std_logic;
signal \N__27918\ : std_logic;
signal \N__27915\ : std_logic;
signal \N__27912\ : std_logic;
signal \N__27909\ : std_logic;
signal \N__27906\ : std_logic;
signal \N__27899\ : std_logic;
signal \N__27896\ : std_logic;
signal \N__27895\ : std_logic;
signal \N__27892\ : std_logic;
signal \N__27889\ : std_logic;
signal \N__27886\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27880\ : std_logic;
signal \N__27875\ : std_logic;
signal \N__27872\ : std_logic;
signal \N__27869\ : std_logic;
signal \N__27866\ : std_logic;
signal \N__27863\ : std_logic;
signal \N__27860\ : std_logic;
signal \N__27859\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27853\ : std_logic;
signal \N__27850\ : std_logic;
signal \N__27847\ : std_logic;
signal \N__27844\ : std_logic;
signal \N__27839\ : std_logic;
signal \N__27836\ : std_logic;
signal \N__27833\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27829\ : std_logic;
signal \N__27826\ : std_logic;
signal \N__27823\ : std_logic;
signal \N__27820\ : std_logic;
signal \N__27817\ : std_logic;
signal \N__27814\ : std_logic;
signal \N__27809\ : std_logic;
signal \N__27806\ : std_logic;
signal \N__27805\ : std_logic;
signal \N__27804\ : std_logic;
signal \N__27803\ : std_logic;
signal \N__27800\ : std_logic;
signal \N__27797\ : std_logic;
signal \N__27794\ : std_logic;
signal \N__27791\ : std_logic;
signal \N__27784\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27773\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27764\ : std_logic;
signal \N__27761\ : std_logic;
signal \N__27760\ : std_logic;
signal \N__27755\ : std_logic;
signal \N__27754\ : std_logic;
signal \N__27751\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27744\ : std_logic;
signal \N__27741\ : std_logic;
signal \N__27738\ : std_logic;
signal \N__27735\ : std_logic;
signal \N__27728\ : std_logic;
signal \N__27725\ : std_logic;
signal \N__27722\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27718\ : std_logic;
signal \N__27715\ : std_logic;
signal \N__27712\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27701\ : std_logic;
signal \N__27698\ : std_logic;
signal \N__27695\ : std_logic;
signal \N__27692\ : std_logic;
signal \N__27691\ : std_logic;
signal \N__27690\ : std_logic;
signal \N__27687\ : std_logic;
signal \N__27684\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27678\ : std_logic;
signal \N__27677\ : std_logic;
signal \N__27672\ : std_logic;
signal \N__27669\ : std_logic;
signal \N__27666\ : std_logic;
signal \N__27663\ : std_logic;
signal \N__27656\ : std_logic;
signal \N__27655\ : std_logic;
signal \N__27652\ : std_logic;
signal \N__27649\ : std_logic;
signal \N__27646\ : std_logic;
signal \N__27643\ : std_logic;
signal \N__27640\ : std_logic;
signal \N__27637\ : std_logic;
signal \N__27634\ : std_logic;
signal \N__27631\ : std_logic;
signal \N__27626\ : std_logic;
signal \N__27623\ : std_logic;
signal \N__27620\ : std_logic;
signal \N__27617\ : std_logic;
signal \N__27614\ : std_logic;
signal \N__27613\ : std_logic;
signal \N__27612\ : std_logic;
signal \N__27609\ : std_logic;
signal \N__27606\ : std_logic;
signal \N__27603\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27601\ : std_logic;
signal \N__27598\ : std_logic;
signal \N__27595\ : std_logic;
signal \N__27590\ : std_logic;
signal \N__27587\ : std_logic;
signal \N__27584\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27572\ : std_logic;
signal \N__27569\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27567\ : std_logic;
signal \N__27564\ : std_logic;
signal \N__27563\ : std_logic;
signal \N__27560\ : std_logic;
signal \N__27557\ : std_logic;
signal \N__27554\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27541\ : std_logic;
signal \N__27540\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27533\ : std_logic;
signal \N__27530\ : std_logic;
signal \N__27527\ : std_logic;
signal \N__27518\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27511\ : std_logic;
signal \N__27508\ : std_logic;
signal \N__27507\ : std_logic;
signal \N__27506\ : std_logic;
signal \N__27503\ : std_logic;
signal \N__27500\ : std_logic;
signal \N__27497\ : std_logic;
signal \N__27494\ : std_logic;
signal \N__27491\ : std_logic;
signal \N__27488\ : std_logic;
signal \N__27485\ : std_logic;
signal \N__27482\ : std_logic;
signal \N__27473\ : std_logic;
signal \N__27472\ : std_logic;
signal \N__27471\ : std_logic;
signal \N__27470\ : std_logic;
signal \N__27467\ : std_logic;
signal \N__27462\ : std_logic;
signal \N__27459\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27451\ : std_logic;
signal \N__27450\ : std_logic;
signal \N__27447\ : std_logic;
signal \N__27446\ : std_logic;
signal \N__27443\ : std_logic;
signal \N__27440\ : std_logic;
signal \N__27437\ : std_logic;
signal \N__27434\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27419\ : std_logic;
signal \N__27416\ : std_logic;
signal \N__27413\ : std_logic;
signal \N__27410\ : std_logic;
signal \N__27407\ : std_logic;
signal \N__27404\ : std_logic;
signal \N__27401\ : std_logic;
signal \N__27398\ : std_logic;
signal \N__27395\ : std_logic;
signal \N__27392\ : std_logic;
signal \N__27389\ : std_logic;
signal \N__27386\ : std_logic;
signal \N__27383\ : std_logic;
signal \N__27380\ : std_logic;
signal \N__27377\ : std_logic;
signal \N__27374\ : std_logic;
signal \N__27371\ : std_logic;
signal \N__27368\ : std_logic;
signal \N__27365\ : std_logic;
signal \N__27362\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27358\ : std_logic;
signal \N__27357\ : std_logic;
signal \N__27356\ : std_logic;
signal \N__27355\ : std_logic;
signal \N__27354\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27352\ : std_logic;
signal \N__27351\ : std_logic;
signal \N__27350\ : std_logic;
signal \N__27349\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27346\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27344\ : std_logic;
signal \N__27343\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27341\ : std_logic;
signal \N__27340\ : std_logic;
signal \N__27339\ : std_logic;
signal \N__27338\ : std_logic;
signal \N__27337\ : std_logic;
signal \N__27336\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27334\ : std_logic;
signal \N__27333\ : std_logic;
signal \N__27332\ : std_logic;
signal \N__27331\ : std_logic;
signal \N__27330\ : std_logic;
signal \N__27325\ : std_logic;
signal \N__27316\ : std_logic;
signal \N__27307\ : std_logic;
signal \N__27298\ : std_logic;
signal \N__27289\ : std_logic;
signal \N__27280\ : std_logic;
signal \N__27271\ : std_logic;
signal \N__27262\ : std_logic;
signal \N__27255\ : std_logic;
signal \N__27242\ : std_logic;
signal \N__27239\ : std_logic;
signal \N__27236\ : std_logic;
signal \N__27233\ : std_logic;
signal \N__27230\ : std_logic;
signal \N__27227\ : std_logic;
signal \N__27224\ : std_logic;
signal \N__27221\ : std_logic;
signal \N__27218\ : std_logic;
signal \N__27215\ : std_logic;
signal \N__27212\ : std_logic;
signal \N__27209\ : std_logic;
signal \N__27206\ : std_logic;
signal \N__27203\ : std_logic;
signal \N__27200\ : std_logic;
signal \N__27197\ : std_logic;
signal \N__27194\ : std_logic;
signal \N__27191\ : std_logic;
signal \N__27188\ : std_logic;
signal \N__27185\ : std_logic;
signal \N__27182\ : std_logic;
signal \N__27179\ : std_logic;
signal \N__27176\ : std_logic;
signal \N__27173\ : std_logic;
signal \N__27170\ : std_logic;
signal \N__27169\ : std_logic;
signal \N__27164\ : std_logic;
signal \N__27161\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27157\ : std_logic;
signal \N__27154\ : std_logic;
signal \N__27149\ : std_logic;
signal \N__27146\ : std_logic;
signal \N__27143\ : std_logic;
signal \N__27142\ : std_logic;
signal \N__27139\ : std_logic;
signal \N__27136\ : std_logic;
signal \N__27135\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27133\ : std_logic;
signal \N__27132\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27112\ : std_logic;
signal \N__27109\ : std_logic;
signal \N__27106\ : std_logic;
signal \N__27103\ : std_logic;
signal \N__27100\ : std_logic;
signal \N__27097\ : std_logic;
signal \N__27094\ : std_logic;
signal \N__27087\ : std_logic;
signal \N__27082\ : std_logic;
signal \N__27079\ : std_logic;
signal \N__27068\ : std_logic;
signal \N__27065\ : std_logic;
signal \N__27064\ : std_logic;
signal \N__27059\ : std_logic;
signal \N__27056\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27052\ : std_logic;
signal \N__27049\ : std_logic;
signal \N__27044\ : std_logic;
signal \N__27043\ : std_logic;
signal \N__27042\ : std_logic;
signal \N__27039\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27033\ : std_logic;
signal \N__27030\ : std_logic;
signal \N__27027\ : std_logic;
signal \N__27024\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27011\ : std_logic;
signal \N__27008\ : std_logic;
signal \N__27007\ : std_logic;
signal \N__27002\ : std_logic;
signal \N__27001\ : std_logic;
signal \N__27000\ : std_logic;
signal \N__26997\ : std_logic;
signal \N__26994\ : std_logic;
signal \N__26991\ : std_logic;
signal \N__26988\ : std_logic;
signal \N__26985\ : std_logic;
signal \N__26978\ : std_logic;
signal \N__26975\ : std_logic;
signal \N__26972\ : std_logic;
signal \N__26969\ : std_logic;
signal \N__26966\ : std_logic;
signal \N__26963\ : std_logic;
signal \N__26960\ : std_logic;
signal \N__26959\ : std_logic;
signal \N__26956\ : std_logic;
signal \N__26953\ : std_logic;
signal \N__26952\ : std_logic;
signal \N__26951\ : std_logic;
signal \N__26948\ : std_logic;
signal \N__26943\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26924\ : std_logic;
signal \N__26921\ : std_logic;
signal \N__26918\ : std_logic;
signal \N__26915\ : std_logic;
signal \N__26914\ : std_logic;
signal \N__26913\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26909\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26896\ : std_logic;
signal \N__26893\ : std_logic;
signal \N__26888\ : std_logic;
signal \N__26885\ : std_logic;
signal \N__26882\ : std_logic;
signal \N__26879\ : std_logic;
signal \N__26878\ : std_logic;
signal \N__26877\ : std_logic;
signal \N__26874\ : std_logic;
signal \N__26869\ : std_logic;
signal \N__26868\ : std_logic;
signal \N__26863\ : std_logic;
signal \N__26860\ : std_logic;
signal \N__26857\ : std_logic;
signal \N__26854\ : std_logic;
signal \N__26849\ : std_logic;
signal \N__26846\ : std_logic;
signal \N__26843\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26841\ : std_logic;
signal \N__26840\ : std_logic;
signal \N__26837\ : std_logic;
signal \N__26832\ : std_logic;
signal \N__26829\ : std_logic;
signal \N__26824\ : std_logic;
signal \N__26821\ : std_logic;
signal \N__26816\ : std_logic;
signal \N__26813\ : std_logic;
signal \N__26812\ : std_logic;
signal \N__26807\ : std_logic;
signal \N__26806\ : std_logic;
signal \N__26803\ : std_logic;
signal \N__26800\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26794\ : std_logic;
signal \N__26791\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26783\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26774\ : std_logic;
signal \N__26771\ : std_logic;
signal \N__26770\ : std_logic;
signal \N__26769\ : std_logic;
signal \N__26766\ : std_logic;
signal \N__26765\ : std_logic;
signal \N__26760\ : std_logic;
signal \N__26757\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26748\ : std_logic;
signal \N__26745\ : std_logic;
signal \N__26738\ : std_logic;
signal \N__26735\ : std_logic;
signal \N__26734\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26730\ : std_logic;
signal \N__26727\ : std_logic;
signal \N__26724\ : std_logic;
signal \N__26721\ : std_logic;
signal \N__26720\ : std_logic;
signal \N__26715\ : std_logic;
signal \N__26712\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26704\ : std_logic;
signal \N__26701\ : std_logic;
signal \N__26696\ : std_logic;
signal \N__26693\ : std_logic;
signal \N__26690\ : std_logic;
signal \N__26689\ : std_logic;
signal \N__26688\ : std_logic;
signal \N__26685\ : std_logic;
signal \N__26682\ : std_logic;
signal \N__26681\ : std_logic;
signal \N__26678\ : std_logic;
signal \N__26673\ : std_logic;
signal \N__26670\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26662\ : std_logic;
signal \N__26657\ : std_logic;
signal \N__26654\ : std_logic;
signal \N__26651\ : std_logic;
signal \N__26648\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26643\ : std_logic;
signal \N__26640\ : std_logic;
signal \N__26635\ : std_logic;
signal \N__26634\ : std_logic;
signal \N__26631\ : std_logic;
signal \N__26628\ : std_logic;
signal \N__26625\ : std_logic;
signal \N__26622\ : std_logic;
signal \N__26619\ : std_logic;
signal \N__26616\ : std_logic;
signal \N__26609\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26600\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26598\ : std_logic;
signal \N__26597\ : std_logic;
signal \N__26594\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26588\ : std_logic;
signal \N__26585\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26570\ : std_logic;
signal \N__26567\ : std_logic;
signal \N__26566\ : std_logic;
signal \N__26565\ : std_logic;
signal \N__26562\ : std_logic;
signal \N__26557\ : std_logic;
signal \N__26556\ : std_logic;
signal \N__26551\ : std_logic;
signal \N__26548\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26539\ : std_logic;
signal \N__26538\ : std_logic;
signal \N__26535\ : std_logic;
signal \N__26530\ : std_logic;
signal \N__26525\ : std_logic;
signal \N__26524\ : std_logic;
signal \N__26521\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26513\ : std_logic;
signal \N__26510\ : std_logic;
signal \N__26507\ : std_logic;
signal \N__26504\ : std_logic;
signal \N__26501\ : std_logic;
signal \N__26500\ : std_logic;
signal \N__26497\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26489\ : std_logic;
signal \N__26488\ : std_logic;
signal \N__26485\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26479\ : std_logic;
signal \N__26476\ : std_logic;
signal \N__26475\ : std_logic;
signal \N__26472\ : std_logic;
signal \N__26469\ : std_logic;
signal \N__26466\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26452\ : std_logic;
signal \N__26449\ : std_logic;
signal \N__26448\ : std_logic;
signal \N__26445\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26439\ : std_logic;
signal \N__26436\ : std_logic;
signal \N__26433\ : std_logic;
signal \N__26430\ : std_logic;
signal \N__26423\ : std_logic;
signal \N__26420\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26414\ : std_logic;
signal \N__26413\ : std_logic;
signal \N__26410\ : std_logic;
signal \N__26407\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26398\ : std_logic;
signal \N__26397\ : std_logic;
signal \N__26394\ : std_logic;
signal \N__26389\ : std_logic;
signal \N__26388\ : std_logic;
signal \N__26383\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26369\ : std_logic;
signal \N__26368\ : std_logic;
signal \N__26367\ : std_logic;
signal \N__26366\ : std_logic;
signal \N__26359\ : std_logic;
signal \N__26356\ : std_logic;
signal \N__26353\ : std_logic;
signal \N__26350\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26342\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26338\ : std_logic;
signal \N__26337\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26331\ : std_logic;
signal \N__26328\ : std_logic;
signal \N__26325\ : std_logic;
signal \N__26320\ : std_logic;
signal \N__26317\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26306\ : std_logic;
signal \N__26305\ : std_logic;
signal \N__26304\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26300\ : std_logic;
signal \N__26295\ : std_logic;
signal \N__26292\ : std_logic;
signal \N__26287\ : std_logic;
signal \N__26284\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26261\ : std_logic;
signal \N__26258\ : std_logic;
signal \N__26255\ : std_logic;
signal \N__26252\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26246\ : std_logic;
signal \N__26243\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26239\ : std_logic;
signal \N__26236\ : std_logic;
signal \N__26233\ : std_logic;
signal \N__26232\ : std_logic;
signal \N__26229\ : std_logic;
signal \N__26224\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26218\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26212\ : std_logic;
signal \N__26209\ : std_logic;
signal \N__26206\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26198\ : std_logic;
signal \N__26195\ : std_logic;
signal \N__26194\ : std_logic;
signal \N__26189\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26187\ : std_logic;
signal \N__26184\ : std_logic;
signal \N__26181\ : std_logic;
signal \N__26178\ : std_logic;
signal \N__26175\ : std_logic;
signal \N__26172\ : std_logic;
signal \N__26169\ : std_logic;
signal \N__26166\ : std_logic;
signal \N__26161\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26150\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26146\ : std_logic;
signal \N__26141\ : std_logic;
signal \N__26140\ : std_logic;
signal \N__26139\ : std_logic;
signal \N__26136\ : std_logic;
signal \N__26133\ : std_logic;
signal \N__26130\ : std_logic;
signal \N__26127\ : std_logic;
signal \N__26124\ : std_logic;
signal \N__26121\ : std_logic;
signal \N__26118\ : std_logic;
signal \N__26113\ : std_logic;
signal \N__26108\ : std_logic;
signal \N__26105\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26101\ : std_logic;
signal \N__26098\ : std_logic;
signal \N__26097\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26086\ : std_logic;
signal \N__26083\ : std_logic;
signal \N__26080\ : std_logic;
signal \N__26077\ : std_logic;
signal \N__26074\ : std_logic;
signal \N__26069\ : std_logic;
signal \N__26068\ : std_logic;
signal \N__26067\ : std_logic;
signal \N__26062\ : std_logic;
signal \N__26059\ : std_logic;
signal \N__26056\ : std_logic;
signal \N__26053\ : std_logic;
signal \N__26050\ : std_logic;
signal \N__26049\ : std_logic;
signal \N__26044\ : std_logic;
signal \N__26041\ : std_logic;
signal \N__26038\ : std_logic;
signal \N__26035\ : std_logic;
signal \N__26030\ : std_logic;
signal \N__26027\ : std_logic;
signal \N__26024\ : std_logic;
signal \N__26023\ : std_logic;
signal \N__26020\ : std_logic;
signal \N__26019\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26006\ : std_logic;
signal \N__26005\ : std_logic;
signal \N__26002\ : std_logic;
signal \N__25999\ : std_logic;
signal \N__25994\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25990\ : std_logic;
signal \N__25989\ : std_logic;
signal \N__25984\ : std_logic;
signal \N__25981\ : std_logic;
signal \N__25978\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25972\ : std_logic;
signal \N__25971\ : std_logic;
signal \N__25968\ : std_logic;
signal \N__25965\ : std_logic;
signal \N__25962\ : std_logic;
signal \N__25955\ : std_logic;
signal \N__25952\ : std_logic;
signal \N__25949\ : std_logic;
signal \N__25946\ : std_logic;
signal \N__25943\ : std_logic;
signal \N__25940\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25933\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25929\ : std_logic;
signal \N__25926\ : std_logic;
signal \N__25923\ : std_logic;
signal \N__25918\ : std_logic;
signal \N__25915\ : std_logic;
signal \N__25910\ : std_logic;
signal \N__25909\ : std_logic;
signal \N__25906\ : std_logic;
signal \N__25903\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25895\ : std_logic;
signal \N__25892\ : std_logic;
signal \N__25891\ : std_logic;
signal \N__25890\ : std_logic;
signal \N__25887\ : std_logic;
signal \N__25884\ : std_logic;
signal \N__25881\ : std_logic;
signal \N__25880\ : std_logic;
signal \N__25877\ : std_logic;
signal \N__25872\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25863\ : std_logic;
signal \N__25860\ : std_logic;
signal \N__25855\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25847\ : std_logic;
signal \N__25844\ : std_logic;
signal \N__25841\ : std_logic;
signal \N__25838\ : std_logic;
signal \N__25837\ : std_logic;
signal \N__25836\ : std_logic;
signal \N__25833\ : std_logic;
signal \N__25830\ : std_logic;
signal \N__25827\ : std_logic;
signal \N__25826\ : std_logic;
signal \N__25821\ : std_logic;
signal \N__25818\ : std_logic;
signal \N__25815\ : std_logic;
signal \N__25812\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25806\ : std_logic;
signal \N__25803\ : std_logic;
signal \N__25798\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25790\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25781\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25777\ : std_logic;
signal \N__25774\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25770\ : std_logic;
signal \N__25765\ : std_logic;
signal \N__25762\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25753\ : std_logic;
signal \N__25750\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25742\ : std_logic;
signal \N__25741\ : std_logic;
signal \N__25740\ : std_logic;
signal \N__25739\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25731\ : std_logic;
signal \N__25728\ : std_logic;
signal \N__25725\ : std_logic;
signal \N__25722\ : std_logic;
signal \N__25719\ : std_logic;
signal \N__25716\ : std_logic;
signal \N__25711\ : std_logic;
signal \N__25706\ : std_logic;
signal \N__25703\ : std_logic;
signal \N__25700\ : std_logic;
signal \N__25697\ : std_logic;
signal \N__25694\ : std_logic;
signal \N__25691\ : std_logic;
signal \N__25688\ : std_logic;
signal \N__25685\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25681\ : std_logic;
signal \N__25680\ : std_logic;
signal \N__25677\ : std_logic;
signal \N__25676\ : std_logic;
signal \N__25671\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25665\ : std_logic;
signal \N__25662\ : std_logic;
signal \N__25657\ : std_logic;
signal \N__25652\ : std_logic;
signal \N__25649\ : std_logic;
signal \N__25646\ : std_logic;
signal \N__25643\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25641\ : std_logic;
signal \N__25634\ : std_logic;
signal \N__25631\ : std_logic;
signal \N__25630\ : std_logic;
signal \N__25627\ : std_logic;
signal \N__25624\ : std_logic;
signal \N__25621\ : std_logic;
signal \N__25618\ : std_logic;
signal \N__25613\ : std_logic;
signal \N__25612\ : std_logic;
signal \N__25609\ : std_logic;
signal \N__25606\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25602\ : std_logic;
signal \N__25597\ : std_logic;
signal \N__25594\ : std_logic;
signal \N__25591\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25587\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25573\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25562\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25556\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25535\ : std_logic;
signal \N__25532\ : std_logic;
signal \N__25529\ : std_logic;
signal \N__25526\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25520\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25508\ : std_logic;
signal \N__25505\ : std_logic;
signal \N__25504\ : std_logic;
signal \N__25503\ : std_logic;
signal \N__25498\ : std_logic;
signal \N__25495\ : std_logic;
signal \N__25492\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25488\ : std_logic;
signal \N__25483\ : std_logic;
signal \N__25480\ : std_logic;
signal \N__25477\ : std_logic;
signal \N__25474\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25466\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25459\ : std_logic;
signal \N__25456\ : std_logic;
signal \N__25453\ : std_logic;
signal \N__25450\ : std_logic;
signal \N__25447\ : std_logic;
signal \N__25442\ : std_logic;
signal \N__25439\ : std_logic;
signal \N__25436\ : std_logic;
signal \N__25433\ : std_logic;
signal \N__25430\ : std_logic;
signal \N__25427\ : std_logic;
signal \N__25424\ : std_logic;
signal \N__25421\ : std_logic;
signal \N__25418\ : std_logic;
signal \N__25415\ : std_logic;
signal \N__25412\ : std_logic;
signal \N__25409\ : std_logic;
signal \N__25406\ : std_logic;
signal \N__25403\ : std_logic;
signal \N__25400\ : std_logic;
signal \N__25397\ : std_logic;
signal \N__25394\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25388\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25376\ : std_logic;
signal \N__25373\ : std_logic;
signal \N__25370\ : std_logic;
signal \N__25367\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25358\ : std_logic;
signal \N__25355\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25349\ : std_logic;
signal \N__25346\ : std_logic;
signal \N__25343\ : std_logic;
signal \N__25340\ : std_logic;
signal \N__25337\ : std_logic;
signal \N__25334\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25319\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25304\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25297\ : std_logic;
signal \N__25294\ : std_logic;
signal \N__25291\ : std_logic;
signal \N__25288\ : std_logic;
signal \N__25285\ : std_logic;
signal \N__25282\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25274\ : std_logic;
signal \N__25271\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25265\ : std_logic;
signal \N__25264\ : std_logic;
signal \N__25263\ : std_logic;
signal \N__25260\ : std_logic;
signal \N__25257\ : std_logic;
signal \N__25254\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25244\ : std_logic;
signal \N__25241\ : std_logic;
signal \N__25238\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25226\ : std_logic;
signal \N__25223\ : std_logic;
signal \N__25220\ : std_logic;
signal \N__25217\ : std_logic;
signal \N__25214\ : std_logic;
signal \N__25211\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25193\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25184\ : std_logic;
signal \N__25181\ : std_logic;
signal \N__25178\ : std_logic;
signal \N__25175\ : std_logic;
signal \N__25172\ : std_logic;
signal \N__25169\ : std_logic;
signal \N__25166\ : std_logic;
signal \N__25163\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25157\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25151\ : std_logic;
signal \N__25148\ : std_logic;
signal \N__25145\ : std_logic;
signal \N__25142\ : std_logic;
signal \N__25139\ : std_logic;
signal \N__25136\ : std_logic;
signal \N__25133\ : std_logic;
signal \N__25130\ : std_logic;
signal \N__25127\ : std_logic;
signal \N__25124\ : std_logic;
signal \N__25121\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25115\ : std_logic;
signal \N__25112\ : std_logic;
signal \N__25109\ : std_logic;
signal \N__25106\ : std_logic;
signal \N__25103\ : std_logic;
signal \N__25100\ : std_logic;
signal \N__25097\ : std_logic;
signal \N__25094\ : std_logic;
signal \N__25091\ : std_logic;
signal \N__25088\ : std_logic;
signal \N__25085\ : std_logic;
signal \N__25082\ : std_logic;
signal \N__25079\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25070\ : std_logic;
signal \N__25067\ : std_logic;
signal \N__25064\ : std_logic;
signal \N__25061\ : std_logic;
signal \N__25058\ : std_logic;
signal \N__25055\ : std_logic;
signal \N__25052\ : std_logic;
signal \N__25049\ : std_logic;
signal \N__25046\ : std_logic;
signal \N__25043\ : std_logic;
signal \N__25040\ : std_logic;
signal \N__25037\ : std_logic;
signal \N__25034\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25028\ : std_logic;
signal \N__25027\ : std_logic;
signal \N__25024\ : std_logic;
signal \N__25021\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25015\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__25001\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24977\ : std_logic;
signal \N__24974\ : std_logic;
signal \N__24971\ : std_logic;
signal \N__24968\ : std_logic;
signal \N__24967\ : std_logic;
signal \N__24966\ : std_logic;
signal \N__24963\ : std_logic;
signal \N__24960\ : std_logic;
signal \N__24959\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24953\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24949\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24941\ : std_logic;
signal \N__24938\ : std_logic;
signal \N__24935\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24923\ : std_logic;
signal \N__24920\ : std_logic;
signal \N__24917\ : std_logic;
signal \N__24914\ : std_logic;
signal \N__24913\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24908\ : std_logic;
signal \N__24907\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24900\ : std_logic;
signal \N__24897\ : std_logic;
signal \N__24892\ : std_logic;
signal \N__24887\ : std_logic;
signal \N__24884\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24869\ : std_logic;
signal \N__24866\ : std_logic;
signal \N__24863\ : std_logic;
signal \N__24860\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24854\ : std_logic;
signal \N__24851\ : std_logic;
signal \N__24848\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24842\ : std_logic;
signal \N__24839\ : std_logic;
signal \N__24836\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24827\ : std_logic;
signal \N__24824\ : std_logic;
signal \N__24821\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24791\ : std_logic;
signal \N__24788\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24782\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24773\ : std_logic;
signal \N__24770\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24761\ : std_logic;
signal \N__24758\ : std_logic;
signal \N__24755\ : std_logic;
signal \N__24752\ : std_logic;
signal \N__24749\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24734\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24728\ : std_logic;
signal \N__24725\ : std_logic;
signal \N__24722\ : std_logic;
signal \N__24719\ : std_logic;
signal \N__24716\ : std_logic;
signal \N__24713\ : std_logic;
signal \N__24710\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24701\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24692\ : std_logic;
signal \N__24689\ : std_logic;
signal \N__24686\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24668\ : std_logic;
signal \N__24665\ : std_logic;
signal \N__24662\ : std_logic;
signal \N__24659\ : std_logic;
signal \N__24656\ : std_logic;
signal \N__24653\ : std_logic;
signal \N__24650\ : std_logic;
signal \N__24647\ : std_logic;
signal \N__24644\ : std_logic;
signal \N__24641\ : std_logic;
signal \N__24638\ : std_logic;
signal \N__24635\ : std_logic;
signal \N__24632\ : std_logic;
signal \N__24629\ : std_logic;
signal \N__24626\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24620\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24599\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24593\ : std_logic;
signal \N__24590\ : std_logic;
signal \N__24587\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24578\ : std_logic;
signal \N__24575\ : std_logic;
signal \N__24572\ : std_logic;
signal \N__24569\ : std_logic;
signal \N__24566\ : std_logic;
signal \N__24563\ : std_logic;
signal \N__24560\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24554\ : std_logic;
signal \N__24551\ : std_logic;
signal \N__24548\ : std_logic;
signal \N__24545\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24539\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24518\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24512\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24503\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24497\ : std_logic;
signal \N__24494\ : std_logic;
signal \N__24491\ : std_logic;
signal \N__24490\ : std_logic;
signal \N__24489\ : std_logic;
signal \N__24486\ : std_logic;
signal \N__24483\ : std_logic;
signal \N__24480\ : std_logic;
signal \N__24477\ : std_logic;
signal \N__24470\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24465\ : std_logic;
signal \N__24462\ : std_logic;
signal \N__24459\ : std_logic;
signal \N__24456\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24440\ : std_logic;
signal \N__24437\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24431\ : std_logic;
signal \N__24428\ : std_logic;
signal \N__24425\ : std_logic;
signal \N__24422\ : std_logic;
signal \N__24419\ : std_logic;
signal \N__24416\ : std_logic;
signal \N__24413\ : std_logic;
signal \N__24410\ : std_logic;
signal \N__24409\ : std_logic;
signal \N__24406\ : std_logic;
signal \N__24405\ : std_logic;
signal \N__24402\ : std_logic;
signal \N__24399\ : std_logic;
signal \N__24396\ : std_logic;
signal \N__24389\ : std_logic;
signal \N__24388\ : std_logic;
signal \N__24385\ : std_logic;
signal \N__24384\ : std_logic;
signal \N__24381\ : std_logic;
signal \N__24378\ : std_logic;
signal \N__24375\ : std_logic;
signal \N__24368\ : std_logic;
signal \N__24365\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24360\ : std_logic;
signal \N__24357\ : std_logic;
signal \N__24354\ : std_logic;
signal \N__24351\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24341\ : std_logic;
signal \N__24340\ : std_logic;
signal \N__24339\ : std_logic;
signal \N__24336\ : std_logic;
signal \N__24333\ : std_logic;
signal \N__24330\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24316\ : std_logic;
signal \N__24315\ : std_logic;
signal \N__24312\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24299\ : std_logic;
signal \N__24298\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24296\ : std_logic;
signal \N__24295\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24293\ : std_logic;
signal \N__24292\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24290\ : std_logic;
signal \N__24281\ : std_logic;
signal \N__24272\ : std_logic;
signal \N__24267\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24256\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24252\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24243\ : std_logic;
signal \N__24236\ : std_logic;
signal \N__24235\ : std_logic;
signal \N__24234\ : std_logic;
signal \N__24231\ : std_logic;
signal \N__24228\ : std_logic;
signal \N__24225\ : std_logic;
signal \N__24218\ : std_logic;
signal \N__24217\ : std_logic;
signal \N__24214\ : std_logic;
signal \N__24213\ : std_logic;
signal \N__24210\ : std_logic;
signal \N__24207\ : std_logic;
signal \N__24204\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24188\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24182\ : std_logic;
signal \N__24179\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24161\ : std_logic;
signal \N__24158\ : std_logic;
signal \N__24155\ : std_logic;
signal \N__24152\ : std_logic;
signal \N__24149\ : std_logic;
signal \N__24148\ : std_logic;
signal \N__24145\ : std_logic;
signal \N__24142\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24129\ : std_logic;
signal \N__24126\ : std_logic;
signal \N__24123\ : std_logic;
signal \N__24116\ : std_logic;
signal \N__24113\ : std_logic;
signal \N__24112\ : std_logic;
signal \N__24109\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24105\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24094\ : std_logic;
signal \N__24089\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24083\ : std_logic;
signal \N__24082\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24076\ : std_logic;
signal \N__24073\ : std_logic;
signal \N__24070\ : std_logic;
signal \N__24065\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24059\ : std_logic;
signal \N__24058\ : std_logic;
signal \N__24055\ : std_logic;
signal \N__24052\ : std_logic;
signal \N__24049\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24035\ : std_logic;
signal \N__24034\ : std_logic;
signal \N__24031\ : std_logic;
signal \N__24028\ : std_logic;
signal \N__24025\ : std_logic;
signal \N__24020\ : std_logic;
signal \N__24017\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24008\ : std_logic;
signal \N__24005\ : std_logic;
signal \N__24002\ : std_logic;
signal \N__24001\ : std_logic;
signal \N__24000\ : std_logic;
signal \N__23997\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23985\ : std_logic;
signal \N__23982\ : std_logic;
signal \N__23979\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23967\ : std_logic;
signal \N__23966\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23964\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23962\ : std_logic;
signal \N__23961\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23958\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23955\ : std_logic;
signal \N__23954\ : std_logic;
signal \N__23953\ : std_logic;
signal \N__23952\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23949\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23947\ : std_logic;
signal \N__23946\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23944\ : std_logic;
signal \N__23943\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23941\ : std_logic;
signal \N__23940\ : std_logic;
signal \N__23931\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23913\ : std_logic;
signal \N__23904\ : std_logic;
signal \N__23895\ : std_logic;
signal \N__23886\ : std_logic;
signal \N__23881\ : std_logic;
signal \N__23872\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23858\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23843\ : std_logic;
signal \N__23840\ : std_logic;
signal \N__23837\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23833\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23826\ : std_logic;
signal \N__23823\ : std_logic;
signal \N__23820\ : std_logic;
signal \N__23817\ : std_logic;
signal \N__23812\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23799\ : std_logic;
signal \N__23796\ : std_logic;
signal \N__23793\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23774\ : std_logic;
signal \N__23771\ : std_logic;
signal \N__23770\ : std_logic;
signal \N__23769\ : std_logic;
signal \N__23764\ : std_logic;
signal \N__23761\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23750\ : std_logic;
signal \N__23747\ : std_logic;
signal \N__23746\ : std_logic;
signal \N__23743\ : std_logic;
signal \N__23740\ : std_logic;
signal \N__23735\ : std_logic;
signal \N__23734\ : std_logic;
signal \N__23731\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23725\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23716\ : std_logic;
signal \N__23713\ : std_logic;
signal \N__23710\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23701\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23686\ : std_logic;
signal \N__23681\ : std_logic;
signal \N__23680\ : std_logic;
signal \N__23677\ : std_logic;
signal \N__23674\ : std_logic;
signal \N__23671\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23662\ : std_logic;
signal \N__23661\ : std_logic;
signal \N__23656\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23642\ : std_logic;
signal \N__23639\ : std_logic;
signal \N__23638\ : std_logic;
signal \N__23635\ : std_logic;
signal \N__23634\ : std_logic;
signal \N__23631\ : std_logic;
signal \N__23628\ : std_logic;
signal \N__23625\ : std_logic;
signal \N__23620\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23611\ : std_logic;
signal \N__23608\ : std_logic;
signal \N__23605\ : std_logic;
signal \N__23602\ : std_logic;
signal \N__23601\ : std_logic;
signal \N__23598\ : std_logic;
signal \N__23595\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23586\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23575\ : std_logic;
signal \N__23572\ : std_logic;
signal \N__23571\ : std_logic;
signal \N__23568\ : std_logic;
signal \N__23565\ : std_logic;
signal \N__23562\ : std_logic;
signal \N__23557\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23549\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23539\ : std_logic;
signal \N__23536\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23515\ : std_logic;
signal \N__23512\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23504\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23497\ : std_logic;
signal \N__23494\ : std_logic;
signal \N__23489\ : std_logic;
signal \N__23488\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23479\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23467\ : std_logic;
signal \N__23464\ : std_logic;
signal \N__23461\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23455\ : std_logic;
signal \N__23452\ : std_logic;
signal \N__23449\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23440\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23434\ : std_logic;
signal \N__23431\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23420\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23416\ : std_logic;
signal \N__23415\ : std_logic;
signal \N__23410\ : std_logic;
signal \N__23407\ : std_logic;
signal \N__23404\ : std_logic;
signal \N__23399\ : std_logic;
signal \N__23396\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23392\ : std_logic;
signal \N__23389\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23382\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23374\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23362\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23356\ : std_logic;
signal \N__23355\ : std_logic;
signal \N__23350\ : std_logic;
signal \N__23347\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23335\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23329\ : std_logic;
signal \N__23328\ : std_logic;
signal \N__23323\ : std_logic;
signal \N__23320\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23307\ : std_logic;
signal \N__23304\ : std_logic;
signal \N__23301\ : std_logic;
signal \N__23298\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23281\ : std_logic;
signal \N__23278\ : std_logic;
signal \N__23275\ : std_logic;
signal \N__23274\ : std_logic;
signal \N__23269\ : std_logic;
signal \N__23266\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23258\ : std_logic;
signal \N__23255\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23243\ : std_logic;
signal \N__23242\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23236\ : std_logic;
signal \N__23233\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23219\ : std_logic;
signal \N__23218\ : std_logic;
signal \N__23215\ : std_logic;
signal \N__23212\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23200\ : std_logic;
signal \N__23195\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23191\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23180\ : std_logic;
signal \N__23177\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23173\ : std_logic;
signal \N__23170\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23162\ : std_logic;
signal \N__23161\ : std_logic;
signal \N__23158\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23147\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23135\ : std_logic;
signal \N__23132\ : std_logic;
signal \N__23129\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23122\ : std_logic;
signal \N__23121\ : std_logic;
signal \N__23116\ : std_logic;
signal \N__23113\ : std_logic;
signal \N__23110\ : std_logic;
signal \N__23107\ : std_logic;
signal \N__23102\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23094\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23091\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23088\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23085\ : std_logic;
signal \N__23084\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23064\ : std_logic;
signal \N__23063\ : std_logic;
signal \N__23062\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23050\ : std_logic;
signal \N__23047\ : std_logic;
signal \N__23044\ : std_logic;
signal \N__23043\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23035\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23033\ : std_logic;
signal \N__23032\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23029\ : std_logic;
signal \N__23028\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23010\ : std_logic;
signal \N__23001\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22993\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22974\ : std_logic;
signal \N__22971\ : std_logic;
signal \N__22968\ : std_logic;
signal \N__22967\ : std_logic;
signal \N__22964\ : std_logic;
signal \N__22961\ : std_logic;
signal \N__22958\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22940\ : std_logic;
signal \N__22937\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22921\ : std_logic;
signal \N__22918\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22877\ : std_logic;
signal \N__22876\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22874\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22860\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22845\ : std_logic;
signal \N__22842\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22838\ : std_logic;
signal \N__22835\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22829\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22804\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22781\ : std_logic;
signal \N__22774\ : std_logic;
signal \N__22771\ : std_logic;
signal \N__22768\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22762\ : std_logic;
signal \N__22759\ : std_logic;
signal \N__22754\ : std_logic;
signal \N__22749\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22741\ : std_logic;
signal \N__22740\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22731\ : std_logic;
signal \N__22728\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22715\ : std_logic;
signal \N__22712\ : std_logic;
signal \N__22709\ : std_logic;
signal \N__22706\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22700\ : std_logic;
signal \N__22697\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22664\ : std_logic;
signal \N__22661\ : std_logic;
signal \N__22658\ : std_logic;
signal \N__22655\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22635\ : std_logic;
signal \N__22634\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22626\ : std_logic;
signal \N__22623\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22613\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22608\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22600\ : std_logic;
signal \N__22595\ : std_logic;
signal \N__22592\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22586\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22547\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22526\ : std_logic;
signal \N__22523\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22517\ : std_logic;
signal \N__22514\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22490\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22457\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22442\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22436\ : std_logic;
signal \N__22433\ : std_logic;
signal \N__22430\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22424\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22394\ : std_logic;
signal \N__22391\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22387\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22292\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22268\ : std_logic;
signal \N__22265\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22238\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22214\ : std_logic;
signal \N__22211\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22181\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22150\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22148\ : std_logic;
signal \N__22147\ : std_logic;
signal \N__22144\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22140\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22136\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22103\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22093\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22082\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22071\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21931\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21916\ : std_logic;
signal \N__21913\ : std_logic;
signal \N__21910\ : std_logic;
signal \N__21907\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21895\ : std_logic;
signal \N__21894\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21892\ : std_logic;
signal \N__21891\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21878\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21863\ : std_logic;
signal \N__21862\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21855\ : std_logic;
signal \N__21850\ : std_logic;
signal \N__21847\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21841\ : std_logic;
signal \N__21836\ : std_logic;
signal \N__21833\ : std_logic;
signal \N__21830\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21798\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21743\ : std_logic;
signal \N__21740\ : std_logic;
signal \N__21737\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21694\ : std_logic;
signal \N__21691\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21682\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21664\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21658\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21626\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21610\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21587\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21575\ : std_logic;
signal \N__21574\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21560\ : std_logic;
signal \N__21557\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21532\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21515\ : std_logic;
signal \N__21514\ : std_logic;
signal \N__21509\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21503\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21488\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21476\ : std_logic;
signal \N__21473\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21460\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21452\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21445\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21425\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21415\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21386\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21382\ : std_logic;
signal \N__21379\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21373\ : std_logic;
signal \N__21370\ : std_logic;
signal \N__21367\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21343\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21329\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21323\ : std_logic;
signal \N__21322\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21316\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21302\ : std_logic;
signal \N__21299\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21286\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21279\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21266\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21257\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21241\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21237\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21223\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21217\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21208\ : std_logic;
signal \N__21205\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21201\ : std_logic;
signal \N__21198\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21192\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21184\ : std_logic;
signal \N__21181\ : std_logic;
signal \N__21178\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21160\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21133\ : std_logic;
signal \N__21130\ : std_logic;
signal \N__21127\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21091\ : std_logic;
signal \N__21090\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21071\ : std_logic;
signal \N__21068\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21058\ : std_logic;
signal \N__21057\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21055\ : std_logic;
signal \N__21054\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21046\ : std_logic;
signal \N__21043\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21025\ : std_logic;
signal \N__21024\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21022\ : std_logic;
signal \N__21021\ : std_logic;
signal \N__21018\ : std_logic;
signal \N__21015\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__20998\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20954\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20945\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20918\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20896\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20890\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20884\ : std_logic;
signal \N__20881\ : std_logic;
signal \N__20878\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20870\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20863\ : std_logic;
signal \N__20860\ : std_logic;
signal \N__20859\ : std_logic;
signal \N__20854\ : std_logic;
signal \N__20851\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20845\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20819\ : std_logic;
signal \N__20816\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20800\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20791\ : std_logic;
signal \N__20788\ : std_logic;
signal \N__20785\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20779\ : std_logic;
signal \N__20776\ : std_logic;
signal \N__20773\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20747\ : std_logic;
signal \N__20744\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20737\ : std_logic;
signal \N__20734\ : std_logic;
signal \N__20729\ : std_logic;
signal \N__20726\ : std_logic;
signal \N__20723\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20710\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20703\ : std_logic;
signal \N__20700\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20673\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20667\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20657\ : std_logic;
signal \N__20654\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20648\ : std_logic;
signal \N__20645\ : std_logic;
signal \N__20642\ : std_logic;
signal \N__20639\ : std_logic;
signal \N__20636\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20630\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20626\ : std_logic;
signal \N__20623\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20613\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20610\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20604\ : std_logic;
signal \N__20603\ : std_logic;
signal \N__20602\ : std_logic;
signal \N__20601\ : std_logic;
signal \N__20600\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20598\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20559\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20557\ : std_logic;
signal \N__20556\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20553\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20540\ : std_logic;
signal \N__20537\ : std_logic;
signal \N__20532\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20530\ : std_logic;
signal \N__20529\ : std_logic;
signal \N__20526\ : std_logic;
signal \N__20523\ : std_logic;
signal \N__20520\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20503\ : std_logic;
signal \N__20500\ : std_logic;
signal \N__20493\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20474\ : std_logic;
signal \N__20471\ : std_logic;
signal \N__20466\ : std_logic;
signal \N__20463\ : std_logic;
signal \N__20450\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20448\ : std_logic;
signal \N__20447\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20445\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20431\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20421\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20402\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20400\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20398\ : std_logic;
signal \N__20397\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20383\ : std_logic;
signal \N__20380\ : std_logic;
signal \N__20379\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20362\ : std_logic;
signal \N__20361\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20311\ : std_logic;
signal \N__20308\ : std_logic;
signal \N__20305\ : std_logic;
signal \N__20302\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20293\ : std_logic;
signal \N__20290\ : std_logic;
signal \N__20285\ : std_logic;
signal \N__20284\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20278\ : std_logic;
signal \N__20275\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20260\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20243\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20231\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20201\ : std_logic;
signal \N__20198\ : std_logic;
signal \N__20195\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20163\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20154\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20140\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20126\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20117\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20108\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20094\ : std_logic;
signal \N__20091\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20082\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20054\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20048\ : std_logic;
signal \N__20045\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20041\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20036\ : std_logic;
signal \N__20035\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20032\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20007\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19996\ : std_logic;
signal \N__19995\ : std_logic;
signal \N__19990\ : std_logic;
signal \N__19987\ : std_logic;
signal \N__19984\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19943\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19890\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19887\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19882\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19872\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19864\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19858\ : std_logic;
signal \N__19855\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19839\ : std_logic;
signal \N__19836\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19828\ : std_logic;
signal \N__19827\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19815\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19813\ : std_logic;
signal \N__19810\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19791\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19780\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19688\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19679\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19675\ : std_logic;
signal \N__19674\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19666\ : std_logic;
signal \N__19665\ : std_logic;
signal \N__19662\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19657\ : std_logic;
signal \N__19654\ : std_logic;
signal \N__19651\ : std_logic;
signal \N__19638\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19583\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19576\ : std_logic;
signal \N__19575\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19567\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19555\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19551\ : std_logic;
signal \N__19548\ : std_logic;
signal \N__19545\ : std_logic;
signal \N__19542\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19525\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19518\ : std_logic;
signal \N__19515\ : std_logic;
signal \N__19512\ : std_logic;
signal \N__19509\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19436\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19406\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19400\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19391\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19304\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19280\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19262\ : std_logic;
signal \N__19259\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19244\ : std_logic;
signal \N__19241\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19223\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19196\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19169\ : std_logic;
signal \N__19166\ : std_logic;
signal \N__19163\ : std_logic;
signal \N__19160\ : std_logic;
signal \N__19157\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19145\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19136\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19130\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19103\ : std_logic;
signal \N__19100\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19091\ : std_logic;
signal \N__19088\ : std_logic;
signal \N__19085\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19079\ : std_logic;
signal \N__19076\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19052\ : std_logic;
signal \N__19049\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19043\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19034\ : std_logic;
signal \N__19031\ : std_logic;
signal \N__19028\ : std_logic;
signal \N__19025\ : std_logic;
signal \N__19022\ : std_logic;
signal \N__19019\ : std_logic;
signal \N__19016\ : std_logic;
signal \N__19015\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19007\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__18998\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18986\ : std_logic;
signal \N__18985\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18977\ : std_logic;
signal \N__18974\ : std_logic;
signal \N__18971\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18967\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18961\ : std_logic;
signal \N__18958\ : std_logic;
signal \N__18953\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18935\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18931\ : std_logic;
signal \N__18928\ : std_logic;
signal \N__18925\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18910\ : std_logic;
signal \N__18909\ : std_logic;
signal \N__18906\ : std_logic;
signal \N__18901\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18889\ : std_logic;
signal \N__18886\ : std_logic;
signal \N__18883\ : std_logic;
signal \N__18880\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18868\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18857\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18850\ : std_logic;
signal \N__18847\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18839\ : std_logic;
signal \N__18838\ : std_logic;
signal \N__18837\ : std_logic;
signal \N__18834\ : std_logic;
signal \N__18831\ : std_logic;
signal \N__18828\ : std_logic;
signal \N__18821\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18808\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18802\ : std_logic;
signal \N__18799\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18790\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18775\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18766\ : std_logic;
signal \N__18763\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18757\ : std_logic;
signal \N__18756\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18748\ : std_logic;
signal \N__18745\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18739\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18733\ : std_logic;
signal \N__18732\ : std_logic;
signal \N__18729\ : std_logic;
signal \N__18724\ : std_logic;
signal \N__18721\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18712\ : std_logic;
signal \N__18711\ : std_logic;
signal \N__18708\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18691\ : std_logic;
signal \N__18690\ : std_logic;
signal \N__18687\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18676\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18668\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18666\ : std_logic;
signal \N__18659\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18652\ : std_logic;
signal \N__18649\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18643\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18632\ : std_logic;
signal \N__18631\ : std_logic;
signal \N__18628\ : std_logic;
signal \N__18625\ : std_logic;
signal \N__18620\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18614\ : std_logic;
signal \N__18613\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18607\ : std_logic;
signal \N__18602\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18596\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18587\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18581\ : std_logic;
signal \N__18580\ : std_logic;
signal \N__18577\ : std_logic;
signal \N__18574\ : std_logic;
signal \N__18569\ : std_logic;
signal \N__18566\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18548\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18542\ : std_logic;
signal \N__18539\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18470\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18458\ : std_logic;
signal \N__18455\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18425\ : std_logic;
signal \N__18422\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18416\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18350\ : std_logic;
signal \N__18349\ : std_logic;
signal \N__18344\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18340\ : std_logic;
signal \N__18339\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18329\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18323\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18314\ : std_logic;
signal \N__18311\ : std_logic;
signal \N__18308\ : std_logic;
signal \N__18305\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18293\ : std_logic;
signal \N__18290\ : std_logic;
signal \N__18287\ : std_logic;
signal \N__18284\ : std_logic;
signal \N__18281\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18275\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_27_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_96_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_0_3_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_0_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_96\ : std_logic;
signal \pwm_generator_inst.O_0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_0\ : std_logic;
signal \bfn_1_7_0_\ : std_logic;
signal \pwm_generator_inst.O_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_0\ : std_logic;
signal \pwm_generator_inst.O_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_1\ : std_logic;
signal \pwm_generator_inst.O_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_2\ : std_logic;
signal \pwm_generator_inst.O_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_3\ : std_logic;
signal \pwm_generator_inst.O_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_4\ : std_logic;
signal \pwm_generator_inst.O_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_5\ : std_logic;
signal \pwm_generator_inst.O_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_7\ : std_logic;
signal \pwm_generator_inst.O_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_8\ : std_logic;
signal \bfn_1_8_0_\ : std_logic;
signal \pwm_generator_inst.O_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_15\ : std_logic;
signal \bfn_1_9_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_18\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc\ : std_logic;
signal \bfn_1_10_0_\ : std_logic;
signal \pwm_generator_inst.O_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_0\ : std_logic;
signal \pwm_generator_inst.O_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_1\ : std_logic;
signal \pwm_generator_inst.O_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_2\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_3\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_4\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_5\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_6\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_7\ : std_logic;
signal \bfn_1_11_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_9\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_10\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_15\ : std_logic;
signal \bfn_1_12_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_16\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_17\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_18\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_19\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_1_15\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_1_16\ : std_logic;
signal un7_start_stop_0_a3 : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\ : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_\ : std_logic;
signal pwm_duty_input_7 : std_logic;
signal pwm_duty_input_5 : std_logic;
signal pwm_duty_input_8 : std_logic;
signal pwm_duty_input_9 : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\ : std_logic;
signal pwm_duty_input_6 : std_logic;
signal \current_shift_inst.PI_CTRL.N_97\ : std_logic;
signal pwm_duty_input_0 : std_logic;
signal pwm_duty_input_2 : std_logic;
signal pwm_duty_input_1 : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_18\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO\ : std_logic;
signal \pwm_generator_inst.O_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_10_cascade_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_15_cascade_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_16\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_16_cascade_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_17\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4\ : std_logic;
signal \bfn_2_11_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_17\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_18\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_19\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_20\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_21\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_22\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_23\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0\ : std_logic;
signal \bfn_2_12_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_24\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_25\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16\ : std_logic;
signal \bfn_2_13_0_\ : std_logic;
signal \N_32_i_i\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_91\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_31\ : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\ : std_logic;
signal pwm_duty_input_3 : std_logic;
signal \pwm_generator_inst.un1_duty_inputlt3\ : std_logic;
signal pwm_duty_input_4 : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_0\ : std_logic;
signal \bfn_3_8_0_\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_0\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_1\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_7\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_7\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_8\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8\ : std_logic;
signal \bfn_3_9_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_8\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_178\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_118\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_9_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_2\ : std_logic;
signal \bfn_4_5_0_\ : std_logic;
signal un5_counter_cry_1 : std_logic;
signal un5_counter_cry_2 : std_logic;
signal un5_counter_cry_3 : std_logic;
signal un5_counter_cry_4 : std_logic;
signal un5_counter_cry_5 : std_logic;
signal un5_counter_cry_6 : std_logic;
signal un5_counter_cry_7 : std_logic;
signal un5_counter_cry_8 : std_logic;
signal \bfn_4_6_0_\ : std_logic;
signal un5_counter_cry_9 : std_logic;
signal un5_counter_cry_10 : std_logic;
signal un5_counter_cry_11 : std_logic;
signal \counterZ0Z_11\ : std_logic;
signal \counterZ0Z_9\ : std_logic;
signal \counterZ0Z_8\ : std_logic;
signal \counterZ0Z_2\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6\ : std_logic;
signal \counter_RNO_0Z0Z_7\ : std_logic;
signal \counterZ0Z_7\ : std_logic;
signal \N_19_1\ : std_logic;
signal \pwm_generator_inst.N_17\ : std_logic;
signal \pwm_generator_inst.N_16\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\ : std_logic;
signal clk_12mhz : std_logic;
signal \GB_BUFFER_clk_12mhz_THRU_CO\ : std_logic;
signal \counterZ0Z_4\ : std_logic;
signal \counterZ0Z_3\ : std_logic;
signal \counterZ0Z_5\ : std_logic;
signal \counterZ0Z_6\ : std_logic;
signal \un2_counter_5_cascade_\ : std_logic;
signal \counter_RNO_0Z0Z_12\ : std_logic;
signal \counterZ0Z_12\ : std_logic;
signal \counter_RNO_0Z0Z_10\ : std_logic;
signal \counterZ0Z_10\ : std_logic;
signal \counterZ0Z_1\ : std_logic;
signal \counterZ0Z_0\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_3\ : std_logic;
signal un2_counter_8 : std_logic;
signal un2_counter_7 : std_logic;
signal un2_counter_9 : std_logic;
signal \clk_10khz_RNIIENAZ0Z2_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_98\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\ : std_logic;
signal \bfn_5_9_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\ : std_logic;
signal \bfn_5_10_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\ : std_logic;
signal \bfn_5_11_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\ : std_logic;
signal \bfn_5_12_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un8_enablelto31\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_19\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_6\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_2\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_0\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_5\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_7\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_1\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_4\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_9\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_23\ : std_logic;
signal clk_10khz_i : std_logic;
signal \clk_10khz_RNIIENAZ0Z2\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lt19_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lt19_0_cascade_\ : std_logic;
signal \bfn_7_19_0_\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \bfn_7_20_0_\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \bfn_7_21_0_\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \bfn_7_22_0_\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \current_shift_inst.timer_phase.N_188_i_g\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_0\ : std_logic;
signal \pwm_generator_inst.counter_i_0\ : std_logic;
signal \bfn_8_8_0_\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_1\ : std_logic;
signal \pwm_generator_inst.counter_i_1\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_0\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counter_i_2\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_1\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_3\ : std_logic;
signal \pwm_generator_inst.counter_i_3\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_2\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_4\ : std_logic;
signal \pwm_generator_inst.counter_i_4\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_3\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_5\ : std_logic;
signal \pwm_generator_inst.counter_i_5\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_4\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_6\ : std_logic;
signal \pwm_generator_inst.counter_i_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_5\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_7\ : std_logic;
signal \pwm_generator_inst.counter_i_7\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_7\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_8\ : std_logic;
signal \pwm_generator_inst.counter_i_8\ : std_logic;
signal \bfn_8_9_0_\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_9\ : std_logic;
signal \pwm_generator_inst.counter_i_9\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_8\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_9\ : std_logic;
signal pwm_output_c : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_12_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_enablelt3_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto31_5_0\ : std_logic;
signal \bfn_8_13_0_\ : std_logic;
signal \current_shift_inst.control_input_1_cry_0\ : std_logic;
signal \current_shift_inst.control_input_1_cry_1\ : std_logic;
signal \current_shift_inst.control_input_1_cry_2\ : std_logic;
signal \current_shift_inst.control_input_1_cry_3\ : std_logic;
signal \current_shift_inst.control_input_1_cry_4\ : std_logic;
signal \current_shift_inst.control_input_1_cry_5\ : std_logic;
signal \current_shift_inst.control_input_1_cry_6\ : std_logic;
signal \current_shift_inst.control_input_1_cry_7\ : std_logic;
signal \bfn_8_14_0_\ : std_logic;
signal \current_shift_inst.control_input_1_cry_8\ : std_logic;
signal \current_shift_inst.control_input_1_cry_9\ : std_logic;
signal \current_shift_inst.control_input_1_cry_10\ : std_logic;
signal \current_shift_inst.control_input_1_cry_11\ : std_logic;
signal \current_shift_inst.control_input_1_cry_12\ : std_logic;
signal \current_shift_inst.control_input_1_cry_13\ : std_logic;
signal \current_shift_inst.control_input_1_cry_14\ : std_logic;
signal \current_shift_inst.control_input_1_cry_15\ : std_logic;
signal \bfn_8_15_0_\ : std_logic;
signal \current_shift_inst.control_input_1_cry_16\ : std_logic;
signal \current_shift_inst.control_input_1_cry_17\ : std_logic;
signal \current_shift_inst.control_input_1_cry_18\ : std_logic;
signal \current_shift_inst.control_input_1_cry_19\ : std_logic;
signal \current_shift_inst.control_input_1_cry_20\ : std_logic;
signal \current_shift_inst.control_input_1_cry_21\ : std_logic;
signal \current_shift_inst.control_input_1_cry_22\ : std_logic;
signal \current_shift_inst.control_input_1_cry_23\ : std_logic;
signal \bfn_8_16_0_\ : std_logic;
signal \current_shift_inst.control_input_1_cry_24\ : std_logic;
signal \bfn_8_17_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_2\ : std_logic;
signal \current_shift_inst.z_5_cry_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_3\ : std_logic;
signal \current_shift_inst.z_5_cry_2\ : std_logic;
signal \current_shift_inst.z_5_cry_3\ : std_logic;
signal \current_shift_inst.z_5_cry_4\ : std_logic;
signal \current_shift_inst.z_5_cry_5\ : std_logic;
signal \current_shift_inst.z_5_cry_6\ : std_logic;
signal \current_shift_inst.z_5_cry_7\ : std_logic;
signal \current_shift_inst.z_5_cry_8\ : std_logic;
signal \bfn_8_18_0_\ : std_logic;
signal \current_shift_inst.z_5_cry_9\ : std_logic;
signal \current_shift_inst.z_5_cry_10\ : std_logic;
signal \current_shift_inst.z_5_cry_11\ : std_logic;
signal \current_shift_inst.z_5_cry_12\ : std_logic;
signal \current_shift_inst.z_5_cry_13\ : std_logic;
signal \current_shift_inst.z_5_cry_14\ : std_logic;
signal \current_shift_inst.z_5_cry_15\ : std_logic;
signal \current_shift_inst.z_5_cry_16\ : std_logic;
signal \bfn_8_19_0_\ : std_logic;
signal \current_shift_inst.z_5_cry_17\ : std_logic;
signal \current_shift_inst.z_5_cry_18\ : std_logic;
signal \current_shift_inst.z_5_cry_19\ : std_logic;
signal \current_shift_inst.z_5_cry_20\ : std_logic;
signal \current_shift_inst.z_5_cry_21\ : std_logic;
signal \current_shift_inst.z_5_cry_22\ : std_logic;
signal \current_shift_inst.z_5_cry_23\ : std_logic;
signal \current_shift_inst.z_5_cry_24\ : std_logic;
signal \bfn_8_20_0_\ : std_logic;
signal \current_shift_inst.z_5_cry_25\ : std_logic;
signal \current_shift_inst.z_5_cry_26\ : std_logic;
signal \current_shift_inst.z_5_cry_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_29\ : std_logic;
signal \current_shift_inst.z_5_cry_28\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_30\ : std_logic;
signal \current_shift_inst.z_5_cry_29\ : std_logic;
signal \current_shift_inst.z_5_cry_30\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_0\ : std_logic;
signal \bfn_8_21_0_\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_1\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_0\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_2\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_1\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_3\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_2\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_4\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_3\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_5\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_4\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_6\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_5\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_7\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_6\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_7\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_8\ : std_logic;
signal \bfn_8_22_0_\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_9\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_8\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_10\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_9\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_11\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_10\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_12\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_11\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_13\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_12\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_14\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_13\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_15\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_14\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_15\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_16\ : std_logic;
signal \bfn_8_23_0_\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_17\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_16\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_18\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_17\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_19\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_18\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_20\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_19\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_21\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_20\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_22\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_21\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_23\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_22\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_23\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_24\ : std_logic;
signal \bfn_8_24_0_\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_25\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_24\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_26\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_25\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_27\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_26\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_28\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_27\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_28\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_29\ : std_logic;
signal \current_shift_inst.timer_s1.N_187_i\ : std_logic;
signal \current_shift_inst.timer_phase.N_193_i\ : std_logic;
signal \current_shift_inst.timer_phase.running_i\ : std_logic;
signal il_max_comp1_c : std_logic;
signal \bfn_9_7_0_\ : std_logic;
signal \pwm_generator_inst.counter_cry_0\ : std_logic;
signal \pwm_generator_inst.counter_cry_1\ : std_logic;
signal \pwm_generator_inst.counter_cry_2\ : std_logic;
signal \pwm_generator_inst.counter_cry_3\ : std_logic;
signal \pwm_generator_inst.counter_cry_4\ : std_logic;
signal \pwm_generator_inst.counter_cry_5\ : std_logic;
signal \pwm_generator_inst.counter_cry_6\ : std_logic;
signal \pwm_generator_inst.counter_cry_7\ : std_logic;
signal \bfn_9_8_0_\ : std_logic;
signal \pwm_generator_inst.counter_cry_8\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_3\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_1\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_4\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_6\ : std_logic;
signal \pwm_generator_inst.un1_counterlt9_cascade_\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_5\ : std_logic;
signal \pwm_generator_inst.un1_counter_0\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_9\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_8\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_7\ : std_logic;
signal \pwm_generator_inst.un1_counterlto9_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_0\ : std_logic;
signal \pwm_generator_inst.un1_counterlto2_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_11_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_44\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_43\ : std_logic;
signal \bfn_9_13_0_\ : std_logic;
signal \current_shift_inst.z_i_0_31\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CO\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_2_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_1\ : std_logic;
signal \current_shift_inst.N_1620_i\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_3_c_invZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_2\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_3\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_4\ : std_logic;
signal \current_shift_inst.control_input_1_axb_0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_5\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_6\ : std_logic;
signal \current_shift_inst.control_input_1_axb_1\ : std_logic;
signal \bfn_9_14_0_\ : std_logic;
signal \current_shift_inst.control_input_1_axb_2\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_7\ : std_logic;
signal \current_shift_inst.control_input_1_axb_3\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_8\ : std_logic;
signal \current_shift_inst.control_input_1_axb_4\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_9\ : std_logic;
signal \current_shift_inst.control_input_1_axb_5\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_10\ : std_logic;
signal \current_shift_inst.control_input_1_axb_6\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJTQ51_12\ : std_logic;
signal \current_shift_inst.control_input_1_axb_7\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIR0UI_13\ : std_logic;
signal \current_shift_inst.control_input_1_axb_8\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_13\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_14\ : std_logic;
signal \current_shift_inst.control_input_1_axb_9\ : std_logic;
signal \bfn_9_15_0_\ : std_logic;
signal \current_shift_inst.control_input_1_axb_10\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_15\ : std_logic;
signal \current_shift_inst.control_input_1_axb_11\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_16\ : std_logic;
signal \current_shift_inst.control_input_1_axb_12\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_17\ : std_logic;
signal \current_shift_inst.control_input_1_axb_13\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_18\ : std_logic;
signal \current_shift_inst.control_input_1_axb_14\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_19\ : std_logic;
signal \current_shift_inst.control_input_1_axb_15\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_20\ : std_logic;
signal \current_shift_inst.control_input_1_axb_16\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_21\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_22\ : std_logic;
signal \current_shift_inst.control_input_1_axb_17\ : std_logic;
signal \bfn_9_16_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIU73K_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIVJ781_23\ : std_logic;
signal \current_shift_inst.control_input_1_axb_18\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_23\ : std_logic;
signal \current_shift_inst.control_input_1_axb_19\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIB4C81_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI4G5K_25\ : std_logic;
signal \current_shift_inst.control_input_1_axb_20\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_25\ : std_logic;
signal \current_shift_inst.control_input_1_axb_21\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIAO7K_27\ : std_logic;
signal \current_shift_inst.control_input_1_axb_22\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIDS8K_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIKKJ81_29\ : std_logic;
signal \current_shift_inst.control_input_1_axb_23\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIVQF91_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI7OAK_29\ : std_logic;
signal \current_shift_inst.control_input_1_axb_24\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_29\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_30\ : std_logic;
signal \current_shift_inst.un38_control_input_0_axb_31\ : std_logic;
signal \current_shift_inst.control_input_1_cry_24_THRU_CO\ : std_logic;
signal \bfn_9_17_0_\ : std_logic;
signal \current_shift_inst.phase_valid_RNISLORZ0Z2\ : std_logic;
signal \G_406\ : std_logic;
signal \bfn_9_18_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_1\ : std_logic;
signal \G_405\ : std_logic;
signal \current_shift_inst.z_cry_0\ : std_logic;
signal \current_shift_inst.z_5_2\ : std_logic;
signal \current_shift_inst.z_cry_1\ : std_logic;
signal \current_shift_inst.z_5_3\ : std_logic;
signal \current_shift_inst.z_cry_2\ : std_logic;
signal \current_shift_inst.z_5_4\ : std_logic;
signal \current_shift_inst.z_cry_3\ : std_logic;
signal \current_shift_inst.z_5_5\ : std_logic;
signal \current_shift_inst.z_cry_4\ : std_logic;
signal \current_shift_inst.z_5_6\ : std_logic;
signal \current_shift_inst.z_cry_5\ : std_logic;
signal \current_shift_inst.z_5_7\ : std_logic;
signal \current_shift_inst.z_cry_6\ : std_logic;
signal \current_shift_inst.z_cry_7\ : std_logic;
signal \current_shift_inst.z_5_8\ : std_logic;
signal \bfn_9_19_0_\ : std_logic;
signal \current_shift_inst.z_5_9\ : std_logic;
signal \current_shift_inst.z_cry_8\ : std_logic;
signal \current_shift_inst.z_5_10\ : std_logic;
signal \current_shift_inst.z_cry_9\ : std_logic;
signal \current_shift_inst.z_5_11\ : std_logic;
signal \current_shift_inst.z_cry_10\ : std_logic;
signal \current_shift_inst.z_5_12\ : std_logic;
signal \current_shift_inst.z_cry_11\ : std_logic;
signal \current_shift_inst.z_5_13\ : std_logic;
signal \current_shift_inst.z_cry_12\ : std_logic;
signal \current_shift_inst.z_5_14\ : std_logic;
signal \current_shift_inst.z_cry_13\ : std_logic;
signal \current_shift_inst.z_5_15\ : std_logic;
signal \current_shift_inst.z_cry_14\ : std_logic;
signal \current_shift_inst.z_cry_15\ : std_logic;
signal \current_shift_inst.z_5_16\ : std_logic;
signal \bfn_9_20_0_\ : std_logic;
signal \current_shift_inst.z_5_17\ : std_logic;
signal \current_shift_inst.z_cry_16\ : std_logic;
signal \current_shift_inst.z_5_18\ : std_logic;
signal \current_shift_inst.z_cry_17\ : std_logic;
signal \current_shift_inst.z_5_19\ : std_logic;
signal \current_shift_inst.z_cry_18\ : std_logic;
signal \current_shift_inst.z_5_20\ : std_logic;
signal \current_shift_inst.z_cry_19\ : std_logic;
signal \current_shift_inst.z_5_21\ : std_logic;
signal \current_shift_inst.z_cry_20\ : std_logic;
signal \current_shift_inst.z_5_22\ : std_logic;
signal \current_shift_inst.z_cry_21\ : std_logic;
signal \current_shift_inst.z_5_23\ : std_logic;
signal \current_shift_inst.z_cry_22\ : std_logic;
signal \current_shift_inst.z_cry_23\ : std_logic;
signal \current_shift_inst.z_5_24\ : std_logic;
signal \bfn_9_21_0_\ : std_logic;
signal \current_shift_inst.z_5_25\ : std_logic;
signal \current_shift_inst.z_cry_24\ : std_logic;
signal \current_shift_inst.z_5_26\ : std_logic;
signal \current_shift_inst.z_cry_25\ : std_logic;
signal \current_shift_inst.z_5_27\ : std_logic;
signal \current_shift_inst.z_cry_26\ : std_logic;
signal \current_shift_inst.z_5_28\ : std_logic;
signal \current_shift_inst.z_cry_27\ : std_logic;
signal \current_shift_inst.z_5_29\ : std_logic;
signal \current_shift_inst.z_cry_28\ : std_logic;
signal \current_shift_inst.z_5_30\ : std_logic;
signal \current_shift_inst.z_cry_29\ : std_logic;
signal \current_shift_inst.z_5_cry_30_THRU_CO\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_31\ : std_logic;
signal \current_shift_inst.z_cry_30\ : std_logic;
signal \current_shift_inst.stop_timer_s1_RNOZ0Z_0\ : std_logic;
signal \current_shift_inst.start_timer_phaseZ0\ : std_logic;
signal \il_max_comp1_D1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_4_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0Z_0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIVQKU1_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNILORI_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIN7DV_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIOSSI_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI1PG21_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIER9V_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIP5T51_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_4\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5M161_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIIKQI_10\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI4D1J_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIVDV51_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIK3CV_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI53NU1_6\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_6\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIHVAV_6\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI7DM51_10\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI4H5J_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_10\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJDBL1_10\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIBBPU1_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIU4VI_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIO0U12_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIE6961_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJ3381_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIOV0K_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIAL3J_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI7H2J_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNILRVJ_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPC571_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIBU361_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI190J_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIDR081_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIH6661_17\ : std_logic;
signal \current_shift_inst.un38_control_input_0\ : std_logic;
signal \bfn_10_17_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_1\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_2\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_3_c_RNINL4GZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_3\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_4\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_5\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_6\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_7\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_8\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0\ : std_logic;
signal \bfn_10_18_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_9_c_RNIALDJZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_9\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_10_c_RNIJLTGZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_10\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_11\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_12\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_13\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_14\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_15\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_16\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0\ : std_logic;
signal \bfn_10_19_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_17\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_18\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_19\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_20\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_21\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_22\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_23\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_24\ : std_logic;
signal \bfn_10_20_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_25\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_26\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_27\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_28\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_30\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_28\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNINKG81_27\ : std_logic;
signal \bfn_10_21_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_0\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_1\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_7\ : std_logic;
signal \bfn_10_22_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_9\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_15\ : std_logic;
signal \bfn_10_23_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_17\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_23\ : std_logic;
signal \bfn_10_24_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_25\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.running_i\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_28\ : std_logic;
signal \current_shift_inst.start_timer_sZ0Z1\ : std_logic;
signal \current_shift_inst.timer_s1.runningZ0\ : std_logic;
signal \current_shift_inst.stop_timer_sZ0Z1\ : std_logic;
signal \current_shift_inst.timer_s1.N_192_i\ : std_logic;
signal \current_shift_inst.timer_phase.runningZ0\ : std_logic;
signal \current_shift_inst.stop_timer_phaseZ0\ : std_logic;
signal \current_shift_inst.timer_phase.N_188_i\ : std_logic;
signal il_max_comp2_c : std_logic;
signal il_min_comp2_c : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_0\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_axb_0\ : std_logic;
signal \bfn_11_10_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_1\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_0\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_1\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_4\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_5\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_6\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_7\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_8\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\ : std_logic;
signal \bfn_11_11_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_9\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_10\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_11\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_12\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_13\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_14\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_15\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_16\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\ : std_logic;
signal \bfn_11_12_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_17\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_18\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_19\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_18\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_21\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_22\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_23\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_23\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_24\ : std_logic;
signal \bfn_11_13_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_29\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto31_cZ0Z_0_cascade_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_fast_31\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_1\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_1\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_2\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_2\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_14\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_3\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_4\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_5\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_6\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_7\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_8\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_13\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_15\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_9\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_10\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_11\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_12\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_16\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_20\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_18\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_23\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_19\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_25\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_22\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_24\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_17\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_21\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_26\ : std_logic;
signal \current_shift_inst.z_31\ : std_logic;
signal \current_shift_inst.z_i_31\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_30\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_27\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_29\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_28\ : std_logic;
signal \current_shift_inst.S1_sync_prevZ0\ : std_logic;
signal \current_shift_inst.S1_syncZ0Z0\ : std_logic;
signal \current_shift_inst.S1_syncZ0Z1\ : std_logic;
signal \current_shift_inst.meas_stateZ0Z_0\ : std_logic;
signal \current_shift_inst.S1_riseZ0\ : std_logic;
signal \current_shift_inst.phase_validZ0\ : std_logic;
signal il_min_comp1_c : std_logic;
signal \il_min_comp1_D1\ : std_logic;
signal \il_min_comp2_D1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_m5_iZ0Z_1_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_N_4_cascade_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_11\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIDLO51_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI1C4K_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_27\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIHCE81_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_23\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPB581_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_22\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIR32K_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_26\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI7K6K_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_24\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5S981_24\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_0\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_3\ : std_logic;
signal \bfn_12_19_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_1\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_4\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_2\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_5\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_3\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_6\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_4\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_7\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_5\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_6\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_9\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_7\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_10\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_8\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_11\ : std_logic;
signal \bfn_12_20_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_9\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_12\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_10\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_13\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_11\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_14\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_12\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_15\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_13\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_16\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_14\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_17\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_15\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_18\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_16\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_19\ : std_logic;
signal \bfn_12_21_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_17\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_20\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_18\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_21\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_19\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_22\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_20\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_23\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_21\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_24\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_22\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_25\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_23\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_26\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_24\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_27\ : std_logic;
signal \bfn_12_22_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_25\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_28\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_28\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_26\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_29\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_29\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_27\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_30\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.N_187_i_g\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\ : std_logic;
signal s1_phy_c : std_logic;
signal \current_shift_inst.S3_riseZ0\ : std_logic;
signal \current_shift_inst.S3_sync_prevZ0\ : std_logic;
signal \current_shift_inst.S3_syncZ0Z0\ : std_logic;
signal \current_shift_inst.S3_syncZ0Z1\ : std_logic;
signal \il_max_comp2_D1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_47\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_79\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_27\ : std_logic;
signal \N_605_g\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto13_3Z0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto30_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto8Z0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_m2_eZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_11_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlt31_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_0\ : std_logic;
signal \bfn_13_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ1Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \bfn_13_14_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_16\ : std_logic;
signal \bfn_13_15_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\ : std_logic;
signal \phase_controller_slave.stoper_tr.time_passed_1_sqmuxa\ : std_logic;
signal \phase_controller_slave.tr_time_passed\ : std_logic;
signal \phase_controller_slave.stateZ0Z_0\ : std_logic;
signal \phase_controller_slave.state_RNIVDE2Z0Z_0_cascade_\ : std_logic;
signal state_ns_i_a2_1 : std_logic;
signal start_stop_c : std_logic;
signal s4_phy_c : std_logic;
signal \il_min_comp2_D2\ : std_logic;
signal \phase_controller_slave.stateZ0Z_1\ : std_logic;
signal \phase_controller_slave.start_timer_tr_0_sqmuxa\ : std_logic;
signal \phase_controller_slave.state_RNIVDE2Z0Z_0\ : std_logic;
signal s3_phy_c : std_logic;
signal shift_flag_start : std_logic;
signal \phase_controller_inst1.state_RNI7NN7Z0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa\ : std_logic;
signal \phase_controller_inst1.start_timer_tr_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.tr_time_passed\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_0\ : std_logic;
signal \bfn_13_24_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7\ : std_logic;
signal \bfn_13_25_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15\ : std_logic;
signal \bfn_13_26_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0\ : std_logic;
signal s2_phy_c : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_335_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_2_cascade_\ : std_logic;
signal \il_min_comp1_D2\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.time_passed11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_m2_eZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_m2_eZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8\ : std_logic;
signal measured_delay_hc_23 : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_3\ : std_logic;
signal \phase_controller_inst1.start_timer_hc_0_sqmuxa_cascade_\ : std_logic;
signal \phase_controller_inst1.start_timer_hc_RNOZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_3\ : std_logic;
signal \il_max_comp1_D2\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa\ : std_logic;
signal \phase_controller_inst1.hc_time_passed\ : std_logic;
signal \phase_controller_inst1.stoper_hc.time_passed11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.time_passed11_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_N_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto31_dZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_start_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto31_dZ0Z_0_cascade_\ : std_logic;
signal measured_delay_hc_16 : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto31_cZ0Z_0\ : std_logic;
signal measured_delay_hc_17 : std_logic;
signal measured_delay_hc_10 : std_logic;
signal measured_delay_hc_11 : std_logic;
signal measured_delay_hc_2 : std_logic;
signal measured_delay_hc_7 : std_logic;
signal measured_delay_hc_5 : std_logic;
signal measured_delay_hc_12 : std_logic;
signal measured_delay_hc_1 : std_logic;
signal measured_delay_hc_3 : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_2\ : std_logic;
signal measured_delay_hc_15 : std_logic;
signal measured_delay_hc_13 : std_logic;
signal measured_delay_hc_18 : std_logic;
signal measured_delay_hc_6 : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlt31_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlt31\ : std_logic;
signal measured_delay_hc_8 : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_start\ : std_logic;
signal \bfn_14_18_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7\ : std_logic;
signal \bfn_14_19_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15\ : std_logic;
signal \bfn_14_20_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\ : std_logic;
signal delay_tr_input_c : std_logic;
signal delay_tr_d1 : std_logic;
signal red_c_i : std_logic;
signal \delay_measurement_inst.prev_hc_sigZ0\ : std_logic;
signal \delay_measurement_inst.hc_stateZ0Z_0\ : std_logic;
signal delay_tr_d2 : std_logic;
signal \delay_measurement_inst.tr_stateZ0Z_0\ : std_logic;
signal \delay_measurement_inst.prev_tr_sigZ0\ : std_logic;
signal delay_hc_input_c : std_logic;
signal delay_hc_d1 : std_logic;
signal delay_hc_d2 : std_logic;
signal measured_delay_hc_9 : std_logic;
signal \delay_measurement_inst.start_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6_cascade_\ : std_logic;
signal \delay_measurement_inst.stop_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt15_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto6_c_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto6_0_0_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt9\ : std_logic;
signal measured_delay_hc_21 : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1\ : std_logic;
signal measured_delay_hc_20 : std_logic;
signal measured_delay_hc_19 : std_logic;
signal measured_delay_hc_22 : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto31_0_0\ : std_logic;
signal measured_delay_hc_29 : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_4\ : std_logic;
signal measured_delay_hc_27 : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_15_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9\ : std_logic;
signal \bfn_15_14_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17\ : std_logic;
signal \bfn_15_15_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_0\ : std_logic;
signal \bfn_15_16_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ1Z_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \bfn_15_17_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_16\ : std_logic;
signal \bfn_15_18_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_18\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_19\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.time_passed11\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_slave.start_timer_trZ0\ : std_logic;
signal \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_15_21_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_15_22_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_17\ : std_logic;
signal \bfn_15_23_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_19\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_15_24_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_15_25_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_17\ : std_logic;
signal \bfn_15_26_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \delay_measurement_inst.start_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.stop_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.runningZ0\ : std_logic;
signal \bfn_16_7_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_7\ : std_logic;
signal \bfn_16_8_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_15\ : std_logic;
signal \bfn_16_9_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_23\ : std_logic;
signal \bfn_16_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_336_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_a1_2_0_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_a1_2_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto30_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto30_2_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3_cascade_\ : std_logic;
signal measured_delay_hc_4 : std_logic;
signal measured_delay_hc_14 : std_logic;
signal measured_delay_hc_24 : std_logic;
signal measured_delay_hc_25 : std_logic;
signal measured_delay_hc_26 : std_logic;
signal measured_delay_hc_28 : std_logic;
signal measured_delay_hc_30 : std_logic;
signal measured_delay_hc_0 : std_logic;
signal \delay_measurement_inst.delay_hc_reg3\ : std_logic;
signal \delay_measurement_inst.un1_elapsed_time_hc\ : std_logic;
signal measured_delay_hc_31 : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6_cascade_\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal measured_delay_tr_10 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal measured_delay_tr_9 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal measured_delay_tr_12 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\ : std_logic;
signal \bfn_17_8_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_11\ : std_logic;
signal \bfn_17_9_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\ : std_logic;
signal \bfn_17_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\ : std_logic;
signal \bfn_17_11_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_4\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto5_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIB3GH4Z0Z_3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_7_0\ : std_logic;
signal \bfn_17_13_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_7\ : std_logic;
signal \bfn_17_14_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_15\ : std_logic;
signal \bfn_17_15_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_23\ : std_logic;
signal \bfn_17_16_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_338_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_293\ : std_logic;
signal \delay_measurement_inst.N_358_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19\ : std_logic;
signal \delay_measurement_inst.N_307\ : std_logic;
signal \phase_controller_slave.start_timer_hc_RNO_0_0\ : std_logic;
signal \phase_controller_slave.start_timer_hc_0_sqmuxa_cascade_\ : std_logic;
signal phase_controller_inst1_state_4 : std_logic;
signal \il_max_comp2_D2\ : std_logic;
signal \phase_controller_slave.stateZ0Z_3\ : std_logic;
signal \phase_controller_slave.stateZ0Z_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.time_passed11\ : std_logic;
signal \phase_controller_slave.stoper_hc.time_passed_1_sqmuxa\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_slave.hc_time_passed\ : std_logic;
signal \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_slave.start_timer_hcZ0\ : std_logic;
signal \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4Z0Z_3_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_279\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_262\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_335_i_g\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_18\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_17\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_19\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_16\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_a0_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto9\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_a0_1_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto19_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_a0_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\ : std_logic;
signal \bfn_18_15_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\ : std_logic;
signal \bfn_18_16_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\ : std_logic;
signal \bfn_18_17_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\ : std_logic;
signal \bfn_18_18_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_337_i\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_18_19_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9\ : std_logic;
signal \bfn_18_20_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17\ : std_logic;
signal \bfn_18_21_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_reg3lto9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_320_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_320_4_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_12\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_10\ : std_logic;
signal \delay_measurement_inst.N_328\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_331_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_321_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILUISZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_331\ : std_logic;
signal \delay_measurement_inst.delay_tr_reg_esr_RNO_0Z0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_reg3lto14\ : std_logic;
signal measured_delay_tr_14 : std_logic;
signal \delay_measurement_inst.delay_tr_reg3lto15\ : std_logic;
signal \delay_measurement_inst.elapsed_time_ns_1_RNIM96P1_16\ : std_logic;
signal measured_delay_tr_15 : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_1\ : std_logic;
signal measured_delay_tr_1 : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_5\ : std_logic;
signal measured_delay_tr_5 : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_3\ : std_logic;
signal measured_delay_tr_3 : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_8\ : std_logic;
signal measured_delay_tr_8 : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_7\ : std_logic;
signal measured_delay_tr_7 : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_17\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_13\ : std_logic;
signal measured_delay_tr_13 : std_logic;
signal \delay_measurement_inst.delay_tr_reg3lto6\ : std_logic;
signal measured_delay_tr_6 : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_4\ : std_logic;
signal measured_delay_tr_4 : std_logic;
signal \delay_measurement_inst.N_324\ : std_logic;
signal \delay_measurement_inst.elapsed_time_ns_1_RNI80KG7_6\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_2\ : std_logic;
signal measured_delay_tr_2 : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_16\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_11\ : std_logic;
signal \delay_measurement_inst.N_301\ : std_logic;
signal measured_delay_tr_11 : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_18\ : std_logic;
signal measured_delay_tr_18 : std_logic;
signal measured_delay_tr_17 : std_logic;
signal measured_delay_tr_16 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3Z0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_i\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_31\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_19\ : std_logic;
signal \delay_measurement_inst.N_358\ : std_logic;
signal measured_delay_tr_19 : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_100mhz_0 : std_logic;
signal \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\ : std_logic;
signal red_c_g : std_logic;

signal reset_wire : std_logic;
signal start_stop_wire : std_logic;
signal il_max_comp2_wire : std_logic;
signal pwm_output_wire : std_logic;
signal il_max_comp1_wire : std_logic;
signal s2_phy_wire : std_logic;
signal delay_hc_input_wire : std_logic;
signal delay_tr_input_wire : std_logic;
signal il_min_comp2_wire : std_logic;
signal s1_phy_wire : std_logic;
signal s4_phy_wire : std_logic;
signal il_min_comp1_wire : std_logic;
signal s3_phy_wire : std_logic;
signal rgb_b_wire : std_logic;
signal rgb_g_wire : std_logic;
signal rgb_r_wire : std_logic;
signal \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);

begin
    reset_wire <= reset;
    start_stop_wire <= start_stop;
    il_max_comp2_wire <= il_max_comp2;
    pwm_output <= pwm_output_wire;
    il_max_comp1_wire <= il_max_comp1;
    s2_phy <= s2_phy_wire;
    delay_hc_input_wire <= delay_hc_input;
    delay_tr_input_wire <= delay_tr_input;
    il_min_comp2_wire <= il_min_comp2;
    s1_phy <= s1_phy_wire;
    s4_phy <= s4_phy_wire;
    il_min_comp1_wire <= il_min_comp1;
    s3_phy <= s3_phy_wire;
    rgb_b <= rgb_b_wire;
    rgb_g <= rgb_g_wire;
    rgb_r <= rgb_r_wire;
    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_A_wire\ <= '0'&\N__20529\&\N__20557\&\N__20530\&\N__20558\&\N__20531\&\N__18716\&\N__18740\&\N__18779\&\N__18692\&\N__18758\&\N__19525\&\N__19551\&\N__18643\&\N__18631\&\N__18655\;
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__23095\&\N__23092\&'0'&'0'&'0'&\N__23090\&\N__23094\&\N__23091\&\N__23093\;
    \pwm_generator_inst.un2_threshold_acc_1_25\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(25);
    \pwm_generator_inst.un2_threshold_acc_1_24\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(24);
    \pwm_generator_inst.un2_threshold_acc_1_23\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(23);
    \pwm_generator_inst.un2_threshold_acc_1_22\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(22);
    \pwm_generator_inst.un2_threshold_acc_1_21\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(21);
    \pwm_generator_inst.un2_threshold_acc_1_20\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(20);
    \pwm_generator_inst.un2_threshold_acc_1_19\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(19);
    \pwm_generator_inst.un2_threshold_acc_1_18\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(18);
    \pwm_generator_inst.un2_threshold_acc_1_17\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(17);
    \pwm_generator_inst.un2_threshold_acc_1_16\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_acc_1_15\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.O_14\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.O_13\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.O_12\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un3_threshold_acc\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.O_10\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.O_9\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.O_8\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.O_7\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.O_6\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.O_5\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.O_4\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.O_3\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.O_2\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.O_1\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.O_0\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_A_wire\ <= '0'&\N__20612\&\N__20605\&\N__20610\&\N__20604\&\N__20611\&\N__20603\&\N__20613\&\N__20600\&\N__20606\&\N__20599\&\N__20607\&\N__20601\&\N__20608\&\N__20602\&\N__20609\;
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__23063\&\N__23060\&'0'&'0'&'0'&\N__23058\&\N__23062\&\N__23059\&\N__23061\;
    \pwm_generator_inst.un2_threshold_acc_2_1_16\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_acc_2_1_15\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.un2_threshold_acc_2_14\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.un2_threshold_acc_2_13\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.un2_threshold_acc_2_12\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un2_threshold_acc_2_11\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.un2_threshold_acc_2_10\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.un2_threshold_acc_2_9\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.un2_threshold_acc_2_8\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.un2_threshold_acc_2_7\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.un2_threshold_acc_2_6\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.un2_threshold_acc_2_5\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.un2_threshold_acc_2_4\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.un2_threshold_acc_2_3\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.un2_threshold_acc_2_2\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.un2_threshold_acc_2_1\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.un2_threshold_acc_2_0\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(0);

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__20819\,
            RESETB => \N__35880\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => clk_100mhz_0
        );

    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__23099\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__23089\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__23064\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__23057\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\
        );

    \reset_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__48678\,
            GLOBALBUFFEROUTPUT => red_c_g
        );

    \reset_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48680\,
            DIN => \N__48679\,
            DOUT => \N__48678\,
            PACKAGEPIN => reset_wire
        );

    \reset_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48680\,
            PADOUT => \N__48679\,
            PADIN => \N__48678\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \start_stop_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48669\,
            DIN => \N__48668\,
            DOUT => \N__48667\,
            PACKAGEPIN => start_stop_wire
        );

    \start_stop_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48669\,
            PADOUT => \N__48668\,
            PADIN => \N__48667\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => start_stop_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48660\,
            DIN => \N__48659\,
            DOUT => \N__48658\,
            PACKAGEPIN => il_max_comp2_wire
        );

    \il_max_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48660\,
            PADOUT => \N__48659\,
            PADIN => \N__48658\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48651\,
            DIN => \N__48650\,
            DOUT => \N__48649\,
            PACKAGEPIN => pwm_output_wire
        );

    \pwm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48651\,
            PADOUT => \N__48650\,
            PADIN => \N__48649\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__22418\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48642\,
            DIN => \N__48641\,
            DOUT => \N__48640\,
            PACKAGEPIN => il_max_comp1_wire
        );

    \il_max_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48642\,
            PADOUT => \N__48641\,
            PADIN => \N__48640\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s2_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48633\,
            DIN => \N__48632\,
            DOUT => \N__48631\,
            PACKAGEPIN => s2_phy_wire
        );

    \s2_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48633\,
            PADOUT => \N__48632\,
            PADIN => \N__48631\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__34073\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_hc_input_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48624\,
            DIN => \N__48623\,
            DOUT => \N__48622\,
            PACKAGEPIN => delay_hc_input_wire
        );

    \delay_hc_input_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48624\,
            PADOUT => \N__48623\,
            PADIN => \N__48622\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_hc_input_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_tr_input_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48615\,
            DIN => \N__48614\,
            DOUT => \N__48613\,
            PACKAGEPIN => delay_tr_input_wire
        );

    \delay_tr_input_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48615\,
            PADOUT => \N__48614\,
            PADIN => \N__48613\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_tr_input_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48606\,
            DIN => \N__48605\,
            DOUT => \N__48604\,
            PACKAGEPIN => il_min_comp2_wire
        );

    \il_min_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48606\,
            PADOUT => \N__48605\,
            PADIN => \N__48604\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s1_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48597\,
            DIN => \N__48596\,
            DOUT => \N__48595\,
            PACKAGEPIN => s1_phy_wire
        );

    \s1_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48597\,
            PADOUT => \N__48596\,
            PADIN => \N__48595\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__32327\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s4_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48588\,
            DIN => \N__48587\,
            DOUT => \N__48586\,
            PACKAGEPIN => s4_phy_wire
        );

    \s4_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48588\,
            PADOUT => \N__48587\,
            PADIN => \N__48586\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__33641\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48579\,
            DIN => \N__48578\,
            DOUT => \N__48577\,
            PACKAGEPIN => il_min_comp1_wire
        );

    \il_min_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48579\,
            PADOUT => \N__48578\,
            PADIN => \N__48577\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s3_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48570\,
            DIN => \N__48569\,
            DOUT => \N__48568\,
            PACKAGEPIN => s3_phy_wire
        );

    \s3_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48570\,
            PADOUT => \N__48569\,
            PADIN => \N__48568\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__33902\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__11621\ : InMux
    port map (
            O => \N__48551\,
            I => \N__48547\
        );

    \I__11620\ : InMux
    port map (
            O => \N__48550\,
            I => \N__48544\
        );

    \I__11619\ : LocalMux
    port map (
            O => \N__48547\,
            I => \N__48538\
        );

    \I__11618\ : LocalMux
    port map (
            O => \N__48544\,
            I => \N__48538\
        );

    \I__11617\ : InMux
    port map (
            O => \N__48543\,
            I => \N__48535\
        );

    \I__11616\ : Span4Mux_v
    port map (
            O => \N__48538\,
            I => \N__48532\
        );

    \I__11615\ : LocalMux
    port map (
            O => \N__48535\,
            I => \N__48529\
        );

    \I__11614\ : Odrv4
    port map (
            O => \N__48532\,
            I => \delay_measurement_inst.elapsed_time_tr_16\
        );

    \I__11613\ : Odrv4
    port map (
            O => \N__48529\,
            I => \delay_measurement_inst.elapsed_time_tr_16\
        );

    \I__11612\ : InMux
    port map (
            O => \N__48524\,
            I => \N__48521\
        );

    \I__11611\ : LocalMux
    port map (
            O => \N__48521\,
            I => \N__48517\
        );

    \I__11610\ : InMux
    port map (
            O => \N__48520\,
            I => \N__48514\
        );

    \I__11609\ : Span4Mux_v
    port map (
            O => \N__48517\,
            I => \N__48509\
        );

    \I__11608\ : LocalMux
    port map (
            O => \N__48514\,
            I => \N__48509\
        );

    \I__11607\ : Odrv4
    port map (
            O => \N__48509\,
            I => \delay_measurement_inst.elapsed_time_tr_11\
        );

    \I__11606\ : InMux
    port map (
            O => \N__48506\,
            I => \N__48499\
        );

    \I__11605\ : InMux
    port map (
            O => \N__48505\,
            I => \N__48499\
        );

    \I__11604\ : InMux
    port map (
            O => \N__48504\,
            I => \N__48496\
        );

    \I__11603\ : LocalMux
    port map (
            O => \N__48499\,
            I => \N__48491\
        );

    \I__11602\ : LocalMux
    port map (
            O => \N__48496\,
            I => \N__48488\
        );

    \I__11601\ : InMux
    port map (
            O => \N__48495\,
            I => \N__48485\
        );

    \I__11600\ : InMux
    port map (
            O => \N__48494\,
            I => \N__48482\
        );

    \I__11599\ : Span4Mux_h
    port map (
            O => \N__48491\,
            I => \N__48479\
        );

    \I__11598\ : Span4Mux_h
    port map (
            O => \N__48488\,
            I => \N__48472\
        );

    \I__11597\ : LocalMux
    port map (
            O => \N__48485\,
            I => \N__48472\
        );

    \I__11596\ : LocalMux
    port map (
            O => \N__48482\,
            I => \N__48472\
        );

    \I__11595\ : Odrv4
    port map (
            O => \N__48479\,
            I => \delay_measurement_inst.N_301\
        );

    \I__11594\ : Odrv4
    port map (
            O => \N__48472\,
            I => \delay_measurement_inst.N_301\
        );

    \I__11593\ : InMux
    port map (
            O => \N__48467\,
            I => \N__48463\
        );

    \I__11592\ : InMux
    port map (
            O => \N__48466\,
            I => \N__48460\
        );

    \I__11591\ : LocalMux
    port map (
            O => \N__48463\,
            I => \N__48454\
        );

    \I__11590\ : LocalMux
    port map (
            O => \N__48460\,
            I => \N__48454\
        );

    \I__11589\ : InMux
    port map (
            O => \N__48459\,
            I => \N__48451\
        );

    \I__11588\ : Span12Mux_s10_v
    port map (
            O => \N__48454\,
            I => \N__48446\
        );

    \I__11587\ : LocalMux
    port map (
            O => \N__48451\,
            I => \N__48446\
        );

    \I__11586\ : Odrv12
    port map (
            O => \N__48446\,
            I => measured_delay_tr_11
        );

    \I__11585\ : InMux
    port map (
            O => \N__48443\,
            I => \N__48439\
        );

    \I__11584\ : InMux
    port map (
            O => \N__48442\,
            I => \N__48435\
        );

    \I__11583\ : LocalMux
    port map (
            O => \N__48439\,
            I => \N__48432\
        );

    \I__11582\ : InMux
    port map (
            O => \N__48438\,
            I => \N__48429\
        );

    \I__11581\ : LocalMux
    port map (
            O => \N__48435\,
            I => \N__48426\
        );

    \I__11580\ : Span4Mux_v
    port map (
            O => \N__48432\,
            I => \N__48423\
        );

    \I__11579\ : LocalMux
    port map (
            O => \N__48429\,
            I => \N__48420\
        );

    \I__11578\ : Span4Mux_h
    port map (
            O => \N__48426\,
            I => \N__48417\
        );

    \I__11577\ : Odrv4
    port map (
            O => \N__48423\,
            I => \delay_measurement_inst.elapsed_time_tr_18\
        );

    \I__11576\ : Odrv12
    port map (
            O => \N__48420\,
            I => \delay_measurement_inst.elapsed_time_tr_18\
        );

    \I__11575\ : Odrv4
    port map (
            O => \N__48417\,
            I => \delay_measurement_inst.elapsed_time_tr_18\
        );

    \I__11574\ : InMux
    port map (
            O => \N__48410\,
            I => \N__48406\
        );

    \I__11573\ : InMux
    port map (
            O => \N__48409\,
            I => \N__48403\
        );

    \I__11572\ : LocalMux
    port map (
            O => \N__48406\,
            I => \N__48397\
        );

    \I__11571\ : LocalMux
    port map (
            O => \N__48403\,
            I => \N__48397\
        );

    \I__11570\ : InMux
    port map (
            O => \N__48402\,
            I => \N__48394\
        );

    \I__11569\ : Span4Mux_v
    port map (
            O => \N__48397\,
            I => \N__48389\
        );

    \I__11568\ : LocalMux
    port map (
            O => \N__48394\,
            I => \N__48389\
        );

    \I__11567\ : Span4Mux_h
    port map (
            O => \N__48389\,
            I => \N__48385\
        );

    \I__11566\ : InMux
    port map (
            O => \N__48388\,
            I => \N__48382\
        );

    \I__11565\ : Odrv4
    port map (
            O => \N__48385\,
            I => measured_delay_tr_18
        );

    \I__11564\ : LocalMux
    port map (
            O => \N__48382\,
            I => measured_delay_tr_18
        );

    \I__11563\ : InMux
    port map (
            O => \N__48377\,
            I => \N__48374\
        );

    \I__11562\ : LocalMux
    port map (
            O => \N__48374\,
            I => \N__48370\
        );

    \I__11561\ : InMux
    port map (
            O => \N__48373\,
            I => \N__48367\
        );

    \I__11560\ : Span4Mux_v
    port map (
            O => \N__48370\,
            I => \N__48361\
        );

    \I__11559\ : LocalMux
    port map (
            O => \N__48367\,
            I => \N__48361\
        );

    \I__11558\ : InMux
    port map (
            O => \N__48366\,
            I => \N__48358\
        );

    \I__11557\ : Span4Mux_h
    port map (
            O => \N__48361\,
            I => \N__48352\
        );

    \I__11556\ : LocalMux
    port map (
            O => \N__48358\,
            I => \N__48352\
        );

    \I__11555\ : InMux
    port map (
            O => \N__48357\,
            I => \N__48349\
        );

    \I__11554\ : Span4Mux_v
    port map (
            O => \N__48352\,
            I => \N__48346\
        );

    \I__11553\ : LocalMux
    port map (
            O => \N__48349\,
            I => \N__48343\
        );

    \I__11552\ : Odrv4
    port map (
            O => \N__48346\,
            I => measured_delay_tr_17
        );

    \I__11551\ : Odrv4
    port map (
            O => \N__48343\,
            I => measured_delay_tr_17
        );

    \I__11550\ : InMux
    port map (
            O => \N__48338\,
            I => \N__48335\
        );

    \I__11549\ : LocalMux
    port map (
            O => \N__48335\,
            I => \N__48331\
        );

    \I__11548\ : InMux
    port map (
            O => \N__48334\,
            I => \N__48328\
        );

    \I__11547\ : Span4Mux_v
    port map (
            O => \N__48331\,
            I => \N__48322\
        );

    \I__11546\ : LocalMux
    port map (
            O => \N__48328\,
            I => \N__48322\
        );

    \I__11545\ : InMux
    port map (
            O => \N__48327\,
            I => \N__48319\
        );

    \I__11544\ : Span4Mux_h
    port map (
            O => \N__48322\,
            I => \N__48313\
        );

    \I__11543\ : LocalMux
    port map (
            O => \N__48319\,
            I => \N__48313\
        );

    \I__11542\ : InMux
    port map (
            O => \N__48318\,
            I => \N__48310\
        );

    \I__11541\ : Span4Mux_h
    port map (
            O => \N__48313\,
            I => \N__48307\
        );

    \I__11540\ : LocalMux
    port map (
            O => \N__48310\,
            I => \N__48304\
        );

    \I__11539\ : Odrv4
    port map (
            O => \N__48307\,
            I => measured_delay_tr_16
        );

    \I__11538\ : Odrv4
    port map (
            O => \N__48304\,
            I => measured_delay_tr_16
        );

    \I__11537\ : InMux
    port map (
            O => \N__48299\,
            I => \N__48296\
        );

    \I__11536\ : LocalMux
    port map (
            O => \N__48296\,
            I => \N__48293\
        );

    \I__11535\ : Odrv4
    port map (
            O => \N__48293\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3Z0Z_3\
        );

    \I__11534\ : InMux
    port map (
            O => \N__48290\,
            I => \N__48287\
        );

    \I__11533\ : LocalMux
    port map (
            O => \N__48287\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_i\
        );

    \I__11532\ : CascadeMux
    port map (
            O => \N__48284\,
            I => \N__48275\
        );

    \I__11531\ : CascadeMux
    port map (
            O => \N__48283\,
            I => \N__48270\
        );

    \I__11530\ : CascadeMux
    port map (
            O => \N__48282\,
            I => \N__48267\
        );

    \I__11529\ : CascadeMux
    port map (
            O => \N__48281\,
            I => \N__48262\
        );

    \I__11528\ : InMux
    port map (
            O => \N__48280\,
            I => \N__48254\
        );

    \I__11527\ : InMux
    port map (
            O => \N__48279\,
            I => \N__48247\
        );

    \I__11526\ : InMux
    port map (
            O => \N__48278\,
            I => \N__48247\
        );

    \I__11525\ : InMux
    port map (
            O => \N__48275\,
            I => \N__48240\
        );

    \I__11524\ : InMux
    port map (
            O => \N__48274\,
            I => \N__48240\
        );

    \I__11523\ : InMux
    port map (
            O => \N__48273\,
            I => \N__48240\
        );

    \I__11522\ : InMux
    port map (
            O => \N__48270\,
            I => \N__48231\
        );

    \I__11521\ : InMux
    port map (
            O => \N__48267\,
            I => \N__48231\
        );

    \I__11520\ : InMux
    port map (
            O => \N__48266\,
            I => \N__48231\
        );

    \I__11519\ : InMux
    port map (
            O => \N__48265\,
            I => \N__48231\
        );

    \I__11518\ : InMux
    port map (
            O => \N__48262\,
            I => \N__48228\
        );

    \I__11517\ : InMux
    port map (
            O => \N__48261\,
            I => \N__48223\
        );

    \I__11516\ : InMux
    port map (
            O => \N__48260\,
            I => \N__48223\
        );

    \I__11515\ : CascadeMux
    port map (
            O => \N__48259\,
            I => \N__48220\
        );

    \I__11514\ : CascadeMux
    port map (
            O => \N__48258\,
            I => \N__48217\
        );

    \I__11513\ : CascadeMux
    port map (
            O => \N__48257\,
            I => \N__48212\
        );

    \I__11512\ : LocalMux
    port map (
            O => \N__48254\,
            I => \N__48208\
        );

    \I__11511\ : InMux
    port map (
            O => \N__48253\,
            I => \N__48203\
        );

    \I__11510\ : InMux
    port map (
            O => \N__48252\,
            I => \N__48203\
        );

    \I__11509\ : LocalMux
    port map (
            O => \N__48247\,
            I => \N__48196\
        );

    \I__11508\ : LocalMux
    port map (
            O => \N__48240\,
            I => \N__48196\
        );

    \I__11507\ : LocalMux
    port map (
            O => \N__48231\,
            I => \N__48196\
        );

    \I__11506\ : LocalMux
    port map (
            O => \N__48228\,
            I => \N__48191\
        );

    \I__11505\ : LocalMux
    port map (
            O => \N__48223\,
            I => \N__48191\
        );

    \I__11504\ : InMux
    port map (
            O => \N__48220\,
            I => \N__48178\
        );

    \I__11503\ : InMux
    port map (
            O => \N__48217\,
            I => \N__48178\
        );

    \I__11502\ : InMux
    port map (
            O => \N__48216\,
            I => \N__48178\
        );

    \I__11501\ : InMux
    port map (
            O => \N__48215\,
            I => \N__48178\
        );

    \I__11500\ : InMux
    port map (
            O => \N__48212\,
            I => \N__48178\
        );

    \I__11499\ : InMux
    port map (
            O => \N__48211\,
            I => \N__48178\
        );

    \I__11498\ : Span4Mux_v
    port map (
            O => \N__48208\,
            I => \N__48173\
        );

    \I__11497\ : LocalMux
    port map (
            O => \N__48203\,
            I => \N__48173\
        );

    \I__11496\ : Span4Mux_v
    port map (
            O => \N__48196\,
            I => \N__48168\
        );

    \I__11495\ : Span4Mux_v
    port map (
            O => \N__48191\,
            I => \N__48168\
        );

    \I__11494\ : LocalMux
    port map (
            O => \N__48178\,
            I => \N__48165\
        );

    \I__11493\ : Span4Mux_h
    port map (
            O => \N__48173\,
            I => \N__48162\
        );

    \I__11492\ : Odrv4
    port map (
            O => \N__48168\,
            I => \delay_measurement_inst.elapsed_time_tr_31\
        );

    \I__11491\ : Odrv12
    port map (
            O => \N__48165\,
            I => \delay_measurement_inst.elapsed_time_tr_31\
        );

    \I__11490\ : Odrv4
    port map (
            O => \N__48162\,
            I => \delay_measurement_inst.elapsed_time_tr_31\
        );

    \I__11489\ : InMux
    port map (
            O => \N__48155\,
            I => \N__48151\
        );

    \I__11488\ : InMux
    port map (
            O => \N__48154\,
            I => \N__48148\
        );

    \I__11487\ : LocalMux
    port map (
            O => \N__48151\,
            I => \N__48144\
        );

    \I__11486\ : LocalMux
    port map (
            O => \N__48148\,
            I => \N__48141\
        );

    \I__11485\ : CascadeMux
    port map (
            O => \N__48147\,
            I => \N__48138\
        );

    \I__11484\ : Span4Mux_v
    port map (
            O => \N__48144\,
            I => \N__48133\
        );

    \I__11483\ : Span4Mux_v
    port map (
            O => \N__48141\,
            I => \N__48133\
        );

    \I__11482\ : InMux
    port map (
            O => \N__48138\,
            I => \N__48130\
        );

    \I__11481\ : Sp12to4
    port map (
            O => \N__48133\,
            I => \N__48125\
        );

    \I__11480\ : LocalMux
    port map (
            O => \N__48130\,
            I => \N__48125\
        );

    \I__11479\ : Odrv12
    port map (
            O => \N__48125\,
            I => \delay_measurement_inst.elapsed_time_tr_19\
        );

    \I__11478\ : InMux
    port map (
            O => \N__48122\,
            I => \N__48114\
        );

    \I__11477\ : InMux
    port map (
            O => \N__48121\,
            I => \N__48114\
        );

    \I__11476\ : InMux
    port map (
            O => \N__48120\,
            I => \N__48111\
        );

    \I__11475\ : InMux
    port map (
            O => \N__48119\,
            I => \N__48108\
        );

    \I__11474\ : LocalMux
    port map (
            O => \N__48114\,
            I => \N__48103\
        );

    \I__11473\ : LocalMux
    port map (
            O => \N__48111\,
            I => \N__48100\
        );

    \I__11472\ : LocalMux
    port map (
            O => \N__48108\,
            I => \N__48097\
        );

    \I__11471\ : InMux
    port map (
            O => \N__48107\,
            I => \N__48092\
        );

    \I__11470\ : InMux
    port map (
            O => \N__48106\,
            I => \N__48092\
        );

    \I__11469\ : Span4Mux_v
    port map (
            O => \N__48103\,
            I => \N__48081\
        );

    \I__11468\ : Span4Mux_h
    port map (
            O => \N__48100\,
            I => \N__48081\
        );

    \I__11467\ : Span4Mux_v
    port map (
            O => \N__48097\,
            I => \N__48081\
        );

    \I__11466\ : LocalMux
    port map (
            O => \N__48092\,
            I => \N__48081\
        );

    \I__11465\ : InMux
    port map (
            O => \N__48091\,
            I => \N__48075\
        );

    \I__11464\ : InMux
    port map (
            O => \N__48090\,
            I => \N__48075\
        );

    \I__11463\ : Span4Mux_h
    port map (
            O => \N__48081\,
            I => \N__48072\
        );

    \I__11462\ : InMux
    port map (
            O => \N__48080\,
            I => \N__48069\
        );

    \I__11461\ : LocalMux
    port map (
            O => \N__48075\,
            I => \N__48066\
        );

    \I__11460\ : Odrv4
    port map (
            O => \N__48072\,
            I => \delay_measurement_inst.N_358\
        );

    \I__11459\ : LocalMux
    port map (
            O => \N__48069\,
            I => \delay_measurement_inst.N_358\
        );

    \I__11458\ : Odrv12
    port map (
            O => \N__48066\,
            I => \delay_measurement_inst.N_358\
        );

    \I__11457\ : InMux
    port map (
            O => \N__48059\,
            I => \N__48056\
        );

    \I__11456\ : LocalMux
    port map (
            O => \N__48056\,
            I => \N__48051\
        );

    \I__11455\ : CascadeMux
    port map (
            O => \N__48055\,
            I => \N__48048\
        );

    \I__11454\ : InMux
    port map (
            O => \N__48054\,
            I => \N__48045\
        );

    \I__11453\ : Span4Mux_v
    port map (
            O => \N__48051\,
            I => \N__48041\
        );

    \I__11452\ : InMux
    port map (
            O => \N__48048\,
            I => \N__48038\
        );

    \I__11451\ : LocalMux
    port map (
            O => \N__48045\,
            I => \N__48035\
        );

    \I__11450\ : CascadeMux
    port map (
            O => \N__48044\,
            I => \N__48032\
        );

    \I__11449\ : Span4Mux_h
    port map (
            O => \N__48041\,
            I => \N__48027\
        );

    \I__11448\ : LocalMux
    port map (
            O => \N__48038\,
            I => \N__48027\
        );

    \I__11447\ : Span4Mux_v
    port map (
            O => \N__48035\,
            I => \N__48024\
        );

    \I__11446\ : InMux
    port map (
            O => \N__48032\,
            I => \N__48021\
        );

    \I__11445\ : Span4Mux_v
    port map (
            O => \N__48027\,
            I => \N__48018\
        );

    \I__11444\ : Span4Mux_h
    port map (
            O => \N__48024\,
            I => \N__48013\
        );

    \I__11443\ : LocalMux
    port map (
            O => \N__48021\,
            I => \N__48013\
        );

    \I__11442\ : Odrv4
    port map (
            O => \N__48018\,
            I => measured_delay_tr_19
        );

    \I__11441\ : Odrv4
    port map (
            O => \N__48013\,
            I => measured_delay_tr_19
        );

    \I__11440\ : ClkMux
    port map (
            O => \N__48008\,
            I => \N__47522\
        );

    \I__11439\ : ClkMux
    port map (
            O => \N__48007\,
            I => \N__47522\
        );

    \I__11438\ : ClkMux
    port map (
            O => \N__48006\,
            I => \N__47522\
        );

    \I__11437\ : ClkMux
    port map (
            O => \N__48005\,
            I => \N__47522\
        );

    \I__11436\ : ClkMux
    port map (
            O => \N__48004\,
            I => \N__47522\
        );

    \I__11435\ : ClkMux
    port map (
            O => \N__48003\,
            I => \N__47522\
        );

    \I__11434\ : ClkMux
    port map (
            O => \N__48002\,
            I => \N__47522\
        );

    \I__11433\ : ClkMux
    port map (
            O => \N__48001\,
            I => \N__47522\
        );

    \I__11432\ : ClkMux
    port map (
            O => \N__48000\,
            I => \N__47522\
        );

    \I__11431\ : ClkMux
    port map (
            O => \N__47999\,
            I => \N__47522\
        );

    \I__11430\ : ClkMux
    port map (
            O => \N__47998\,
            I => \N__47522\
        );

    \I__11429\ : ClkMux
    port map (
            O => \N__47997\,
            I => \N__47522\
        );

    \I__11428\ : ClkMux
    port map (
            O => \N__47996\,
            I => \N__47522\
        );

    \I__11427\ : ClkMux
    port map (
            O => \N__47995\,
            I => \N__47522\
        );

    \I__11426\ : ClkMux
    port map (
            O => \N__47994\,
            I => \N__47522\
        );

    \I__11425\ : ClkMux
    port map (
            O => \N__47993\,
            I => \N__47522\
        );

    \I__11424\ : ClkMux
    port map (
            O => \N__47992\,
            I => \N__47522\
        );

    \I__11423\ : ClkMux
    port map (
            O => \N__47991\,
            I => \N__47522\
        );

    \I__11422\ : ClkMux
    port map (
            O => \N__47990\,
            I => \N__47522\
        );

    \I__11421\ : ClkMux
    port map (
            O => \N__47989\,
            I => \N__47522\
        );

    \I__11420\ : ClkMux
    port map (
            O => \N__47988\,
            I => \N__47522\
        );

    \I__11419\ : ClkMux
    port map (
            O => \N__47987\,
            I => \N__47522\
        );

    \I__11418\ : ClkMux
    port map (
            O => \N__47986\,
            I => \N__47522\
        );

    \I__11417\ : ClkMux
    port map (
            O => \N__47985\,
            I => \N__47522\
        );

    \I__11416\ : ClkMux
    port map (
            O => \N__47984\,
            I => \N__47522\
        );

    \I__11415\ : ClkMux
    port map (
            O => \N__47983\,
            I => \N__47522\
        );

    \I__11414\ : ClkMux
    port map (
            O => \N__47982\,
            I => \N__47522\
        );

    \I__11413\ : ClkMux
    port map (
            O => \N__47981\,
            I => \N__47522\
        );

    \I__11412\ : ClkMux
    port map (
            O => \N__47980\,
            I => \N__47522\
        );

    \I__11411\ : ClkMux
    port map (
            O => \N__47979\,
            I => \N__47522\
        );

    \I__11410\ : ClkMux
    port map (
            O => \N__47978\,
            I => \N__47522\
        );

    \I__11409\ : ClkMux
    port map (
            O => \N__47977\,
            I => \N__47522\
        );

    \I__11408\ : ClkMux
    port map (
            O => \N__47976\,
            I => \N__47522\
        );

    \I__11407\ : ClkMux
    port map (
            O => \N__47975\,
            I => \N__47522\
        );

    \I__11406\ : ClkMux
    port map (
            O => \N__47974\,
            I => \N__47522\
        );

    \I__11405\ : ClkMux
    port map (
            O => \N__47973\,
            I => \N__47522\
        );

    \I__11404\ : ClkMux
    port map (
            O => \N__47972\,
            I => \N__47522\
        );

    \I__11403\ : ClkMux
    port map (
            O => \N__47971\,
            I => \N__47522\
        );

    \I__11402\ : ClkMux
    port map (
            O => \N__47970\,
            I => \N__47522\
        );

    \I__11401\ : ClkMux
    port map (
            O => \N__47969\,
            I => \N__47522\
        );

    \I__11400\ : ClkMux
    port map (
            O => \N__47968\,
            I => \N__47522\
        );

    \I__11399\ : ClkMux
    port map (
            O => \N__47967\,
            I => \N__47522\
        );

    \I__11398\ : ClkMux
    port map (
            O => \N__47966\,
            I => \N__47522\
        );

    \I__11397\ : ClkMux
    port map (
            O => \N__47965\,
            I => \N__47522\
        );

    \I__11396\ : ClkMux
    port map (
            O => \N__47964\,
            I => \N__47522\
        );

    \I__11395\ : ClkMux
    port map (
            O => \N__47963\,
            I => \N__47522\
        );

    \I__11394\ : ClkMux
    port map (
            O => \N__47962\,
            I => \N__47522\
        );

    \I__11393\ : ClkMux
    port map (
            O => \N__47961\,
            I => \N__47522\
        );

    \I__11392\ : ClkMux
    port map (
            O => \N__47960\,
            I => \N__47522\
        );

    \I__11391\ : ClkMux
    port map (
            O => \N__47959\,
            I => \N__47522\
        );

    \I__11390\ : ClkMux
    port map (
            O => \N__47958\,
            I => \N__47522\
        );

    \I__11389\ : ClkMux
    port map (
            O => \N__47957\,
            I => \N__47522\
        );

    \I__11388\ : ClkMux
    port map (
            O => \N__47956\,
            I => \N__47522\
        );

    \I__11387\ : ClkMux
    port map (
            O => \N__47955\,
            I => \N__47522\
        );

    \I__11386\ : ClkMux
    port map (
            O => \N__47954\,
            I => \N__47522\
        );

    \I__11385\ : ClkMux
    port map (
            O => \N__47953\,
            I => \N__47522\
        );

    \I__11384\ : ClkMux
    port map (
            O => \N__47952\,
            I => \N__47522\
        );

    \I__11383\ : ClkMux
    port map (
            O => \N__47951\,
            I => \N__47522\
        );

    \I__11382\ : ClkMux
    port map (
            O => \N__47950\,
            I => \N__47522\
        );

    \I__11381\ : ClkMux
    port map (
            O => \N__47949\,
            I => \N__47522\
        );

    \I__11380\ : ClkMux
    port map (
            O => \N__47948\,
            I => \N__47522\
        );

    \I__11379\ : ClkMux
    port map (
            O => \N__47947\,
            I => \N__47522\
        );

    \I__11378\ : ClkMux
    port map (
            O => \N__47946\,
            I => \N__47522\
        );

    \I__11377\ : ClkMux
    port map (
            O => \N__47945\,
            I => \N__47522\
        );

    \I__11376\ : ClkMux
    port map (
            O => \N__47944\,
            I => \N__47522\
        );

    \I__11375\ : ClkMux
    port map (
            O => \N__47943\,
            I => \N__47522\
        );

    \I__11374\ : ClkMux
    port map (
            O => \N__47942\,
            I => \N__47522\
        );

    \I__11373\ : ClkMux
    port map (
            O => \N__47941\,
            I => \N__47522\
        );

    \I__11372\ : ClkMux
    port map (
            O => \N__47940\,
            I => \N__47522\
        );

    \I__11371\ : ClkMux
    port map (
            O => \N__47939\,
            I => \N__47522\
        );

    \I__11370\ : ClkMux
    port map (
            O => \N__47938\,
            I => \N__47522\
        );

    \I__11369\ : ClkMux
    port map (
            O => \N__47937\,
            I => \N__47522\
        );

    \I__11368\ : ClkMux
    port map (
            O => \N__47936\,
            I => \N__47522\
        );

    \I__11367\ : ClkMux
    port map (
            O => \N__47935\,
            I => \N__47522\
        );

    \I__11366\ : ClkMux
    port map (
            O => \N__47934\,
            I => \N__47522\
        );

    \I__11365\ : ClkMux
    port map (
            O => \N__47933\,
            I => \N__47522\
        );

    \I__11364\ : ClkMux
    port map (
            O => \N__47932\,
            I => \N__47522\
        );

    \I__11363\ : ClkMux
    port map (
            O => \N__47931\,
            I => \N__47522\
        );

    \I__11362\ : ClkMux
    port map (
            O => \N__47930\,
            I => \N__47522\
        );

    \I__11361\ : ClkMux
    port map (
            O => \N__47929\,
            I => \N__47522\
        );

    \I__11360\ : ClkMux
    port map (
            O => \N__47928\,
            I => \N__47522\
        );

    \I__11359\ : ClkMux
    port map (
            O => \N__47927\,
            I => \N__47522\
        );

    \I__11358\ : ClkMux
    port map (
            O => \N__47926\,
            I => \N__47522\
        );

    \I__11357\ : ClkMux
    port map (
            O => \N__47925\,
            I => \N__47522\
        );

    \I__11356\ : ClkMux
    port map (
            O => \N__47924\,
            I => \N__47522\
        );

    \I__11355\ : ClkMux
    port map (
            O => \N__47923\,
            I => \N__47522\
        );

    \I__11354\ : ClkMux
    port map (
            O => \N__47922\,
            I => \N__47522\
        );

    \I__11353\ : ClkMux
    port map (
            O => \N__47921\,
            I => \N__47522\
        );

    \I__11352\ : ClkMux
    port map (
            O => \N__47920\,
            I => \N__47522\
        );

    \I__11351\ : ClkMux
    port map (
            O => \N__47919\,
            I => \N__47522\
        );

    \I__11350\ : ClkMux
    port map (
            O => \N__47918\,
            I => \N__47522\
        );

    \I__11349\ : ClkMux
    port map (
            O => \N__47917\,
            I => \N__47522\
        );

    \I__11348\ : ClkMux
    port map (
            O => \N__47916\,
            I => \N__47522\
        );

    \I__11347\ : ClkMux
    port map (
            O => \N__47915\,
            I => \N__47522\
        );

    \I__11346\ : ClkMux
    port map (
            O => \N__47914\,
            I => \N__47522\
        );

    \I__11345\ : ClkMux
    port map (
            O => \N__47913\,
            I => \N__47522\
        );

    \I__11344\ : ClkMux
    port map (
            O => \N__47912\,
            I => \N__47522\
        );

    \I__11343\ : ClkMux
    port map (
            O => \N__47911\,
            I => \N__47522\
        );

    \I__11342\ : ClkMux
    port map (
            O => \N__47910\,
            I => \N__47522\
        );

    \I__11341\ : ClkMux
    port map (
            O => \N__47909\,
            I => \N__47522\
        );

    \I__11340\ : ClkMux
    port map (
            O => \N__47908\,
            I => \N__47522\
        );

    \I__11339\ : ClkMux
    port map (
            O => \N__47907\,
            I => \N__47522\
        );

    \I__11338\ : ClkMux
    port map (
            O => \N__47906\,
            I => \N__47522\
        );

    \I__11337\ : ClkMux
    port map (
            O => \N__47905\,
            I => \N__47522\
        );

    \I__11336\ : ClkMux
    port map (
            O => \N__47904\,
            I => \N__47522\
        );

    \I__11335\ : ClkMux
    port map (
            O => \N__47903\,
            I => \N__47522\
        );

    \I__11334\ : ClkMux
    port map (
            O => \N__47902\,
            I => \N__47522\
        );

    \I__11333\ : ClkMux
    port map (
            O => \N__47901\,
            I => \N__47522\
        );

    \I__11332\ : ClkMux
    port map (
            O => \N__47900\,
            I => \N__47522\
        );

    \I__11331\ : ClkMux
    port map (
            O => \N__47899\,
            I => \N__47522\
        );

    \I__11330\ : ClkMux
    port map (
            O => \N__47898\,
            I => \N__47522\
        );

    \I__11329\ : ClkMux
    port map (
            O => \N__47897\,
            I => \N__47522\
        );

    \I__11328\ : ClkMux
    port map (
            O => \N__47896\,
            I => \N__47522\
        );

    \I__11327\ : ClkMux
    port map (
            O => \N__47895\,
            I => \N__47522\
        );

    \I__11326\ : ClkMux
    port map (
            O => \N__47894\,
            I => \N__47522\
        );

    \I__11325\ : ClkMux
    port map (
            O => \N__47893\,
            I => \N__47522\
        );

    \I__11324\ : ClkMux
    port map (
            O => \N__47892\,
            I => \N__47522\
        );

    \I__11323\ : ClkMux
    port map (
            O => \N__47891\,
            I => \N__47522\
        );

    \I__11322\ : ClkMux
    port map (
            O => \N__47890\,
            I => \N__47522\
        );

    \I__11321\ : ClkMux
    port map (
            O => \N__47889\,
            I => \N__47522\
        );

    \I__11320\ : ClkMux
    port map (
            O => \N__47888\,
            I => \N__47522\
        );

    \I__11319\ : ClkMux
    port map (
            O => \N__47887\,
            I => \N__47522\
        );

    \I__11318\ : ClkMux
    port map (
            O => \N__47886\,
            I => \N__47522\
        );

    \I__11317\ : ClkMux
    port map (
            O => \N__47885\,
            I => \N__47522\
        );

    \I__11316\ : ClkMux
    port map (
            O => \N__47884\,
            I => \N__47522\
        );

    \I__11315\ : ClkMux
    port map (
            O => \N__47883\,
            I => \N__47522\
        );

    \I__11314\ : ClkMux
    port map (
            O => \N__47882\,
            I => \N__47522\
        );

    \I__11313\ : ClkMux
    port map (
            O => \N__47881\,
            I => \N__47522\
        );

    \I__11312\ : ClkMux
    port map (
            O => \N__47880\,
            I => \N__47522\
        );

    \I__11311\ : ClkMux
    port map (
            O => \N__47879\,
            I => \N__47522\
        );

    \I__11310\ : ClkMux
    port map (
            O => \N__47878\,
            I => \N__47522\
        );

    \I__11309\ : ClkMux
    port map (
            O => \N__47877\,
            I => \N__47522\
        );

    \I__11308\ : ClkMux
    port map (
            O => \N__47876\,
            I => \N__47522\
        );

    \I__11307\ : ClkMux
    port map (
            O => \N__47875\,
            I => \N__47522\
        );

    \I__11306\ : ClkMux
    port map (
            O => \N__47874\,
            I => \N__47522\
        );

    \I__11305\ : ClkMux
    port map (
            O => \N__47873\,
            I => \N__47522\
        );

    \I__11304\ : ClkMux
    port map (
            O => \N__47872\,
            I => \N__47522\
        );

    \I__11303\ : ClkMux
    port map (
            O => \N__47871\,
            I => \N__47522\
        );

    \I__11302\ : ClkMux
    port map (
            O => \N__47870\,
            I => \N__47522\
        );

    \I__11301\ : ClkMux
    port map (
            O => \N__47869\,
            I => \N__47522\
        );

    \I__11300\ : ClkMux
    port map (
            O => \N__47868\,
            I => \N__47522\
        );

    \I__11299\ : ClkMux
    port map (
            O => \N__47867\,
            I => \N__47522\
        );

    \I__11298\ : ClkMux
    port map (
            O => \N__47866\,
            I => \N__47522\
        );

    \I__11297\ : ClkMux
    port map (
            O => \N__47865\,
            I => \N__47522\
        );

    \I__11296\ : ClkMux
    port map (
            O => \N__47864\,
            I => \N__47522\
        );

    \I__11295\ : ClkMux
    port map (
            O => \N__47863\,
            I => \N__47522\
        );

    \I__11294\ : ClkMux
    port map (
            O => \N__47862\,
            I => \N__47522\
        );

    \I__11293\ : ClkMux
    port map (
            O => \N__47861\,
            I => \N__47522\
        );

    \I__11292\ : ClkMux
    port map (
            O => \N__47860\,
            I => \N__47522\
        );

    \I__11291\ : ClkMux
    port map (
            O => \N__47859\,
            I => \N__47522\
        );

    \I__11290\ : ClkMux
    port map (
            O => \N__47858\,
            I => \N__47522\
        );

    \I__11289\ : ClkMux
    port map (
            O => \N__47857\,
            I => \N__47522\
        );

    \I__11288\ : ClkMux
    port map (
            O => \N__47856\,
            I => \N__47522\
        );

    \I__11287\ : ClkMux
    port map (
            O => \N__47855\,
            I => \N__47522\
        );

    \I__11286\ : ClkMux
    port map (
            O => \N__47854\,
            I => \N__47522\
        );

    \I__11285\ : ClkMux
    port map (
            O => \N__47853\,
            I => \N__47522\
        );

    \I__11284\ : ClkMux
    port map (
            O => \N__47852\,
            I => \N__47522\
        );

    \I__11283\ : ClkMux
    port map (
            O => \N__47851\,
            I => \N__47522\
        );

    \I__11282\ : ClkMux
    port map (
            O => \N__47850\,
            I => \N__47522\
        );

    \I__11281\ : ClkMux
    port map (
            O => \N__47849\,
            I => \N__47522\
        );

    \I__11280\ : ClkMux
    port map (
            O => \N__47848\,
            I => \N__47522\
        );

    \I__11279\ : ClkMux
    port map (
            O => \N__47847\,
            I => \N__47522\
        );

    \I__11278\ : GlobalMux
    port map (
            O => \N__47522\,
            I => clk_100mhz_0
        );

    \I__11277\ : CEMux
    port map (
            O => \N__47519\,
            I => \N__47515\
        );

    \I__11276\ : CEMux
    port map (
            O => \N__47518\,
            I => \N__47512\
        );

    \I__11275\ : LocalMux
    port map (
            O => \N__47515\,
            I => \N__47508\
        );

    \I__11274\ : LocalMux
    port map (
            O => \N__47512\,
            I => \N__47505\
        );

    \I__11273\ : CEMux
    port map (
            O => \N__47511\,
            I => \N__47502\
        );

    \I__11272\ : Span4Mux_v
    port map (
            O => \N__47508\,
            I => \N__47499\
        );

    \I__11271\ : Span4Mux_v
    port map (
            O => \N__47505\,
            I => \N__47496\
        );

    \I__11270\ : LocalMux
    port map (
            O => \N__47502\,
            I => \N__47493\
        );

    \I__11269\ : Span4Mux_h
    port map (
            O => \N__47499\,
            I => \N__47483\
        );

    \I__11268\ : Span4Mux_h
    port map (
            O => \N__47496\,
            I => \N__47483\
        );

    \I__11267\ : Span4Mux_v
    port map (
            O => \N__47493\,
            I => \N__47483\
        );

    \I__11266\ : CEMux
    port map (
            O => \N__47492\,
            I => \N__47480\
        );

    \I__11265\ : CEMux
    port map (
            O => \N__47491\,
            I => \N__47477\
        );

    \I__11264\ : CEMux
    port map (
            O => \N__47490\,
            I => \N__47474\
        );

    \I__11263\ : Odrv4
    port map (
            O => \N__47483\,
            I => \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\
        );

    \I__11262\ : LocalMux
    port map (
            O => \N__47480\,
            I => \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\
        );

    \I__11261\ : LocalMux
    port map (
            O => \N__47477\,
            I => \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\
        );

    \I__11260\ : LocalMux
    port map (
            O => \N__47474\,
            I => \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\
        );

    \I__11259\ : CascadeMux
    port map (
            O => \N__47465\,
            I => \N__47456\
        );

    \I__11258\ : CascadeMux
    port map (
            O => \N__47464\,
            I => \N__47453\
        );

    \I__11257\ : InMux
    port map (
            O => \N__47463\,
            I => \N__47450\
        );

    \I__11256\ : InMux
    port map (
            O => \N__47462\,
            I => \N__47447\
        );

    \I__11255\ : InMux
    port map (
            O => \N__47461\,
            I => \N__47444\
        );

    \I__11254\ : InMux
    port map (
            O => \N__47460\,
            I => \N__47441\
        );

    \I__11253\ : InMux
    port map (
            O => \N__47459\,
            I => \N__47438\
        );

    \I__11252\ : InMux
    port map (
            O => \N__47456\,
            I => \N__47435\
        );

    \I__11251\ : InMux
    port map (
            O => \N__47453\,
            I => \N__47432\
        );

    \I__11250\ : LocalMux
    port map (
            O => \N__47450\,
            I => \N__47429\
        );

    \I__11249\ : LocalMux
    port map (
            O => \N__47447\,
            I => \N__47426\
        );

    \I__11248\ : LocalMux
    port map (
            O => \N__47444\,
            I => \N__47423\
        );

    \I__11247\ : LocalMux
    port map (
            O => \N__47441\,
            I => \N__47418\
        );

    \I__11246\ : LocalMux
    port map (
            O => \N__47438\,
            I => \N__47332\
        );

    \I__11245\ : LocalMux
    port map (
            O => \N__47435\,
            I => \N__47283\
        );

    \I__11244\ : LocalMux
    port map (
            O => \N__47432\,
            I => \N__47280\
        );

    \I__11243\ : Glb2LocalMux
    port map (
            O => \N__47429\,
            I => \N__46979\
        );

    \I__11242\ : Glb2LocalMux
    port map (
            O => \N__47426\,
            I => \N__46979\
        );

    \I__11241\ : Glb2LocalMux
    port map (
            O => \N__47423\,
            I => \N__46979\
        );

    \I__11240\ : SRMux
    port map (
            O => \N__47422\,
            I => \N__46979\
        );

    \I__11239\ : SRMux
    port map (
            O => \N__47421\,
            I => \N__46979\
        );

    \I__11238\ : Glb2LocalMux
    port map (
            O => \N__47418\,
            I => \N__46979\
        );

    \I__11237\ : SRMux
    port map (
            O => \N__47417\,
            I => \N__46979\
        );

    \I__11236\ : SRMux
    port map (
            O => \N__47416\,
            I => \N__46979\
        );

    \I__11235\ : SRMux
    port map (
            O => \N__47415\,
            I => \N__46979\
        );

    \I__11234\ : SRMux
    port map (
            O => \N__47414\,
            I => \N__46979\
        );

    \I__11233\ : SRMux
    port map (
            O => \N__47413\,
            I => \N__46979\
        );

    \I__11232\ : SRMux
    port map (
            O => \N__47412\,
            I => \N__46979\
        );

    \I__11231\ : SRMux
    port map (
            O => \N__47411\,
            I => \N__46979\
        );

    \I__11230\ : SRMux
    port map (
            O => \N__47410\,
            I => \N__46979\
        );

    \I__11229\ : SRMux
    port map (
            O => \N__47409\,
            I => \N__46979\
        );

    \I__11228\ : SRMux
    port map (
            O => \N__47408\,
            I => \N__46979\
        );

    \I__11227\ : SRMux
    port map (
            O => \N__47407\,
            I => \N__46979\
        );

    \I__11226\ : SRMux
    port map (
            O => \N__47406\,
            I => \N__46979\
        );

    \I__11225\ : SRMux
    port map (
            O => \N__47405\,
            I => \N__46979\
        );

    \I__11224\ : SRMux
    port map (
            O => \N__47404\,
            I => \N__46979\
        );

    \I__11223\ : SRMux
    port map (
            O => \N__47403\,
            I => \N__46979\
        );

    \I__11222\ : SRMux
    port map (
            O => \N__47402\,
            I => \N__46979\
        );

    \I__11221\ : SRMux
    port map (
            O => \N__47401\,
            I => \N__46979\
        );

    \I__11220\ : SRMux
    port map (
            O => \N__47400\,
            I => \N__46979\
        );

    \I__11219\ : SRMux
    port map (
            O => \N__47399\,
            I => \N__46979\
        );

    \I__11218\ : SRMux
    port map (
            O => \N__47398\,
            I => \N__46979\
        );

    \I__11217\ : SRMux
    port map (
            O => \N__47397\,
            I => \N__46979\
        );

    \I__11216\ : SRMux
    port map (
            O => \N__47396\,
            I => \N__46979\
        );

    \I__11215\ : SRMux
    port map (
            O => \N__47395\,
            I => \N__46979\
        );

    \I__11214\ : SRMux
    port map (
            O => \N__47394\,
            I => \N__46979\
        );

    \I__11213\ : SRMux
    port map (
            O => \N__47393\,
            I => \N__46979\
        );

    \I__11212\ : SRMux
    port map (
            O => \N__47392\,
            I => \N__46979\
        );

    \I__11211\ : SRMux
    port map (
            O => \N__47391\,
            I => \N__46979\
        );

    \I__11210\ : SRMux
    port map (
            O => \N__47390\,
            I => \N__46979\
        );

    \I__11209\ : SRMux
    port map (
            O => \N__47389\,
            I => \N__46979\
        );

    \I__11208\ : SRMux
    port map (
            O => \N__47388\,
            I => \N__46979\
        );

    \I__11207\ : SRMux
    port map (
            O => \N__47387\,
            I => \N__46979\
        );

    \I__11206\ : SRMux
    port map (
            O => \N__47386\,
            I => \N__46979\
        );

    \I__11205\ : SRMux
    port map (
            O => \N__47385\,
            I => \N__46979\
        );

    \I__11204\ : SRMux
    port map (
            O => \N__47384\,
            I => \N__46979\
        );

    \I__11203\ : SRMux
    port map (
            O => \N__47383\,
            I => \N__46979\
        );

    \I__11202\ : SRMux
    port map (
            O => \N__47382\,
            I => \N__46979\
        );

    \I__11201\ : SRMux
    port map (
            O => \N__47381\,
            I => \N__46979\
        );

    \I__11200\ : SRMux
    port map (
            O => \N__47380\,
            I => \N__46979\
        );

    \I__11199\ : SRMux
    port map (
            O => \N__47379\,
            I => \N__46979\
        );

    \I__11198\ : SRMux
    port map (
            O => \N__47378\,
            I => \N__46979\
        );

    \I__11197\ : SRMux
    port map (
            O => \N__47377\,
            I => \N__46979\
        );

    \I__11196\ : SRMux
    port map (
            O => \N__47376\,
            I => \N__46979\
        );

    \I__11195\ : SRMux
    port map (
            O => \N__47375\,
            I => \N__46979\
        );

    \I__11194\ : SRMux
    port map (
            O => \N__47374\,
            I => \N__46979\
        );

    \I__11193\ : SRMux
    port map (
            O => \N__47373\,
            I => \N__46979\
        );

    \I__11192\ : SRMux
    port map (
            O => \N__47372\,
            I => \N__46979\
        );

    \I__11191\ : SRMux
    port map (
            O => \N__47371\,
            I => \N__46979\
        );

    \I__11190\ : SRMux
    port map (
            O => \N__47370\,
            I => \N__46979\
        );

    \I__11189\ : SRMux
    port map (
            O => \N__47369\,
            I => \N__46979\
        );

    \I__11188\ : SRMux
    port map (
            O => \N__47368\,
            I => \N__46979\
        );

    \I__11187\ : SRMux
    port map (
            O => \N__47367\,
            I => \N__46979\
        );

    \I__11186\ : SRMux
    port map (
            O => \N__47366\,
            I => \N__46979\
        );

    \I__11185\ : SRMux
    port map (
            O => \N__47365\,
            I => \N__46979\
        );

    \I__11184\ : SRMux
    port map (
            O => \N__47364\,
            I => \N__46979\
        );

    \I__11183\ : SRMux
    port map (
            O => \N__47363\,
            I => \N__46979\
        );

    \I__11182\ : SRMux
    port map (
            O => \N__47362\,
            I => \N__46979\
        );

    \I__11181\ : SRMux
    port map (
            O => \N__47361\,
            I => \N__46979\
        );

    \I__11180\ : SRMux
    port map (
            O => \N__47360\,
            I => \N__46979\
        );

    \I__11179\ : SRMux
    port map (
            O => \N__47359\,
            I => \N__46979\
        );

    \I__11178\ : SRMux
    port map (
            O => \N__47358\,
            I => \N__46979\
        );

    \I__11177\ : SRMux
    port map (
            O => \N__47357\,
            I => \N__46979\
        );

    \I__11176\ : SRMux
    port map (
            O => \N__47356\,
            I => \N__46979\
        );

    \I__11175\ : SRMux
    port map (
            O => \N__47355\,
            I => \N__46979\
        );

    \I__11174\ : SRMux
    port map (
            O => \N__47354\,
            I => \N__46979\
        );

    \I__11173\ : SRMux
    port map (
            O => \N__47353\,
            I => \N__46979\
        );

    \I__11172\ : SRMux
    port map (
            O => \N__47352\,
            I => \N__46979\
        );

    \I__11171\ : SRMux
    port map (
            O => \N__47351\,
            I => \N__46979\
        );

    \I__11170\ : SRMux
    port map (
            O => \N__47350\,
            I => \N__46979\
        );

    \I__11169\ : SRMux
    port map (
            O => \N__47349\,
            I => \N__46979\
        );

    \I__11168\ : SRMux
    port map (
            O => \N__47348\,
            I => \N__46979\
        );

    \I__11167\ : SRMux
    port map (
            O => \N__47347\,
            I => \N__46979\
        );

    \I__11166\ : SRMux
    port map (
            O => \N__47346\,
            I => \N__46979\
        );

    \I__11165\ : SRMux
    port map (
            O => \N__47345\,
            I => \N__46979\
        );

    \I__11164\ : SRMux
    port map (
            O => \N__47344\,
            I => \N__46979\
        );

    \I__11163\ : SRMux
    port map (
            O => \N__47343\,
            I => \N__46979\
        );

    \I__11162\ : SRMux
    port map (
            O => \N__47342\,
            I => \N__46979\
        );

    \I__11161\ : SRMux
    port map (
            O => \N__47341\,
            I => \N__46979\
        );

    \I__11160\ : SRMux
    port map (
            O => \N__47340\,
            I => \N__46979\
        );

    \I__11159\ : SRMux
    port map (
            O => \N__47339\,
            I => \N__46979\
        );

    \I__11158\ : SRMux
    port map (
            O => \N__47338\,
            I => \N__46979\
        );

    \I__11157\ : SRMux
    port map (
            O => \N__47337\,
            I => \N__46979\
        );

    \I__11156\ : SRMux
    port map (
            O => \N__47336\,
            I => \N__46979\
        );

    \I__11155\ : SRMux
    port map (
            O => \N__47335\,
            I => \N__46979\
        );

    \I__11154\ : Glb2LocalMux
    port map (
            O => \N__47332\,
            I => \N__46979\
        );

    \I__11153\ : SRMux
    port map (
            O => \N__47331\,
            I => \N__46979\
        );

    \I__11152\ : SRMux
    port map (
            O => \N__47330\,
            I => \N__46979\
        );

    \I__11151\ : SRMux
    port map (
            O => \N__47329\,
            I => \N__46979\
        );

    \I__11150\ : SRMux
    port map (
            O => \N__47328\,
            I => \N__46979\
        );

    \I__11149\ : SRMux
    port map (
            O => \N__47327\,
            I => \N__46979\
        );

    \I__11148\ : SRMux
    port map (
            O => \N__47326\,
            I => \N__46979\
        );

    \I__11147\ : SRMux
    port map (
            O => \N__47325\,
            I => \N__46979\
        );

    \I__11146\ : SRMux
    port map (
            O => \N__47324\,
            I => \N__46979\
        );

    \I__11145\ : SRMux
    port map (
            O => \N__47323\,
            I => \N__46979\
        );

    \I__11144\ : SRMux
    port map (
            O => \N__47322\,
            I => \N__46979\
        );

    \I__11143\ : SRMux
    port map (
            O => \N__47321\,
            I => \N__46979\
        );

    \I__11142\ : SRMux
    port map (
            O => \N__47320\,
            I => \N__46979\
        );

    \I__11141\ : SRMux
    port map (
            O => \N__47319\,
            I => \N__46979\
        );

    \I__11140\ : SRMux
    port map (
            O => \N__47318\,
            I => \N__46979\
        );

    \I__11139\ : SRMux
    port map (
            O => \N__47317\,
            I => \N__46979\
        );

    \I__11138\ : SRMux
    port map (
            O => \N__47316\,
            I => \N__46979\
        );

    \I__11137\ : SRMux
    port map (
            O => \N__47315\,
            I => \N__46979\
        );

    \I__11136\ : SRMux
    port map (
            O => \N__47314\,
            I => \N__46979\
        );

    \I__11135\ : SRMux
    port map (
            O => \N__47313\,
            I => \N__46979\
        );

    \I__11134\ : SRMux
    port map (
            O => \N__47312\,
            I => \N__46979\
        );

    \I__11133\ : SRMux
    port map (
            O => \N__47311\,
            I => \N__46979\
        );

    \I__11132\ : SRMux
    port map (
            O => \N__47310\,
            I => \N__46979\
        );

    \I__11131\ : SRMux
    port map (
            O => \N__47309\,
            I => \N__46979\
        );

    \I__11130\ : SRMux
    port map (
            O => \N__47308\,
            I => \N__46979\
        );

    \I__11129\ : SRMux
    port map (
            O => \N__47307\,
            I => \N__46979\
        );

    \I__11128\ : SRMux
    port map (
            O => \N__47306\,
            I => \N__46979\
        );

    \I__11127\ : SRMux
    port map (
            O => \N__47305\,
            I => \N__46979\
        );

    \I__11126\ : SRMux
    port map (
            O => \N__47304\,
            I => \N__46979\
        );

    \I__11125\ : SRMux
    port map (
            O => \N__47303\,
            I => \N__46979\
        );

    \I__11124\ : SRMux
    port map (
            O => \N__47302\,
            I => \N__46979\
        );

    \I__11123\ : SRMux
    port map (
            O => \N__47301\,
            I => \N__46979\
        );

    \I__11122\ : SRMux
    port map (
            O => \N__47300\,
            I => \N__46979\
        );

    \I__11121\ : SRMux
    port map (
            O => \N__47299\,
            I => \N__46979\
        );

    \I__11120\ : SRMux
    port map (
            O => \N__47298\,
            I => \N__46979\
        );

    \I__11119\ : SRMux
    port map (
            O => \N__47297\,
            I => \N__46979\
        );

    \I__11118\ : SRMux
    port map (
            O => \N__47296\,
            I => \N__46979\
        );

    \I__11117\ : SRMux
    port map (
            O => \N__47295\,
            I => \N__46979\
        );

    \I__11116\ : SRMux
    port map (
            O => \N__47294\,
            I => \N__46979\
        );

    \I__11115\ : SRMux
    port map (
            O => \N__47293\,
            I => \N__46979\
        );

    \I__11114\ : SRMux
    port map (
            O => \N__47292\,
            I => \N__46979\
        );

    \I__11113\ : SRMux
    port map (
            O => \N__47291\,
            I => \N__46979\
        );

    \I__11112\ : SRMux
    port map (
            O => \N__47290\,
            I => \N__46979\
        );

    \I__11111\ : SRMux
    port map (
            O => \N__47289\,
            I => \N__46979\
        );

    \I__11110\ : SRMux
    port map (
            O => \N__47288\,
            I => \N__46979\
        );

    \I__11109\ : SRMux
    port map (
            O => \N__47287\,
            I => \N__46979\
        );

    \I__11108\ : SRMux
    port map (
            O => \N__47286\,
            I => \N__46979\
        );

    \I__11107\ : Glb2LocalMux
    port map (
            O => \N__47283\,
            I => \N__46979\
        );

    \I__11106\ : Glb2LocalMux
    port map (
            O => \N__47280\,
            I => \N__46979\
        );

    \I__11105\ : SRMux
    port map (
            O => \N__47279\,
            I => \N__46979\
        );

    \I__11104\ : SRMux
    port map (
            O => \N__47278\,
            I => \N__46979\
        );

    \I__11103\ : SRMux
    port map (
            O => \N__47277\,
            I => \N__46979\
        );

    \I__11102\ : SRMux
    port map (
            O => \N__47276\,
            I => \N__46979\
        );

    \I__11101\ : SRMux
    port map (
            O => \N__47275\,
            I => \N__46979\
        );

    \I__11100\ : SRMux
    port map (
            O => \N__47274\,
            I => \N__46979\
        );

    \I__11099\ : SRMux
    port map (
            O => \N__47273\,
            I => \N__46979\
        );

    \I__11098\ : SRMux
    port map (
            O => \N__47272\,
            I => \N__46979\
        );

    \I__11097\ : GlobalMux
    port map (
            O => \N__46979\,
            I => \N__46976\
        );

    \I__11096\ : gio2CtrlBuf
    port map (
            O => \N__46976\,
            I => red_c_g
        );

    \I__11095\ : CascadeMux
    port map (
            O => \N__46973\,
            I => \N__46970\
        );

    \I__11094\ : InMux
    port map (
            O => \N__46970\,
            I => \N__46966\
        );

    \I__11093\ : InMux
    port map (
            O => \N__46969\,
            I => \N__46963\
        );

    \I__11092\ : LocalMux
    port map (
            O => \N__46966\,
            I => \N__46960\
        );

    \I__11091\ : LocalMux
    port map (
            O => \N__46963\,
            I => \N__46957\
        );

    \I__11090\ : Span4Mux_h
    port map (
            O => \N__46960\,
            I => \N__46954\
        );

    \I__11089\ : Span4Mux_h
    port map (
            O => \N__46957\,
            I => \N__46951\
        );

    \I__11088\ : Odrv4
    port map (
            O => \N__46954\,
            I => \delay_measurement_inst.elapsed_time_tr_5\
        );

    \I__11087\ : Odrv4
    port map (
            O => \N__46951\,
            I => \delay_measurement_inst.elapsed_time_tr_5\
        );

    \I__11086\ : InMux
    port map (
            O => \N__46946\,
            I => \N__46942\
        );

    \I__11085\ : InMux
    port map (
            O => \N__46945\,
            I => \N__46938\
        );

    \I__11084\ : LocalMux
    port map (
            O => \N__46942\,
            I => \N__46935\
        );

    \I__11083\ : InMux
    port map (
            O => \N__46941\,
            I => \N__46932\
        );

    \I__11082\ : LocalMux
    port map (
            O => \N__46938\,
            I => \N__46929\
        );

    \I__11081\ : Span4Mux_v
    port map (
            O => \N__46935\,
            I => \N__46924\
        );

    \I__11080\ : LocalMux
    port map (
            O => \N__46932\,
            I => \N__46924\
        );

    \I__11079\ : Span4Mux_h
    port map (
            O => \N__46929\,
            I => \N__46919\
        );

    \I__11078\ : Span4Mux_h
    port map (
            O => \N__46924\,
            I => \N__46919\
        );

    \I__11077\ : Odrv4
    port map (
            O => \N__46919\,
            I => measured_delay_tr_5
        );

    \I__11076\ : InMux
    port map (
            O => \N__46916\,
            I => \N__46911\
        );

    \I__11075\ : InMux
    port map (
            O => \N__46915\,
            I => \N__46906\
        );

    \I__11074\ : InMux
    port map (
            O => \N__46914\,
            I => \N__46906\
        );

    \I__11073\ : LocalMux
    port map (
            O => \N__46911\,
            I => \N__46903\
        );

    \I__11072\ : LocalMux
    port map (
            O => \N__46906\,
            I => \N__46900\
        );

    \I__11071\ : Span4Mux_v
    port map (
            O => \N__46903\,
            I => \N__46897\
        );

    \I__11070\ : Span4Mux_h
    port map (
            O => \N__46900\,
            I => \N__46894\
        );

    \I__11069\ : Odrv4
    port map (
            O => \N__46897\,
            I => \delay_measurement_inst.elapsed_time_tr_3\
        );

    \I__11068\ : Odrv4
    port map (
            O => \N__46894\,
            I => \delay_measurement_inst.elapsed_time_tr_3\
        );

    \I__11067\ : CascadeMux
    port map (
            O => \N__46889\,
            I => \N__46885\
        );

    \I__11066\ : CascadeMux
    port map (
            O => \N__46888\,
            I => \N__46881\
        );

    \I__11065\ : InMux
    port map (
            O => \N__46885\,
            I => \N__46878\
        );

    \I__11064\ : InMux
    port map (
            O => \N__46884\,
            I => \N__46875\
        );

    \I__11063\ : InMux
    port map (
            O => \N__46881\,
            I => \N__46872\
        );

    \I__11062\ : LocalMux
    port map (
            O => \N__46878\,
            I => \N__46867\
        );

    \I__11061\ : LocalMux
    port map (
            O => \N__46875\,
            I => \N__46867\
        );

    \I__11060\ : LocalMux
    port map (
            O => \N__46872\,
            I => \N__46864\
        );

    \I__11059\ : Span4Mux_h
    port map (
            O => \N__46867\,
            I => \N__46861\
        );

    \I__11058\ : Span4Mux_h
    port map (
            O => \N__46864\,
            I => \N__46858\
        );

    \I__11057\ : Span4Mux_v
    port map (
            O => \N__46861\,
            I => \N__46855\
        );

    \I__11056\ : Odrv4
    port map (
            O => \N__46858\,
            I => measured_delay_tr_3
        );

    \I__11055\ : Odrv4
    port map (
            O => \N__46855\,
            I => measured_delay_tr_3
        );

    \I__11054\ : CascadeMux
    port map (
            O => \N__46850\,
            I => \N__46846\
        );

    \I__11053\ : InMux
    port map (
            O => \N__46849\,
            I => \N__46843\
        );

    \I__11052\ : InMux
    port map (
            O => \N__46846\,
            I => \N__46840\
        );

    \I__11051\ : LocalMux
    port map (
            O => \N__46843\,
            I => \N__46837\
        );

    \I__11050\ : LocalMux
    port map (
            O => \N__46840\,
            I => \N__46834\
        );

    \I__11049\ : Span4Mux_h
    port map (
            O => \N__46837\,
            I => \N__46831\
        );

    \I__11048\ : Span4Mux_h
    port map (
            O => \N__46834\,
            I => \N__46828\
        );

    \I__11047\ : Odrv4
    port map (
            O => \N__46831\,
            I => \delay_measurement_inst.elapsed_time_tr_8\
        );

    \I__11046\ : Odrv4
    port map (
            O => \N__46828\,
            I => \delay_measurement_inst.elapsed_time_tr_8\
        );

    \I__11045\ : InMux
    port map (
            O => \N__46823\,
            I => \N__46819\
        );

    \I__11044\ : InMux
    port map (
            O => \N__46822\,
            I => \N__46816\
        );

    \I__11043\ : LocalMux
    port map (
            O => \N__46819\,
            I => \N__46812\
        );

    \I__11042\ : LocalMux
    port map (
            O => \N__46816\,
            I => \N__46809\
        );

    \I__11041\ : InMux
    port map (
            O => \N__46815\,
            I => \N__46806\
        );

    \I__11040\ : Span4Mux_v
    port map (
            O => \N__46812\,
            I => \N__46803\
        );

    \I__11039\ : Span4Mux_v
    port map (
            O => \N__46809\,
            I => \N__46798\
        );

    \I__11038\ : LocalMux
    port map (
            O => \N__46806\,
            I => \N__46798\
        );

    \I__11037\ : Span4Mux_h
    port map (
            O => \N__46803\,
            I => \N__46795\
        );

    \I__11036\ : Span4Mux_h
    port map (
            O => \N__46798\,
            I => \N__46792\
        );

    \I__11035\ : Odrv4
    port map (
            O => \N__46795\,
            I => measured_delay_tr_8
        );

    \I__11034\ : Odrv4
    port map (
            O => \N__46792\,
            I => measured_delay_tr_8
        );

    \I__11033\ : InMux
    port map (
            O => \N__46787\,
            I => \N__46783\
        );

    \I__11032\ : InMux
    port map (
            O => \N__46786\,
            I => \N__46780\
        );

    \I__11031\ : LocalMux
    port map (
            O => \N__46783\,
            I => \N__46777\
        );

    \I__11030\ : LocalMux
    port map (
            O => \N__46780\,
            I => \N__46774\
        );

    \I__11029\ : Span4Mux_v
    port map (
            O => \N__46777\,
            I => \N__46771\
        );

    \I__11028\ : Span4Mux_h
    port map (
            O => \N__46774\,
            I => \N__46768\
        );

    \I__11027\ : Odrv4
    port map (
            O => \N__46771\,
            I => \delay_measurement_inst.elapsed_time_tr_7\
        );

    \I__11026\ : Odrv4
    port map (
            O => \N__46768\,
            I => \delay_measurement_inst.elapsed_time_tr_7\
        );

    \I__11025\ : InMux
    port map (
            O => \N__46763\,
            I => \N__46760\
        );

    \I__11024\ : LocalMux
    port map (
            O => \N__46760\,
            I => \N__46755\
        );

    \I__11023\ : InMux
    port map (
            O => \N__46759\,
            I => \N__46752\
        );

    \I__11022\ : InMux
    port map (
            O => \N__46758\,
            I => \N__46749\
        );

    \I__11021\ : Span4Mux_v
    port map (
            O => \N__46755\,
            I => \N__46742\
        );

    \I__11020\ : LocalMux
    port map (
            O => \N__46752\,
            I => \N__46742\
        );

    \I__11019\ : LocalMux
    port map (
            O => \N__46749\,
            I => \N__46742\
        );

    \I__11018\ : Span4Mux_h
    port map (
            O => \N__46742\,
            I => \N__46739\
        );

    \I__11017\ : Odrv4
    port map (
            O => \N__46739\,
            I => measured_delay_tr_7
        );

    \I__11016\ : InMux
    port map (
            O => \N__46736\,
            I => \N__46731\
        );

    \I__11015\ : InMux
    port map (
            O => \N__46735\,
            I => \N__46728\
        );

    \I__11014\ : CascadeMux
    port map (
            O => \N__46734\,
            I => \N__46725\
        );

    \I__11013\ : LocalMux
    port map (
            O => \N__46731\,
            I => \N__46722\
        );

    \I__11012\ : LocalMux
    port map (
            O => \N__46728\,
            I => \N__46719\
        );

    \I__11011\ : InMux
    port map (
            O => \N__46725\,
            I => \N__46716\
        );

    \I__11010\ : Span4Mux_h
    port map (
            O => \N__46722\,
            I => \N__46713\
        );

    \I__11009\ : Span4Mux_h
    port map (
            O => \N__46719\,
            I => \N__46710\
        );

    \I__11008\ : LocalMux
    port map (
            O => \N__46716\,
            I => \N__46707\
        );

    \I__11007\ : Odrv4
    port map (
            O => \N__46713\,
            I => \delay_measurement_inst.elapsed_time_tr_17\
        );

    \I__11006\ : Odrv4
    port map (
            O => \N__46710\,
            I => \delay_measurement_inst.elapsed_time_tr_17\
        );

    \I__11005\ : Odrv12
    port map (
            O => \N__46707\,
            I => \delay_measurement_inst.elapsed_time_tr_17\
        );

    \I__11004\ : InMux
    port map (
            O => \N__46700\,
            I => \N__46696\
        );

    \I__11003\ : CascadeMux
    port map (
            O => \N__46699\,
            I => \N__46693\
        );

    \I__11002\ : LocalMux
    port map (
            O => \N__46696\,
            I => \N__46690\
        );

    \I__11001\ : InMux
    port map (
            O => \N__46693\,
            I => \N__46687\
        );

    \I__11000\ : Span4Mux_v
    port map (
            O => \N__46690\,
            I => \N__46682\
        );

    \I__10999\ : LocalMux
    port map (
            O => \N__46687\,
            I => \N__46682\
        );

    \I__10998\ : Odrv4
    port map (
            O => \N__46682\,
            I => \delay_measurement_inst.elapsed_time_tr_13\
        );

    \I__10997\ : InMux
    port map (
            O => \N__46679\,
            I => \N__46675\
        );

    \I__10996\ : CascadeMux
    port map (
            O => \N__46678\,
            I => \N__46671\
        );

    \I__10995\ : LocalMux
    port map (
            O => \N__46675\,
            I => \N__46668\
        );

    \I__10994\ : InMux
    port map (
            O => \N__46674\,
            I => \N__46665\
        );

    \I__10993\ : InMux
    port map (
            O => \N__46671\,
            I => \N__46662\
        );

    \I__10992\ : Span4Mux_v
    port map (
            O => \N__46668\,
            I => \N__46655\
        );

    \I__10991\ : LocalMux
    port map (
            O => \N__46665\,
            I => \N__46655\
        );

    \I__10990\ : LocalMux
    port map (
            O => \N__46662\,
            I => \N__46655\
        );

    \I__10989\ : Span4Mux_v
    port map (
            O => \N__46655\,
            I => \N__46652\
        );

    \I__10988\ : Odrv4
    port map (
            O => \N__46652\,
            I => measured_delay_tr_13
        );

    \I__10987\ : InMux
    port map (
            O => \N__46649\,
            I => \N__46644\
        );

    \I__10986\ : InMux
    port map (
            O => \N__46648\,
            I => \N__46641\
        );

    \I__10985\ : InMux
    port map (
            O => \N__46647\,
            I => \N__46638\
        );

    \I__10984\ : LocalMux
    port map (
            O => \N__46644\,
            I => \N__46630\
        );

    \I__10983\ : LocalMux
    port map (
            O => \N__46641\,
            I => \N__46630\
        );

    \I__10982\ : LocalMux
    port map (
            O => \N__46638\,
            I => \N__46630\
        );

    \I__10981\ : InMux
    port map (
            O => \N__46637\,
            I => \N__46627\
        );

    \I__10980\ : Span4Mux_v
    port map (
            O => \N__46630\,
            I => \N__46622\
        );

    \I__10979\ : LocalMux
    port map (
            O => \N__46627\,
            I => \N__46622\
        );

    \I__10978\ : Odrv4
    port map (
            O => \N__46622\,
            I => \delay_measurement_inst.delay_tr_reg3lto6\
        );

    \I__10977\ : InMux
    port map (
            O => \N__46619\,
            I => \N__46616\
        );

    \I__10976\ : LocalMux
    port map (
            O => \N__46616\,
            I => \N__46611\
        );

    \I__10975\ : InMux
    port map (
            O => \N__46615\,
            I => \N__46608\
        );

    \I__10974\ : InMux
    port map (
            O => \N__46614\,
            I => \N__46605\
        );

    \I__10973\ : Span4Mux_v
    port map (
            O => \N__46611\,
            I => \N__46598\
        );

    \I__10972\ : LocalMux
    port map (
            O => \N__46608\,
            I => \N__46598\
        );

    \I__10971\ : LocalMux
    port map (
            O => \N__46605\,
            I => \N__46598\
        );

    \I__10970\ : Span4Mux_h
    port map (
            O => \N__46598\,
            I => \N__46595\
        );

    \I__10969\ : Odrv4
    port map (
            O => \N__46595\,
            I => measured_delay_tr_6
        );

    \I__10968\ : InMux
    port map (
            O => \N__46592\,
            I => \N__46588\
        );

    \I__10967\ : InMux
    port map (
            O => \N__46591\,
            I => \N__46585\
        );

    \I__10966\ : LocalMux
    port map (
            O => \N__46588\,
            I => \N__46582\
        );

    \I__10965\ : LocalMux
    port map (
            O => \N__46585\,
            I => \N__46579\
        );

    \I__10964\ : Span4Mux_v
    port map (
            O => \N__46582\,
            I => \N__46576\
        );

    \I__10963\ : Span4Mux_h
    port map (
            O => \N__46579\,
            I => \N__46573\
        );

    \I__10962\ : Odrv4
    port map (
            O => \N__46576\,
            I => \delay_measurement_inst.elapsed_time_tr_4\
        );

    \I__10961\ : Odrv4
    port map (
            O => \N__46573\,
            I => \delay_measurement_inst.elapsed_time_tr_4\
        );

    \I__10960\ : InMux
    port map (
            O => \N__46568\,
            I => \N__46565\
        );

    \I__10959\ : LocalMux
    port map (
            O => \N__46565\,
            I => \N__46560\
        );

    \I__10958\ : InMux
    port map (
            O => \N__46564\,
            I => \N__46557\
        );

    \I__10957\ : InMux
    port map (
            O => \N__46563\,
            I => \N__46554\
        );

    \I__10956\ : Span4Mux_v
    port map (
            O => \N__46560\,
            I => \N__46547\
        );

    \I__10955\ : LocalMux
    port map (
            O => \N__46557\,
            I => \N__46547\
        );

    \I__10954\ : LocalMux
    port map (
            O => \N__46554\,
            I => \N__46547\
        );

    \I__10953\ : Span4Mux_h
    port map (
            O => \N__46547\,
            I => \N__46544\
        );

    \I__10952\ : Odrv4
    port map (
            O => \N__46544\,
            I => measured_delay_tr_4
        );

    \I__10951\ : InMux
    port map (
            O => \N__46541\,
            I => \N__46525\
        );

    \I__10950\ : InMux
    port map (
            O => \N__46540\,
            I => \N__46525\
        );

    \I__10949\ : InMux
    port map (
            O => \N__46539\,
            I => \N__46525\
        );

    \I__10948\ : InMux
    port map (
            O => \N__46538\,
            I => \N__46525\
        );

    \I__10947\ : InMux
    port map (
            O => \N__46537\,
            I => \N__46516\
        );

    \I__10946\ : InMux
    port map (
            O => \N__46536\,
            I => \N__46516\
        );

    \I__10945\ : InMux
    port map (
            O => \N__46535\,
            I => \N__46516\
        );

    \I__10944\ : InMux
    port map (
            O => \N__46534\,
            I => \N__46516\
        );

    \I__10943\ : LocalMux
    port map (
            O => \N__46525\,
            I => \N__46513\
        );

    \I__10942\ : LocalMux
    port map (
            O => \N__46516\,
            I => \N__46510\
        );

    \I__10941\ : Span4Mux_h
    port map (
            O => \N__46513\,
            I => \N__46507\
        );

    \I__10940\ : Span4Mux_h
    port map (
            O => \N__46510\,
            I => \N__46504\
        );

    \I__10939\ : Odrv4
    port map (
            O => \N__46507\,
            I => \delay_measurement_inst.N_324\
        );

    \I__10938\ : Odrv4
    port map (
            O => \N__46504\,
            I => \delay_measurement_inst.N_324\
        );

    \I__10937\ : InMux
    port map (
            O => \N__46499\,
            I => \N__46490\
        );

    \I__10936\ : InMux
    port map (
            O => \N__46498\,
            I => \N__46490\
        );

    \I__10935\ : InMux
    port map (
            O => \N__46497\,
            I => \N__46490\
        );

    \I__10934\ : LocalMux
    port map (
            O => \N__46490\,
            I => \N__46484\
        );

    \I__10933\ : InMux
    port map (
            O => \N__46489\,
            I => \N__46477\
        );

    \I__10932\ : InMux
    port map (
            O => \N__46488\,
            I => \N__46477\
        );

    \I__10931\ : InMux
    port map (
            O => \N__46487\,
            I => \N__46477\
        );

    \I__10930\ : Odrv4
    port map (
            O => \N__46484\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNI80KG7_6\
        );

    \I__10929\ : LocalMux
    port map (
            O => \N__46477\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNI80KG7_6\
        );

    \I__10928\ : InMux
    port map (
            O => \N__46472\,
            I => \N__46469\
        );

    \I__10927\ : LocalMux
    port map (
            O => \N__46469\,
            I => \N__46464\
        );

    \I__10926\ : CascadeMux
    port map (
            O => \N__46468\,
            I => \N__46461\
        );

    \I__10925\ : InMux
    port map (
            O => \N__46467\,
            I => \N__46458\
        );

    \I__10924\ : Span4Mux_h
    port map (
            O => \N__46464\,
            I => \N__46455\
        );

    \I__10923\ : InMux
    port map (
            O => \N__46461\,
            I => \N__46452\
        );

    \I__10922\ : LocalMux
    port map (
            O => \N__46458\,
            I => \N__46449\
        );

    \I__10921\ : Span4Mux_v
    port map (
            O => \N__46455\,
            I => \N__46444\
        );

    \I__10920\ : LocalMux
    port map (
            O => \N__46452\,
            I => \N__46444\
        );

    \I__10919\ : Span4Mux_h
    port map (
            O => \N__46449\,
            I => \N__46441\
        );

    \I__10918\ : Span4Mux_h
    port map (
            O => \N__46444\,
            I => \N__46438\
        );

    \I__10917\ : Odrv4
    port map (
            O => \N__46441\,
            I => \delay_measurement_inst.elapsed_time_tr_2\
        );

    \I__10916\ : Odrv4
    port map (
            O => \N__46438\,
            I => \delay_measurement_inst.elapsed_time_tr_2\
        );

    \I__10915\ : CascadeMux
    port map (
            O => \N__46433\,
            I => \N__46429\
        );

    \I__10914\ : CascadeMux
    port map (
            O => \N__46432\,
            I => \N__46426\
        );

    \I__10913\ : InMux
    port map (
            O => \N__46429\,
            I => \N__46423\
        );

    \I__10912\ : InMux
    port map (
            O => \N__46426\,
            I => \N__46419\
        );

    \I__10911\ : LocalMux
    port map (
            O => \N__46423\,
            I => \N__46416\
        );

    \I__10910\ : InMux
    port map (
            O => \N__46422\,
            I => \N__46413\
        );

    \I__10909\ : LocalMux
    port map (
            O => \N__46419\,
            I => \N__46410\
        );

    \I__10908\ : Span4Mux_h
    port map (
            O => \N__46416\,
            I => \N__46405\
        );

    \I__10907\ : LocalMux
    port map (
            O => \N__46413\,
            I => \N__46405\
        );

    \I__10906\ : Span4Mux_h
    port map (
            O => \N__46410\,
            I => \N__46402\
        );

    \I__10905\ : Span4Mux_v
    port map (
            O => \N__46405\,
            I => \N__46399\
        );

    \I__10904\ : Odrv4
    port map (
            O => \N__46402\,
            I => measured_delay_tr_2
        );

    \I__10903\ : Odrv4
    port map (
            O => \N__46399\,
            I => measured_delay_tr_2
        );

    \I__10902\ : CascadeMux
    port map (
            O => \N__46394\,
            I => \delay_measurement_inst.delay_tr_timer.N_331_cascade_\
        );

    \I__10901\ : InMux
    port map (
            O => \N__46391\,
            I => \N__46388\
        );

    \I__10900\ : LocalMux
    port map (
            O => \N__46388\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_5\
        );

    \I__10899\ : InMux
    port map (
            O => \N__46385\,
            I => \N__46382\
        );

    \I__10898\ : LocalMux
    port map (
            O => \N__46382\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_7\
        );

    \I__10897\ : CascadeMux
    port map (
            O => \N__46379\,
            I => \delay_measurement_inst.delay_tr_timer.N_321_cascade_\
        );

    \I__10896\ : InMux
    port map (
            O => \N__46376\,
            I => \N__46372\
        );

    \I__10895\ : InMux
    port map (
            O => \N__46375\,
            I => \N__46369\
        );

    \I__10894\ : LocalMux
    port map (
            O => \N__46372\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILUISZ0Z_14\
        );

    \I__10893\ : LocalMux
    port map (
            O => \N__46369\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILUISZ0Z_14\
        );

    \I__10892\ : InMux
    port map (
            O => \N__46364\,
            I => \N__46358\
        );

    \I__10891\ : InMux
    port map (
            O => \N__46363\,
            I => \N__46358\
        );

    \I__10890\ : LocalMux
    port map (
            O => \N__46358\,
            I => \delay_measurement_inst.delay_tr_timer.N_331\
        );

    \I__10889\ : InMux
    port map (
            O => \N__46355\,
            I => \N__46352\
        );

    \I__10888\ : LocalMux
    port map (
            O => \N__46352\,
            I => \delay_measurement_inst.delay_tr_reg_esr_RNO_0Z0Z_14\
        );

    \I__10887\ : InMux
    port map (
            O => \N__46349\,
            I => \N__46345\
        );

    \I__10886\ : InMux
    port map (
            O => \N__46348\,
            I => \N__46342\
        );

    \I__10885\ : LocalMux
    port map (
            O => \N__46345\,
            I => \N__46337\
        );

    \I__10884\ : LocalMux
    port map (
            O => \N__46342\,
            I => \N__46334\
        );

    \I__10883\ : InMux
    port map (
            O => \N__46341\,
            I => \N__46329\
        );

    \I__10882\ : InMux
    port map (
            O => \N__46340\,
            I => \N__46329\
        );

    \I__10881\ : Span4Mux_v
    port map (
            O => \N__46337\,
            I => \N__46322\
        );

    \I__10880\ : Span4Mux_v
    port map (
            O => \N__46334\,
            I => \N__46322\
        );

    \I__10879\ : LocalMux
    port map (
            O => \N__46329\,
            I => \N__46322\
        );

    \I__10878\ : Odrv4
    port map (
            O => \N__46322\,
            I => \delay_measurement_inst.delay_tr_reg3lto14\
        );

    \I__10877\ : InMux
    port map (
            O => \N__46319\,
            I => \N__46314\
        );

    \I__10876\ : InMux
    port map (
            O => \N__46318\,
            I => \N__46309\
        );

    \I__10875\ : InMux
    port map (
            O => \N__46317\,
            I => \N__46306\
        );

    \I__10874\ : LocalMux
    port map (
            O => \N__46314\,
            I => \N__46303\
        );

    \I__10873\ : InMux
    port map (
            O => \N__46313\,
            I => \N__46298\
        );

    \I__10872\ : InMux
    port map (
            O => \N__46312\,
            I => \N__46298\
        );

    \I__10871\ : LocalMux
    port map (
            O => \N__46309\,
            I => \N__46295\
        );

    \I__10870\ : LocalMux
    port map (
            O => \N__46306\,
            I => \N__46288\
        );

    \I__10869\ : Span4Mux_v
    port map (
            O => \N__46303\,
            I => \N__46288\
        );

    \I__10868\ : LocalMux
    port map (
            O => \N__46298\,
            I => \N__46288\
        );

    \I__10867\ : Span12Mux_v
    port map (
            O => \N__46295\,
            I => \N__46285\
        );

    \I__10866\ : Span4Mux_v
    port map (
            O => \N__46288\,
            I => \N__46282\
        );

    \I__10865\ : Odrv12
    port map (
            O => \N__46285\,
            I => measured_delay_tr_14
        );

    \I__10864\ : Odrv4
    port map (
            O => \N__46282\,
            I => measured_delay_tr_14
        );

    \I__10863\ : InMux
    port map (
            O => \N__46277\,
            I => \N__46269\
        );

    \I__10862\ : CascadeMux
    port map (
            O => \N__46276\,
            I => \N__46266\
        );

    \I__10861\ : InMux
    port map (
            O => \N__46275\,
            I => \N__46263\
        );

    \I__10860\ : InMux
    port map (
            O => \N__46274\,
            I => \N__46260\
        );

    \I__10859\ : InMux
    port map (
            O => \N__46273\,
            I => \N__46255\
        );

    \I__10858\ : InMux
    port map (
            O => \N__46272\,
            I => \N__46255\
        );

    \I__10857\ : LocalMux
    port map (
            O => \N__46269\,
            I => \N__46251\
        );

    \I__10856\ : InMux
    port map (
            O => \N__46266\,
            I => \N__46248\
        );

    \I__10855\ : LocalMux
    port map (
            O => \N__46263\,
            I => \N__46241\
        );

    \I__10854\ : LocalMux
    port map (
            O => \N__46260\,
            I => \N__46241\
        );

    \I__10853\ : LocalMux
    port map (
            O => \N__46255\,
            I => \N__46241\
        );

    \I__10852\ : InMux
    port map (
            O => \N__46254\,
            I => \N__46238\
        );

    \I__10851\ : Span4Mux_v
    port map (
            O => \N__46251\,
            I => \N__46235\
        );

    \I__10850\ : LocalMux
    port map (
            O => \N__46248\,
            I => \N__46232\
        );

    \I__10849\ : Span4Mux_v
    port map (
            O => \N__46241\,
            I => \N__46229\
        );

    \I__10848\ : LocalMux
    port map (
            O => \N__46238\,
            I => \N__46226\
        );

    \I__10847\ : Odrv4
    port map (
            O => \N__46235\,
            I => \delay_measurement_inst.delay_tr_reg3lto15\
        );

    \I__10846\ : Odrv4
    port map (
            O => \N__46232\,
            I => \delay_measurement_inst.delay_tr_reg3lto15\
        );

    \I__10845\ : Odrv4
    port map (
            O => \N__46229\,
            I => \delay_measurement_inst.delay_tr_reg3lto15\
        );

    \I__10844\ : Odrv12
    port map (
            O => \N__46226\,
            I => \delay_measurement_inst.delay_tr_reg3lto15\
        );

    \I__10843\ : CascadeMux
    port map (
            O => \N__46217\,
            I => \N__46214\
        );

    \I__10842\ : InMux
    port map (
            O => \N__46214\,
            I => \N__46210\
        );

    \I__10841\ : InMux
    port map (
            O => \N__46213\,
            I => \N__46207\
        );

    \I__10840\ : LocalMux
    port map (
            O => \N__46210\,
            I => \N__46201\
        );

    \I__10839\ : LocalMux
    port map (
            O => \N__46207\,
            I => \N__46198\
        );

    \I__10838\ : InMux
    port map (
            O => \N__46206\,
            I => \N__46191\
        );

    \I__10837\ : InMux
    port map (
            O => \N__46205\,
            I => \N__46191\
        );

    \I__10836\ : InMux
    port map (
            O => \N__46204\,
            I => \N__46191\
        );

    \I__10835\ : Odrv4
    port map (
            O => \N__46201\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNIM96P1_16\
        );

    \I__10834\ : Odrv12
    port map (
            O => \N__46198\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNIM96P1_16\
        );

    \I__10833\ : LocalMux
    port map (
            O => \N__46191\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNIM96P1_16\
        );

    \I__10832\ : CascadeMux
    port map (
            O => \N__46184\,
            I => \N__46174\
        );

    \I__10831\ : InMux
    port map (
            O => \N__46183\,
            I => \N__46170\
        );

    \I__10830\ : InMux
    port map (
            O => \N__46182\,
            I => \N__46167\
        );

    \I__10829\ : InMux
    port map (
            O => \N__46181\,
            I => \N__46164\
        );

    \I__10828\ : InMux
    port map (
            O => \N__46180\,
            I => \N__46161\
        );

    \I__10827\ : InMux
    port map (
            O => \N__46179\,
            I => \N__46156\
        );

    \I__10826\ : InMux
    port map (
            O => \N__46178\,
            I => \N__46156\
        );

    \I__10825\ : CascadeMux
    port map (
            O => \N__46177\,
            I => \N__46152\
        );

    \I__10824\ : InMux
    port map (
            O => \N__46174\,
            I => \N__46149\
        );

    \I__10823\ : InMux
    port map (
            O => \N__46173\,
            I => \N__46146\
        );

    \I__10822\ : LocalMux
    port map (
            O => \N__46170\,
            I => \N__46143\
        );

    \I__10821\ : LocalMux
    port map (
            O => \N__46167\,
            I => \N__46140\
        );

    \I__10820\ : LocalMux
    port map (
            O => \N__46164\,
            I => \N__46137\
        );

    \I__10819\ : LocalMux
    port map (
            O => \N__46161\,
            I => \N__46132\
        );

    \I__10818\ : LocalMux
    port map (
            O => \N__46156\,
            I => \N__46132\
        );

    \I__10817\ : InMux
    port map (
            O => \N__46155\,
            I => \N__46127\
        );

    \I__10816\ : InMux
    port map (
            O => \N__46152\,
            I => \N__46127\
        );

    \I__10815\ : LocalMux
    port map (
            O => \N__46149\,
            I => \N__46120\
        );

    \I__10814\ : LocalMux
    port map (
            O => \N__46146\,
            I => \N__46120\
        );

    \I__10813\ : Span4Mux_v
    port map (
            O => \N__46143\,
            I => \N__46120\
        );

    \I__10812\ : Span4Mux_v
    port map (
            O => \N__46140\,
            I => \N__46115\
        );

    \I__10811\ : Span4Mux_v
    port map (
            O => \N__46137\,
            I => \N__46115\
        );

    \I__10810\ : Span4Mux_v
    port map (
            O => \N__46132\,
            I => \N__46110\
        );

    \I__10809\ : LocalMux
    port map (
            O => \N__46127\,
            I => \N__46110\
        );

    \I__10808\ : Span4Mux_h
    port map (
            O => \N__46120\,
            I => \N__46105\
        );

    \I__10807\ : Span4Mux_h
    port map (
            O => \N__46115\,
            I => \N__46105\
        );

    \I__10806\ : Span4Mux_v
    port map (
            O => \N__46110\,
            I => \N__46102\
        );

    \I__10805\ : Span4Mux_v
    port map (
            O => \N__46105\,
            I => \N__46099\
        );

    \I__10804\ : Span4Mux_h
    port map (
            O => \N__46102\,
            I => \N__46096\
        );

    \I__10803\ : Odrv4
    port map (
            O => \N__46099\,
            I => measured_delay_tr_15
        );

    \I__10802\ : Odrv4
    port map (
            O => \N__46096\,
            I => measured_delay_tr_15
        );

    \I__10801\ : InMux
    port map (
            O => \N__46091\,
            I => \N__46087\
        );

    \I__10800\ : InMux
    port map (
            O => \N__46090\,
            I => \N__46084\
        );

    \I__10799\ : LocalMux
    port map (
            O => \N__46087\,
            I => \N__46081\
        );

    \I__10798\ : LocalMux
    port map (
            O => \N__46084\,
            I => \N__46078\
        );

    \I__10797\ : Span4Mux_v
    port map (
            O => \N__46081\,
            I => \N__46075\
        );

    \I__10796\ : Span4Mux_h
    port map (
            O => \N__46078\,
            I => \N__46072\
        );

    \I__10795\ : Odrv4
    port map (
            O => \N__46075\,
            I => \delay_measurement_inst.elapsed_time_tr_1\
        );

    \I__10794\ : Odrv4
    port map (
            O => \N__46072\,
            I => \delay_measurement_inst.elapsed_time_tr_1\
        );

    \I__10793\ : CascadeMux
    port map (
            O => \N__46067\,
            I => \N__46064\
        );

    \I__10792\ : InMux
    port map (
            O => \N__46064\,
            I => \N__46061\
        );

    \I__10791\ : LocalMux
    port map (
            O => \N__46061\,
            I => \N__46057\
        );

    \I__10790\ : CascadeMux
    port map (
            O => \N__46060\,
            I => \N__46054\
        );

    \I__10789\ : Span4Mux_v
    port map (
            O => \N__46057\,
            I => \N__46051\
        );

    \I__10788\ : InMux
    port map (
            O => \N__46054\,
            I => \N__46048\
        );

    \I__10787\ : Span4Mux_h
    port map (
            O => \N__46051\,
            I => \N__46043\
        );

    \I__10786\ : LocalMux
    port map (
            O => \N__46048\,
            I => \N__46043\
        );

    \I__10785\ : Span4Mux_h
    port map (
            O => \N__46043\,
            I => \N__46040\
        );

    \I__10784\ : Odrv4
    port map (
            O => \N__46040\,
            I => measured_delay_tr_1
        );

    \I__10783\ : CascadeMux
    port map (
            O => \N__46037\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3_cascade_\
        );

    \I__10782\ : InMux
    port map (
            O => \N__46034\,
            I => \N__46031\
        );

    \I__10781\ : LocalMux
    port map (
            O => \N__46031\,
            I => \N__46025\
        );

    \I__10780\ : InMux
    port map (
            O => \N__46030\,
            I => \N__46022\
        );

    \I__10779\ : InMux
    port map (
            O => \N__46029\,
            I => \N__46018\
        );

    \I__10778\ : InMux
    port map (
            O => \N__46028\,
            I => \N__46015\
        );

    \I__10777\ : Span4Mux_v
    port map (
            O => \N__46025\,
            I => \N__46012\
        );

    \I__10776\ : LocalMux
    port map (
            O => \N__46022\,
            I => \N__46009\
        );

    \I__10775\ : InMux
    port map (
            O => \N__46021\,
            I => \N__46006\
        );

    \I__10774\ : LocalMux
    port map (
            O => \N__46018\,
            I => \N__46003\
        );

    \I__10773\ : LocalMux
    port map (
            O => \N__46015\,
            I => \N__46000\
        );

    \I__10772\ : Span4Mux_v
    port map (
            O => \N__46012\,
            I => \N__45993\
        );

    \I__10771\ : Span4Mux_v
    port map (
            O => \N__46009\,
            I => \N__45993\
        );

    \I__10770\ : LocalMux
    port map (
            O => \N__46006\,
            I => \N__45993\
        );

    \I__10769\ : Odrv4
    port map (
            O => \N__46003\,
            I => \delay_measurement_inst.delay_tr_reg3lto9\
        );

    \I__10768\ : Odrv4
    port map (
            O => \N__46000\,
            I => \delay_measurement_inst.delay_tr_reg3lto9\
        );

    \I__10767\ : Odrv4
    port map (
            O => \N__45993\,
            I => \delay_measurement_inst.delay_tr_reg3lto9\
        );

    \I__10766\ : CascadeMux
    port map (
            O => \N__45986\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6_cascade_\
        );

    \I__10765\ : InMux
    port map (
            O => \N__45983\,
            I => \N__45980\
        );

    \I__10764\ : LocalMux
    port map (
            O => \N__45980\,
            I => \delay_measurement_inst.delay_tr_timer.N_320_4\
        );

    \I__10763\ : CascadeMux
    port map (
            O => \N__45977\,
            I => \delay_measurement_inst.delay_tr_timer.N_320_4_cascade_\
        );

    \I__10762\ : InMux
    port map (
            O => \N__45974\,
            I => \N__45971\
        );

    \I__10761\ : LocalMux
    port map (
            O => \N__45971\,
            I => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3\
        );

    \I__10760\ : InMux
    port map (
            O => \N__45968\,
            I => \N__45965\
        );

    \I__10759\ : LocalMux
    port map (
            O => \N__45965\,
            I => \N__45961\
        );

    \I__10758\ : InMux
    port map (
            O => \N__45964\,
            I => \N__45958\
        );

    \I__10757\ : Span4Mux_v
    port map (
            O => \N__45961\,
            I => \N__45953\
        );

    \I__10756\ : LocalMux
    port map (
            O => \N__45958\,
            I => \N__45953\
        );

    \I__10755\ : Odrv4
    port map (
            O => \N__45953\,
            I => \delay_measurement_inst.elapsed_time_tr_12\
        );

    \I__10754\ : InMux
    port map (
            O => \N__45950\,
            I => \N__45946\
        );

    \I__10753\ : InMux
    port map (
            O => \N__45949\,
            I => \N__45943\
        );

    \I__10752\ : LocalMux
    port map (
            O => \N__45946\,
            I => \N__45940\
        );

    \I__10751\ : LocalMux
    port map (
            O => \N__45943\,
            I => \N__45937\
        );

    \I__10750\ : Span4Mux_v
    port map (
            O => \N__45940\,
            I => \N__45934\
        );

    \I__10749\ : Span4Mux_h
    port map (
            O => \N__45937\,
            I => \N__45931\
        );

    \I__10748\ : Odrv4
    port map (
            O => \N__45934\,
            I => \delay_measurement_inst.elapsed_time_tr_10\
        );

    \I__10747\ : Odrv4
    port map (
            O => \N__45931\,
            I => \delay_measurement_inst.elapsed_time_tr_10\
        );

    \I__10746\ : InMux
    port map (
            O => \N__45926\,
            I => \N__45922\
        );

    \I__10745\ : InMux
    port map (
            O => \N__45925\,
            I => \N__45919\
        );

    \I__10744\ : LocalMux
    port map (
            O => \N__45922\,
            I => \N__45916\
        );

    \I__10743\ : LocalMux
    port map (
            O => \N__45919\,
            I => \N__45913\
        );

    \I__10742\ : Span4Mux_h
    port map (
            O => \N__45916\,
            I => \N__45909\
        );

    \I__10741\ : Span4Mux_h
    port map (
            O => \N__45913\,
            I => \N__45906\
        );

    \I__10740\ : InMux
    port map (
            O => \N__45912\,
            I => \N__45903\
        );

    \I__10739\ : Odrv4
    port map (
            O => \N__45909\,
            I => \delay_measurement_inst.N_328\
        );

    \I__10738\ : Odrv4
    port map (
            O => \N__45906\,
            I => \delay_measurement_inst.N_328\
        );

    \I__10737\ : LocalMux
    port map (
            O => \N__45903\,
            I => \delay_measurement_inst.N_328\
        );

    \I__10736\ : InMux
    port map (
            O => \N__45896\,
            I => \N__45893\
        );

    \I__10735\ : LocalMux
    port map (
            O => \N__45893\,
            I => \N__45890\
        );

    \I__10734\ : Span4Mux_h
    port map (
            O => \N__45890\,
            I => \N__45886\
        );

    \I__10733\ : InMux
    port map (
            O => \N__45889\,
            I => \N__45883\
        );

    \I__10732\ : Odrv4
    port map (
            O => \N__45886\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__10731\ : LocalMux
    port map (
            O => \N__45883\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__10730\ : InMux
    port map (
            O => \N__45878\,
            I => \N__45875\
        );

    \I__10729\ : LocalMux
    port map (
            O => \N__45875\,
            I => \N__45872\
        );

    \I__10728\ : Span4Mux_v
    port map (
            O => \N__45872\,
            I => \N__45869\
        );

    \I__10727\ : Odrv4
    port map (
            O => \N__45869\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14\
        );

    \I__10726\ : InMux
    port map (
            O => \N__45866\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12\
        );

    \I__10725\ : InMux
    port map (
            O => \N__45863\,
            I => \N__45860\
        );

    \I__10724\ : LocalMux
    port map (
            O => \N__45860\,
            I => \N__45856\
        );

    \I__10723\ : InMux
    port map (
            O => \N__45859\,
            I => \N__45853\
        );

    \I__10722\ : Span4Mux_h
    port map (
            O => \N__45856\,
            I => \N__45850\
        );

    \I__10721\ : LocalMux
    port map (
            O => \N__45853\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__10720\ : Odrv4
    port map (
            O => \N__45850\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__10719\ : InMux
    port map (
            O => \N__45845\,
            I => \N__45842\
        );

    \I__10718\ : LocalMux
    port map (
            O => \N__45842\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15\
        );

    \I__10717\ : InMux
    port map (
            O => \N__45839\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13\
        );

    \I__10716\ : InMux
    port map (
            O => \N__45836\,
            I => \N__45833\
        );

    \I__10715\ : LocalMux
    port map (
            O => \N__45833\,
            I => \N__45829\
        );

    \I__10714\ : InMux
    port map (
            O => \N__45832\,
            I => \N__45826\
        );

    \I__10713\ : Span4Mux_v
    port map (
            O => \N__45829\,
            I => \N__45823\
        );

    \I__10712\ : LocalMux
    port map (
            O => \N__45826\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__10711\ : Odrv4
    port map (
            O => \N__45823\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__10710\ : InMux
    port map (
            O => \N__45818\,
            I => \N__45815\
        );

    \I__10709\ : LocalMux
    port map (
            O => \N__45815\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16\
        );

    \I__10708\ : InMux
    port map (
            O => \N__45812\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14\
        );

    \I__10707\ : InMux
    port map (
            O => \N__45809\,
            I => \N__45806\
        );

    \I__10706\ : LocalMux
    port map (
            O => \N__45806\,
            I => \N__45802\
        );

    \I__10705\ : InMux
    port map (
            O => \N__45805\,
            I => \N__45799\
        );

    \I__10704\ : Span4Mux_h
    port map (
            O => \N__45802\,
            I => \N__45796\
        );

    \I__10703\ : LocalMux
    port map (
            O => \N__45799\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__10702\ : Odrv4
    port map (
            O => \N__45796\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__10701\ : InMux
    port map (
            O => \N__45791\,
            I => \N__45788\
        );

    \I__10700\ : LocalMux
    port map (
            O => \N__45788\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17\
        );

    \I__10699\ : InMux
    port map (
            O => \N__45785\,
            I => \bfn_18_21_0_\
        );

    \I__10698\ : InMux
    port map (
            O => \N__45782\,
            I => \N__45779\
        );

    \I__10697\ : LocalMux
    port map (
            O => \N__45779\,
            I => \N__45775\
        );

    \I__10696\ : InMux
    port map (
            O => \N__45778\,
            I => \N__45772\
        );

    \I__10695\ : Span4Mux_h
    port map (
            O => \N__45775\,
            I => \N__45769\
        );

    \I__10694\ : LocalMux
    port map (
            O => \N__45772\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__10693\ : Odrv4
    port map (
            O => \N__45769\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__10692\ : InMux
    port map (
            O => \N__45764\,
            I => \N__45761\
        );

    \I__10691\ : LocalMux
    port map (
            O => \N__45761\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18\
        );

    \I__10690\ : InMux
    port map (
            O => \N__45758\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16\
        );

    \I__10689\ : InMux
    port map (
            O => \N__45755\,
            I => \N__45752\
        );

    \I__10688\ : LocalMux
    port map (
            O => \N__45752\,
            I => \N__45748\
        );

    \I__10687\ : InMux
    port map (
            O => \N__45751\,
            I => \N__45745\
        );

    \I__10686\ : Span4Mux_h
    port map (
            O => \N__45748\,
            I => \N__45742\
        );

    \I__10685\ : LocalMux
    port map (
            O => \N__45745\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__10684\ : Odrv4
    port map (
            O => \N__45742\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__10683\ : InMux
    port map (
            O => \N__45737\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17\
        );

    \I__10682\ : InMux
    port map (
            O => \N__45734\,
            I => \N__45731\
        );

    \I__10681\ : LocalMux
    port map (
            O => \N__45731\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19\
        );

    \I__10680\ : InMux
    port map (
            O => \N__45728\,
            I => \N__45725\
        );

    \I__10679\ : LocalMux
    port map (
            O => \N__45725\,
            I => \N__45721\
        );

    \I__10678\ : InMux
    port map (
            O => \N__45724\,
            I => \N__45718\
        );

    \I__10677\ : Odrv4
    port map (
            O => \N__45721\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6\
        );

    \I__10676\ : LocalMux
    port map (
            O => \N__45718\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6\
        );

    \I__10675\ : InMux
    port map (
            O => \N__45713\,
            I => \N__45709\
        );

    \I__10674\ : InMux
    port map (
            O => \N__45712\,
            I => \N__45705\
        );

    \I__10673\ : LocalMux
    port map (
            O => \N__45709\,
            I => \N__45702\
        );

    \I__10672\ : InMux
    port map (
            O => \N__45708\,
            I => \N__45699\
        );

    \I__10671\ : LocalMux
    port map (
            O => \N__45705\,
            I => \N__45696\
        );

    \I__10670\ : Span4Mux_h
    port map (
            O => \N__45702\,
            I => \N__45686\
        );

    \I__10669\ : LocalMux
    port map (
            O => \N__45699\,
            I => \N__45686\
        );

    \I__10668\ : Span4Mux_h
    port map (
            O => \N__45696\,
            I => \N__45686\
        );

    \I__10667\ : InMux
    port map (
            O => \N__45695\,
            I => \N__45683\
        );

    \I__10666\ : InMux
    port map (
            O => \N__45694\,
            I => \N__45680\
        );

    \I__10665\ : InMux
    port map (
            O => \N__45693\,
            I => \N__45677\
        );

    \I__10664\ : Odrv4
    port map (
            O => \N__45686\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15\
        );

    \I__10663\ : LocalMux
    port map (
            O => \N__45683\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15\
        );

    \I__10662\ : LocalMux
    port map (
            O => \N__45680\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15\
        );

    \I__10661\ : LocalMux
    port map (
            O => \N__45677\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15\
        );

    \I__10660\ : CascadeMux
    port map (
            O => \N__45668\,
            I => \N__45665\
        );

    \I__10659\ : InMux
    port map (
            O => \N__45665\,
            I => \N__45662\
        );

    \I__10658\ : LocalMux
    port map (
            O => \N__45662\,
            I => \N__45659\
        );

    \I__10657\ : Span4Mux_h
    port map (
            O => \N__45659\,
            I => \N__45656\
        );

    \I__10656\ : Odrv4
    port map (
            O => \N__45656\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6\
        );

    \I__10655\ : InMux
    port map (
            O => \N__45653\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4\
        );

    \I__10654\ : InMux
    port map (
            O => \N__45650\,
            I => \N__45647\
        );

    \I__10653\ : LocalMux
    port map (
            O => \N__45647\,
            I => \N__45644\
        );

    \I__10652\ : Span4Mux_v
    port map (
            O => \N__45644\,
            I => \N__45640\
        );

    \I__10651\ : InMux
    port map (
            O => \N__45643\,
            I => \N__45637\
        );

    \I__10650\ : Odrv4
    port map (
            O => \N__45640\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__10649\ : LocalMux
    port map (
            O => \N__45637\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__10648\ : InMux
    port map (
            O => \N__45632\,
            I => \N__45629\
        );

    \I__10647\ : LocalMux
    port map (
            O => \N__45629\,
            I => \N__45626\
        );

    \I__10646\ : Span4Mux_h
    port map (
            O => \N__45626\,
            I => \N__45623\
        );

    \I__10645\ : Odrv4
    port map (
            O => \N__45623\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7\
        );

    \I__10644\ : InMux
    port map (
            O => \N__45620\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5\
        );

    \I__10643\ : InMux
    port map (
            O => \N__45617\,
            I => \N__45614\
        );

    \I__10642\ : LocalMux
    port map (
            O => \N__45614\,
            I => \N__45611\
        );

    \I__10641\ : Span4Mux_h
    port map (
            O => \N__45611\,
            I => \N__45607\
        );

    \I__10640\ : InMux
    port map (
            O => \N__45610\,
            I => \N__45604\
        );

    \I__10639\ : Odrv4
    port map (
            O => \N__45607\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__10638\ : LocalMux
    port map (
            O => \N__45604\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__10637\ : CascadeMux
    port map (
            O => \N__45599\,
            I => \N__45596\
        );

    \I__10636\ : InMux
    port map (
            O => \N__45596\,
            I => \N__45593\
        );

    \I__10635\ : LocalMux
    port map (
            O => \N__45593\,
            I => \N__45590\
        );

    \I__10634\ : Span4Mux_h
    port map (
            O => \N__45590\,
            I => \N__45587\
        );

    \I__10633\ : Odrv4
    port map (
            O => \N__45587\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8\
        );

    \I__10632\ : InMux
    port map (
            O => \N__45584\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6\
        );

    \I__10631\ : InMux
    port map (
            O => \N__45581\,
            I => \N__45578\
        );

    \I__10630\ : LocalMux
    port map (
            O => \N__45578\,
            I => \N__45574\
        );

    \I__10629\ : InMux
    port map (
            O => \N__45577\,
            I => \N__45571\
        );

    \I__10628\ : Span4Mux_h
    port map (
            O => \N__45574\,
            I => \N__45568\
        );

    \I__10627\ : LocalMux
    port map (
            O => \N__45571\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__10626\ : Odrv4
    port map (
            O => \N__45568\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__10625\ : InMux
    port map (
            O => \N__45563\,
            I => \N__45560\
        );

    \I__10624\ : LocalMux
    port map (
            O => \N__45560\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9\
        );

    \I__10623\ : InMux
    port map (
            O => \N__45557\,
            I => \bfn_18_20_0_\
        );

    \I__10622\ : InMux
    port map (
            O => \N__45554\,
            I => \N__45551\
        );

    \I__10621\ : LocalMux
    port map (
            O => \N__45551\,
            I => \N__45548\
        );

    \I__10620\ : Span4Mux_h
    port map (
            O => \N__45548\,
            I => \N__45544\
        );

    \I__10619\ : InMux
    port map (
            O => \N__45547\,
            I => \N__45541\
        );

    \I__10618\ : Odrv4
    port map (
            O => \N__45544\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__10617\ : LocalMux
    port map (
            O => \N__45541\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__10616\ : CascadeMux
    port map (
            O => \N__45536\,
            I => \N__45533\
        );

    \I__10615\ : InMux
    port map (
            O => \N__45533\,
            I => \N__45530\
        );

    \I__10614\ : LocalMux
    port map (
            O => \N__45530\,
            I => \N__45527\
        );

    \I__10613\ : Span4Mux_h
    port map (
            O => \N__45527\,
            I => \N__45524\
        );

    \I__10612\ : Odrv4
    port map (
            O => \N__45524\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10\
        );

    \I__10611\ : InMux
    port map (
            O => \N__45521\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8\
        );

    \I__10610\ : InMux
    port map (
            O => \N__45518\,
            I => \N__45515\
        );

    \I__10609\ : LocalMux
    port map (
            O => \N__45515\,
            I => \N__45511\
        );

    \I__10608\ : InMux
    port map (
            O => \N__45514\,
            I => \N__45508\
        );

    \I__10607\ : Span4Mux_h
    port map (
            O => \N__45511\,
            I => \N__45505\
        );

    \I__10606\ : LocalMux
    port map (
            O => \N__45508\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__10605\ : Odrv4
    port map (
            O => \N__45505\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__10604\ : InMux
    port map (
            O => \N__45500\,
            I => \N__45497\
        );

    \I__10603\ : LocalMux
    port map (
            O => \N__45497\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11\
        );

    \I__10602\ : InMux
    port map (
            O => \N__45494\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9\
        );

    \I__10601\ : InMux
    port map (
            O => \N__45491\,
            I => \N__45488\
        );

    \I__10600\ : LocalMux
    port map (
            O => \N__45488\,
            I => \N__45484\
        );

    \I__10599\ : InMux
    port map (
            O => \N__45487\,
            I => \N__45481\
        );

    \I__10598\ : Span4Mux_h
    port map (
            O => \N__45484\,
            I => \N__45478\
        );

    \I__10597\ : LocalMux
    port map (
            O => \N__45481\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__10596\ : Odrv4
    port map (
            O => \N__45478\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__10595\ : InMux
    port map (
            O => \N__45473\,
            I => \N__45470\
        );

    \I__10594\ : LocalMux
    port map (
            O => \N__45470\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12\
        );

    \I__10593\ : InMux
    port map (
            O => \N__45467\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10\
        );

    \I__10592\ : InMux
    port map (
            O => \N__45464\,
            I => \N__45461\
        );

    \I__10591\ : LocalMux
    port map (
            O => \N__45461\,
            I => \N__45457\
        );

    \I__10590\ : InMux
    port map (
            O => \N__45460\,
            I => \N__45454\
        );

    \I__10589\ : Span4Mux_v
    port map (
            O => \N__45457\,
            I => \N__45451\
        );

    \I__10588\ : LocalMux
    port map (
            O => \N__45454\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__10587\ : Odrv4
    port map (
            O => \N__45451\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__10586\ : InMux
    port map (
            O => \N__45446\,
            I => \N__45443\
        );

    \I__10585\ : LocalMux
    port map (
            O => \N__45443\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13\
        );

    \I__10584\ : InMux
    port map (
            O => \N__45440\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11\
        );

    \I__10583\ : InMux
    port map (
            O => \N__45437\,
            I => \N__45430\
        );

    \I__10582\ : InMux
    port map (
            O => \N__45436\,
            I => \N__45430\
        );

    \I__10581\ : InMux
    port map (
            O => \N__45435\,
            I => \N__45427\
        );

    \I__10580\ : LocalMux
    port map (
            O => \N__45430\,
            I => \N__45424\
        );

    \I__10579\ : LocalMux
    port map (
            O => \N__45427\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__10578\ : Odrv4
    port map (
            O => \N__45424\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__10577\ : CascadeMux
    port map (
            O => \N__45419\,
            I => \N__45416\
        );

    \I__10576\ : InMux
    port map (
            O => \N__45416\,
            I => \N__45412\
        );

    \I__10575\ : InMux
    port map (
            O => \N__45415\,
            I => \N__45409\
        );

    \I__10574\ : LocalMux
    port map (
            O => \N__45412\,
            I => \N__45406\
        );

    \I__10573\ : LocalMux
    port map (
            O => \N__45409\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__10572\ : Odrv4
    port map (
            O => \N__45406\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__10571\ : InMux
    port map (
            O => \N__45401\,
            I => \N__45398\
        );

    \I__10570\ : LocalMux
    port map (
            O => \N__45398\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30\
        );

    \I__10569\ : InMux
    port map (
            O => \N__45395\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__10568\ : InMux
    port map (
            O => \N__45392\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__10567\ : CEMux
    port map (
            O => \N__45389\,
            I => \N__45384\
        );

    \I__10566\ : CEMux
    port map (
            O => \N__45388\,
            I => \N__45381\
        );

    \I__10565\ : CEMux
    port map (
            O => \N__45387\,
            I => \N__45378\
        );

    \I__10564\ : LocalMux
    port map (
            O => \N__45384\,
            I => \N__45374\
        );

    \I__10563\ : LocalMux
    port map (
            O => \N__45381\,
            I => \N__45370\
        );

    \I__10562\ : LocalMux
    port map (
            O => \N__45378\,
            I => \N__45367\
        );

    \I__10561\ : CEMux
    port map (
            O => \N__45377\,
            I => \N__45364\
        );

    \I__10560\ : Span4Mux_v
    port map (
            O => \N__45374\,
            I => \N__45361\
        );

    \I__10559\ : CEMux
    port map (
            O => \N__45373\,
            I => \N__45358\
        );

    \I__10558\ : Span4Mux_v
    port map (
            O => \N__45370\,
            I => \N__45347\
        );

    \I__10557\ : Span4Mux_v
    port map (
            O => \N__45367\,
            I => \N__45347\
        );

    \I__10556\ : LocalMux
    port map (
            O => \N__45364\,
            I => \N__45347\
        );

    \I__10555\ : Span4Mux_v
    port map (
            O => \N__45361\,
            I => \N__45347\
        );

    \I__10554\ : LocalMux
    port map (
            O => \N__45358\,
            I => \N__45347\
        );

    \I__10553\ : Span4Mux_v
    port map (
            O => \N__45347\,
            I => \N__45344\
        );

    \I__10552\ : Span4Mux_h
    port map (
            O => \N__45344\,
            I => \N__45341\
        );

    \I__10551\ : Odrv4
    port map (
            O => \N__45341\,
            I => \delay_measurement_inst.delay_tr_timer.N_337_i\
        );

    \I__10550\ : InMux
    port map (
            O => \N__45338\,
            I => \N__45335\
        );

    \I__10549\ : LocalMux
    port map (
            O => \N__45335\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1\
        );

    \I__10548\ : CascadeMux
    port map (
            O => \N__45332\,
            I => \N__45329\
        );

    \I__10547\ : InMux
    port map (
            O => \N__45329\,
            I => \N__45324\
        );

    \I__10546\ : InMux
    port map (
            O => \N__45328\,
            I => \N__45321\
        );

    \I__10545\ : InMux
    port map (
            O => \N__45327\,
            I => \N__45318\
        );

    \I__10544\ : LocalMux
    port map (
            O => \N__45324\,
            I => \N__45315\
        );

    \I__10543\ : LocalMux
    port map (
            O => \N__45321\,
            I => \N__45310\
        );

    \I__10542\ : LocalMux
    port map (
            O => \N__45318\,
            I => \N__45310\
        );

    \I__10541\ : Span4Mux_h
    port map (
            O => \N__45315\,
            I => \N__45305\
        );

    \I__10540\ : Span4Mux_v
    port map (
            O => \N__45310\,
            I => \N__45305\
        );

    \I__10539\ : Odrv4
    port map (
            O => \N__45305\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__10538\ : InMux
    port map (
            O => \N__45302\,
            I => \N__45299\
        );

    \I__10537\ : LocalMux
    port map (
            O => \N__45299\,
            I => \N__45296\
        );

    \I__10536\ : Span4Mux_h
    port map (
            O => \N__45296\,
            I => \N__45292\
        );

    \I__10535\ : InMux
    port map (
            O => \N__45295\,
            I => \N__45289\
        );

    \I__10534\ : Odrv4
    port map (
            O => \N__45292\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__10533\ : LocalMux
    port map (
            O => \N__45289\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__10532\ : InMux
    port map (
            O => \N__45284\,
            I => \N__45281\
        );

    \I__10531\ : LocalMux
    port map (
            O => \N__45281\,
            I => \N__45278\
        );

    \I__10530\ : Span4Mux_h
    port map (
            O => \N__45278\,
            I => \N__45275\
        );

    \I__10529\ : Odrv4
    port map (
            O => \N__45275\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2\
        );

    \I__10528\ : InMux
    port map (
            O => \N__45272\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0\
        );

    \I__10527\ : InMux
    port map (
            O => \N__45269\,
            I => \N__45266\
        );

    \I__10526\ : LocalMux
    port map (
            O => \N__45266\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0\
        );

    \I__10525\ : CascadeMux
    port map (
            O => \N__45263\,
            I => \N__45260\
        );

    \I__10524\ : InMux
    port map (
            O => \N__45260\,
            I => \N__45257\
        );

    \I__10523\ : LocalMux
    port map (
            O => \N__45257\,
            I => \N__45254\
        );

    \I__10522\ : Span4Mux_v
    port map (
            O => \N__45254\,
            I => \N__45250\
        );

    \I__10521\ : InMux
    port map (
            O => \N__45253\,
            I => \N__45247\
        );

    \I__10520\ : Odrv4
    port map (
            O => \N__45250\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__10519\ : LocalMux
    port map (
            O => \N__45247\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__10518\ : InMux
    port map (
            O => \N__45242\,
            I => \N__45239\
        );

    \I__10517\ : LocalMux
    port map (
            O => \N__45239\,
            I => \N__45236\
        );

    \I__10516\ : Span12Mux_h
    port map (
            O => \N__45236\,
            I => \N__45233\
        );

    \I__10515\ : Odrv12
    port map (
            O => \N__45233\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3\
        );

    \I__10514\ : InMux
    port map (
            O => \N__45230\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1\
        );

    \I__10513\ : InMux
    port map (
            O => \N__45227\,
            I => \N__45224\
        );

    \I__10512\ : LocalMux
    port map (
            O => \N__45224\,
            I => \N__45221\
        );

    \I__10511\ : Span4Mux_h
    port map (
            O => \N__45221\,
            I => \N__45217\
        );

    \I__10510\ : InMux
    port map (
            O => \N__45220\,
            I => \N__45214\
        );

    \I__10509\ : Odrv4
    port map (
            O => \N__45217\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__10508\ : LocalMux
    port map (
            O => \N__45214\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__10507\ : InMux
    port map (
            O => \N__45209\,
            I => \N__45206\
        );

    \I__10506\ : LocalMux
    port map (
            O => \N__45206\,
            I => \N__45203\
        );

    \I__10505\ : Span4Mux_v
    port map (
            O => \N__45203\,
            I => \N__45200\
        );

    \I__10504\ : Odrv4
    port map (
            O => \N__45200\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4\
        );

    \I__10503\ : InMux
    port map (
            O => \N__45197\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2\
        );

    \I__10502\ : InMux
    port map (
            O => \N__45194\,
            I => \N__45191\
        );

    \I__10501\ : LocalMux
    port map (
            O => \N__45191\,
            I => \N__45188\
        );

    \I__10500\ : Span4Mux_v
    port map (
            O => \N__45188\,
            I => \N__45184\
        );

    \I__10499\ : InMux
    port map (
            O => \N__45187\,
            I => \N__45181\
        );

    \I__10498\ : Odrv4
    port map (
            O => \N__45184\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__10497\ : LocalMux
    port map (
            O => \N__45181\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__10496\ : CascadeMux
    port map (
            O => \N__45176\,
            I => \N__45173\
        );

    \I__10495\ : InMux
    port map (
            O => \N__45173\,
            I => \N__45170\
        );

    \I__10494\ : LocalMux
    port map (
            O => \N__45170\,
            I => \N__45167\
        );

    \I__10493\ : Span4Mux_h
    port map (
            O => \N__45167\,
            I => \N__45164\
        );

    \I__10492\ : Odrv4
    port map (
            O => \N__45164\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5\
        );

    \I__10491\ : InMux
    port map (
            O => \N__45161\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3\
        );

    \I__10490\ : InMux
    port map (
            O => \N__45158\,
            I => \N__45155\
        );

    \I__10489\ : LocalMux
    port map (
            O => \N__45155\,
            I => \N__45152\
        );

    \I__10488\ : Span4Mux_h
    port map (
            O => \N__45152\,
            I => \N__45148\
        );

    \I__10487\ : InMux
    port map (
            O => \N__45151\,
            I => \N__45145\
        );

    \I__10486\ : Odrv4
    port map (
            O => \N__45148\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__10485\ : LocalMux
    port map (
            O => \N__45145\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__10484\ : CascadeMux
    port map (
            O => \N__45140\,
            I => \N__45136\
        );

    \I__10483\ : CascadeMux
    port map (
            O => \N__45139\,
            I => \N__45133\
        );

    \I__10482\ : InMux
    port map (
            O => \N__45136\,
            I => \N__45127\
        );

    \I__10481\ : InMux
    port map (
            O => \N__45133\,
            I => \N__45127\
        );

    \I__10480\ : InMux
    port map (
            O => \N__45132\,
            I => \N__45124\
        );

    \I__10479\ : LocalMux
    port map (
            O => \N__45127\,
            I => \N__45121\
        );

    \I__10478\ : LocalMux
    port map (
            O => \N__45124\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__10477\ : Odrv4
    port map (
            O => \N__45121\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__10476\ : InMux
    port map (
            O => \N__45116\,
            I => \N__45113\
        );

    \I__10475\ : LocalMux
    port map (
            O => \N__45113\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__10474\ : InMux
    port map (
            O => \N__45110\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__10473\ : InMux
    port map (
            O => \N__45107\,
            I => \N__45101\
        );

    \I__10472\ : InMux
    port map (
            O => \N__45106\,
            I => \N__45101\
        );

    \I__10471\ : LocalMux
    port map (
            O => \N__45101\,
            I => \N__45097\
        );

    \I__10470\ : InMux
    port map (
            O => \N__45100\,
            I => \N__45094\
        );

    \I__10469\ : Span4Mux_h
    port map (
            O => \N__45097\,
            I => \N__45091\
        );

    \I__10468\ : LocalMux
    port map (
            O => \N__45094\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__10467\ : Odrv4
    port map (
            O => \N__45091\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__10466\ : InMux
    port map (
            O => \N__45086\,
            I => \N__45083\
        );

    \I__10465\ : LocalMux
    port map (
            O => \N__45083\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__10464\ : InMux
    port map (
            O => \N__45080\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__10463\ : CascadeMux
    port map (
            O => \N__45077\,
            I => \N__45074\
        );

    \I__10462\ : InMux
    port map (
            O => \N__45074\,
            I => \N__45070\
        );

    \I__10461\ : InMux
    port map (
            O => \N__45073\,
            I => \N__45067\
        );

    \I__10460\ : LocalMux
    port map (
            O => \N__45070\,
            I => \N__45061\
        );

    \I__10459\ : LocalMux
    port map (
            O => \N__45067\,
            I => \N__45061\
        );

    \I__10458\ : InMux
    port map (
            O => \N__45066\,
            I => \N__45058\
        );

    \I__10457\ : Span4Mux_v
    port map (
            O => \N__45061\,
            I => \N__45055\
        );

    \I__10456\ : LocalMux
    port map (
            O => \N__45058\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__10455\ : Odrv4
    port map (
            O => \N__45055\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__10454\ : CascadeMux
    port map (
            O => \N__45050\,
            I => \N__45047\
        );

    \I__10453\ : InMux
    port map (
            O => \N__45047\,
            I => \N__45044\
        );

    \I__10452\ : LocalMux
    port map (
            O => \N__45044\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__10451\ : InMux
    port map (
            O => \N__45041\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__10450\ : CascadeMux
    port map (
            O => \N__45038\,
            I => \N__45034\
        );

    \I__10449\ : InMux
    port map (
            O => \N__45037\,
            I => \N__45031\
        );

    \I__10448\ : InMux
    port map (
            O => \N__45034\,
            I => \N__45028\
        );

    \I__10447\ : LocalMux
    port map (
            O => \N__45031\,
            I => \N__45022\
        );

    \I__10446\ : LocalMux
    port map (
            O => \N__45028\,
            I => \N__45022\
        );

    \I__10445\ : InMux
    port map (
            O => \N__45027\,
            I => \N__45019\
        );

    \I__10444\ : Span4Mux_v
    port map (
            O => \N__45022\,
            I => \N__45016\
        );

    \I__10443\ : LocalMux
    port map (
            O => \N__45019\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__10442\ : Odrv4
    port map (
            O => \N__45016\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__10441\ : InMux
    port map (
            O => \N__45011\,
            I => \N__45008\
        );

    \I__10440\ : LocalMux
    port map (
            O => \N__45008\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__10439\ : InMux
    port map (
            O => \N__45005\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__10438\ : InMux
    port map (
            O => \N__45002\,
            I => \N__44995\
        );

    \I__10437\ : InMux
    port map (
            O => \N__45001\,
            I => \N__44995\
        );

    \I__10436\ : InMux
    port map (
            O => \N__45000\,
            I => \N__44992\
        );

    \I__10435\ : LocalMux
    port map (
            O => \N__44995\,
            I => \N__44989\
        );

    \I__10434\ : LocalMux
    port map (
            O => \N__44992\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__10433\ : Odrv4
    port map (
            O => \N__44989\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__10432\ : InMux
    port map (
            O => \N__44984\,
            I => \N__44981\
        );

    \I__10431\ : LocalMux
    port map (
            O => \N__44981\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__10430\ : InMux
    port map (
            O => \N__44978\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__10429\ : InMux
    port map (
            O => \N__44975\,
            I => \N__44972\
        );

    \I__10428\ : LocalMux
    port map (
            O => \N__44972\,
            I => \N__44968\
        );

    \I__10427\ : CascadeMux
    port map (
            O => \N__44971\,
            I => \N__44964\
        );

    \I__10426\ : Span4Mux_h
    port map (
            O => \N__44968\,
            I => \N__44961\
        );

    \I__10425\ : InMux
    port map (
            O => \N__44967\,
            I => \N__44958\
        );

    \I__10424\ : InMux
    port map (
            O => \N__44964\,
            I => \N__44955\
        );

    \I__10423\ : Odrv4
    port map (
            O => \N__44961\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__10422\ : LocalMux
    port map (
            O => \N__44958\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__10421\ : LocalMux
    port map (
            O => \N__44955\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__10420\ : InMux
    port map (
            O => \N__44948\,
            I => \N__44945\
        );

    \I__10419\ : LocalMux
    port map (
            O => \N__44945\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__10418\ : InMux
    port map (
            O => \N__44942\,
            I => \bfn_18_18_0_\
        );

    \I__10417\ : CascadeMux
    port map (
            O => \N__44939\,
            I => \N__44936\
        );

    \I__10416\ : InMux
    port map (
            O => \N__44936\,
            I => \N__44933\
        );

    \I__10415\ : LocalMux
    port map (
            O => \N__44933\,
            I => \N__44928\
        );

    \I__10414\ : CascadeMux
    port map (
            O => \N__44932\,
            I => \N__44925\
        );

    \I__10413\ : InMux
    port map (
            O => \N__44931\,
            I => \N__44922\
        );

    \I__10412\ : Span4Mux_h
    port map (
            O => \N__44928\,
            I => \N__44919\
        );

    \I__10411\ : InMux
    port map (
            O => \N__44925\,
            I => \N__44916\
        );

    \I__10410\ : LocalMux
    port map (
            O => \N__44922\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__10409\ : Odrv4
    port map (
            O => \N__44919\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__10408\ : LocalMux
    port map (
            O => \N__44916\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__10407\ : CascadeMux
    port map (
            O => \N__44909\,
            I => \N__44906\
        );

    \I__10406\ : InMux
    port map (
            O => \N__44906\,
            I => \N__44903\
        );

    \I__10405\ : LocalMux
    port map (
            O => \N__44903\,
            I => \N__44900\
        );

    \I__10404\ : Odrv4
    port map (
            O => \N__44900\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__10403\ : InMux
    port map (
            O => \N__44897\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__10402\ : InMux
    port map (
            O => \N__44894\,
            I => \N__44890\
        );

    \I__10401\ : InMux
    port map (
            O => \N__44893\,
            I => \N__44887\
        );

    \I__10400\ : LocalMux
    port map (
            O => \N__44890\,
            I => \N__44884\
        );

    \I__10399\ : LocalMux
    port map (
            O => \N__44887\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__10398\ : Odrv4
    port map (
            O => \N__44884\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__10397\ : CascadeMux
    port map (
            O => \N__44879\,
            I => \N__44875\
        );

    \I__10396\ : CascadeMux
    port map (
            O => \N__44878\,
            I => \N__44872\
        );

    \I__10395\ : InMux
    port map (
            O => \N__44875\,
            I => \N__44866\
        );

    \I__10394\ : InMux
    port map (
            O => \N__44872\,
            I => \N__44866\
        );

    \I__10393\ : InMux
    port map (
            O => \N__44871\,
            I => \N__44863\
        );

    \I__10392\ : LocalMux
    port map (
            O => \N__44866\,
            I => \N__44860\
        );

    \I__10391\ : LocalMux
    port map (
            O => \N__44863\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__10390\ : Odrv4
    port map (
            O => \N__44860\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__10389\ : InMux
    port map (
            O => \N__44855\,
            I => \N__44852\
        );

    \I__10388\ : LocalMux
    port map (
            O => \N__44852\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__10387\ : InMux
    port map (
            O => \N__44849\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__10386\ : CascadeMux
    port map (
            O => \N__44846\,
            I => \N__44842\
        );

    \I__10385\ : InMux
    port map (
            O => \N__44845\,
            I => \N__44839\
        );

    \I__10384\ : InMux
    port map (
            O => \N__44842\,
            I => \N__44836\
        );

    \I__10383\ : LocalMux
    port map (
            O => \N__44839\,
            I => \N__44830\
        );

    \I__10382\ : LocalMux
    port map (
            O => \N__44836\,
            I => \N__44830\
        );

    \I__10381\ : InMux
    port map (
            O => \N__44835\,
            I => \N__44827\
        );

    \I__10380\ : Span4Mux_v
    port map (
            O => \N__44830\,
            I => \N__44824\
        );

    \I__10379\ : LocalMux
    port map (
            O => \N__44827\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__10378\ : Odrv4
    port map (
            O => \N__44824\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__10377\ : InMux
    port map (
            O => \N__44819\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__10376\ : CascadeMux
    port map (
            O => \N__44816\,
            I => \N__44812\
        );

    \I__10375\ : CascadeMux
    port map (
            O => \N__44815\,
            I => \N__44809\
        );

    \I__10374\ : InMux
    port map (
            O => \N__44812\,
            I => \N__44803\
        );

    \I__10373\ : InMux
    port map (
            O => \N__44809\,
            I => \N__44803\
        );

    \I__10372\ : InMux
    port map (
            O => \N__44808\,
            I => \N__44800\
        );

    \I__10371\ : LocalMux
    port map (
            O => \N__44803\,
            I => \N__44797\
        );

    \I__10370\ : LocalMux
    port map (
            O => \N__44800\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__10369\ : Odrv4
    port map (
            O => \N__44797\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__10368\ : InMux
    port map (
            O => \N__44792\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__10367\ : CascadeMux
    port map (
            O => \N__44789\,
            I => \N__44785\
        );

    \I__10366\ : CascadeMux
    port map (
            O => \N__44788\,
            I => \N__44782\
        );

    \I__10365\ : InMux
    port map (
            O => \N__44785\,
            I => \N__44776\
        );

    \I__10364\ : InMux
    port map (
            O => \N__44782\,
            I => \N__44776\
        );

    \I__10363\ : InMux
    port map (
            O => \N__44781\,
            I => \N__44773\
        );

    \I__10362\ : LocalMux
    port map (
            O => \N__44776\,
            I => \N__44770\
        );

    \I__10361\ : LocalMux
    port map (
            O => \N__44773\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__10360\ : Odrv4
    port map (
            O => \N__44770\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__10359\ : InMux
    port map (
            O => \N__44765\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__10358\ : InMux
    port map (
            O => \N__44762\,
            I => \N__44755\
        );

    \I__10357\ : InMux
    port map (
            O => \N__44761\,
            I => \N__44755\
        );

    \I__10356\ : InMux
    port map (
            O => \N__44760\,
            I => \N__44752\
        );

    \I__10355\ : LocalMux
    port map (
            O => \N__44755\,
            I => \N__44749\
        );

    \I__10354\ : LocalMux
    port map (
            O => \N__44752\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__10353\ : Odrv4
    port map (
            O => \N__44749\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__10352\ : InMux
    port map (
            O => \N__44744\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__10351\ : InMux
    port map (
            O => \N__44741\,
            I => \N__44734\
        );

    \I__10350\ : InMux
    port map (
            O => \N__44740\,
            I => \N__44734\
        );

    \I__10349\ : InMux
    port map (
            O => \N__44739\,
            I => \N__44731\
        );

    \I__10348\ : LocalMux
    port map (
            O => \N__44734\,
            I => \N__44728\
        );

    \I__10347\ : LocalMux
    port map (
            O => \N__44731\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__10346\ : Odrv4
    port map (
            O => \N__44728\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__10345\ : InMux
    port map (
            O => \N__44723\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__10344\ : CascadeMux
    port map (
            O => \N__44720\,
            I => \N__44716\
        );

    \I__10343\ : InMux
    port map (
            O => \N__44719\,
            I => \N__44712\
        );

    \I__10342\ : InMux
    port map (
            O => \N__44716\,
            I => \N__44709\
        );

    \I__10341\ : InMux
    port map (
            O => \N__44715\,
            I => \N__44706\
        );

    \I__10340\ : LocalMux
    port map (
            O => \N__44712\,
            I => \N__44701\
        );

    \I__10339\ : LocalMux
    port map (
            O => \N__44709\,
            I => \N__44701\
        );

    \I__10338\ : LocalMux
    port map (
            O => \N__44706\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__10337\ : Odrv4
    port map (
            O => \N__44701\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__10336\ : InMux
    port map (
            O => \N__44696\,
            I => \bfn_18_17_0_\
        );

    \I__10335\ : InMux
    port map (
            O => \N__44693\,
            I => \N__44689\
        );

    \I__10334\ : CascadeMux
    port map (
            O => \N__44692\,
            I => \N__44685\
        );

    \I__10333\ : LocalMux
    port map (
            O => \N__44689\,
            I => \N__44682\
        );

    \I__10332\ : InMux
    port map (
            O => \N__44688\,
            I => \N__44679\
        );

    \I__10331\ : InMux
    port map (
            O => \N__44685\,
            I => \N__44676\
        );

    \I__10330\ : Odrv4
    port map (
            O => \N__44682\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__10329\ : LocalMux
    port map (
            O => \N__44679\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__10328\ : LocalMux
    port map (
            O => \N__44676\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__10327\ : InMux
    port map (
            O => \N__44669\,
            I => \N__44666\
        );

    \I__10326\ : LocalMux
    port map (
            O => \N__44666\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__10325\ : InMux
    port map (
            O => \N__44663\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__10324\ : CascadeMux
    port map (
            O => \N__44660\,
            I => \N__44656\
        );

    \I__10323\ : CascadeMux
    port map (
            O => \N__44659\,
            I => \N__44653\
        );

    \I__10322\ : InMux
    port map (
            O => \N__44656\,
            I => \N__44647\
        );

    \I__10321\ : InMux
    port map (
            O => \N__44653\,
            I => \N__44647\
        );

    \I__10320\ : InMux
    port map (
            O => \N__44652\,
            I => \N__44644\
        );

    \I__10319\ : LocalMux
    port map (
            O => \N__44647\,
            I => \N__44641\
        );

    \I__10318\ : LocalMux
    port map (
            O => \N__44644\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__10317\ : Odrv4
    port map (
            O => \N__44641\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__10316\ : InMux
    port map (
            O => \N__44636\,
            I => \N__44633\
        );

    \I__10315\ : LocalMux
    port map (
            O => \N__44633\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__10314\ : InMux
    port map (
            O => \N__44630\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__10313\ : CascadeMux
    port map (
            O => \N__44627\,
            I => \N__44623\
        );

    \I__10312\ : CascadeMux
    port map (
            O => \N__44626\,
            I => \N__44620\
        );

    \I__10311\ : InMux
    port map (
            O => \N__44623\,
            I => \N__44614\
        );

    \I__10310\ : InMux
    port map (
            O => \N__44620\,
            I => \N__44614\
        );

    \I__10309\ : InMux
    port map (
            O => \N__44619\,
            I => \N__44611\
        );

    \I__10308\ : LocalMux
    port map (
            O => \N__44614\,
            I => \N__44608\
        );

    \I__10307\ : LocalMux
    port map (
            O => \N__44611\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__10306\ : Odrv4
    port map (
            O => \N__44608\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__10305\ : InMux
    port map (
            O => \N__44603\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__10304\ : CascadeMux
    port map (
            O => \N__44600\,
            I => \N__44596\
        );

    \I__10303\ : CascadeMux
    port map (
            O => \N__44599\,
            I => \N__44593\
        );

    \I__10302\ : InMux
    port map (
            O => \N__44596\,
            I => \N__44587\
        );

    \I__10301\ : InMux
    port map (
            O => \N__44593\,
            I => \N__44587\
        );

    \I__10300\ : InMux
    port map (
            O => \N__44592\,
            I => \N__44584\
        );

    \I__10299\ : LocalMux
    port map (
            O => \N__44587\,
            I => \N__44581\
        );

    \I__10298\ : LocalMux
    port map (
            O => \N__44584\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__10297\ : Odrv4
    port map (
            O => \N__44581\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__10296\ : InMux
    port map (
            O => \N__44576\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__10295\ : InMux
    port map (
            O => \N__44573\,
            I => \N__44567\
        );

    \I__10294\ : InMux
    port map (
            O => \N__44572\,
            I => \N__44567\
        );

    \I__10293\ : LocalMux
    port map (
            O => \N__44567\,
            I => \N__44563\
        );

    \I__10292\ : InMux
    port map (
            O => \N__44566\,
            I => \N__44560\
        );

    \I__10291\ : Span4Mux_h
    port map (
            O => \N__44563\,
            I => \N__44557\
        );

    \I__10290\ : LocalMux
    port map (
            O => \N__44560\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__10289\ : Odrv4
    port map (
            O => \N__44557\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__10288\ : InMux
    port map (
            O => \N__44552\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__10287\ : InMux
    port map (
            O => \N__44549\,
            I => \N__44543\
        );

    \I__10286\ : InMux
    port map (
            O => \N__44548\,
            I => \N__44543\
        );

    \I__10285\ : LocalMux
    port map (
            O => \N__44543\,
            I => \N__44539\
        );

    \I__10284\ : InMux
    port map (
            O => \N__44542\,
            I => \N__44536\
        );

    \I__10283\ : Span4Mux_h
    port map (
            O => \N__44539\,
            I => \N__44533\
        );

    \I__10282\ : LocalMux
    port map (
            O => \N__44536\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__10281\ : Odrv4
    port map (
            O => \N__44533\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__10280\ : InMux
    port map (
            O => \N__44528\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__10279\ : CascadeMux
    port map (
            O => \N__44525\,
            I => \N__44521\
        );

    \I__10278\ : InMux
    port map (
            O => \N__44524\,
            I => \N__44518\
        );

    \I__10277\ : InMux
    port map (
            O => \N__44521\,
            I => \N__44515\
        );

    \I__10276\ : LocalMux
    port map (
            O => \N__44518\,
            I => \N__44509\
        );

    \I__10275\ : LocalMux
    port map (
            O => \N__44515\,
            I => \N__44509\
        );

    \I__10274\ : InMux
    port map (
            O => \N__44514\,
            I => \N__44506\
        );

    \I__10273\ : Span4Mux_v
    port map (
            O => \N__44509\,
            I => \N__44503\
        );

    \I__10272\ : LocalMux
    port map (
            O => \N__44506\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__10271\ : Odrv4
    port map (
            O => \N__44503\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__10270\ : InMux
    port map (
            O => \N__44498\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__10269\ : CascadeMux
    port map (
            O => \N__44495\,
            I => \N__44491\
        );

    \I__10268\ : CascadeMux
    port map (
            O => \N__44494\,
            I => \N__44488\
        );

    \I__10267\ : InMux
    port map (
            O => \N__44491\,
            I => \N__44483\
        );

    \I__10266\ : InMux
    port map (
            O => \N__44488\,
            I => \N__44483\
        );

    \I__10265\ : LocalMux
    port map (
            O => \N__44483\,
            I => \N__44479\
        );

    \I__10264\ : InMux
    port map (
            O => \N__44482\,
            I => \N__44476\
        );

    \I__10263\ : Span4Mux_v
    port map (
            O => \N__44479\,
            I => \N__44473\
        );

    \I__10262\ : LocalMux
    port map (
            O => \N__44476\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__10261\ : Odrv4
    port map (
            O => \N__44473\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__10260\ : InMux
    port map (
            O => \N__44468\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__10259\ : InMux
    port map (
            O => \N__44465\,
            I => \N__44462\
        );

    \I__10258\ : LocalMux
    port map (
            O => \N__44462\,
            I => \N__44458\
        );

    \I__10257\ : CascadeMux
    port map (
            O => \N__44461\,
            I => \N__44454\
        );

    \I__10256\ : Span4Mux_h
    port map (
            O => \N__44458\,
            I => \N__44451\
        );

    \I__10255\ : InMux
    port map (
            O => \N__44457\,
            I => \N__44448\
        );

    \I__10254\ : InMux
    port map (
            O => \N__44454\,
            I => \N__44445\
        );

    \I__10253\ : Odrv4
    port map (
            O => \N__44451\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__10252\ : LocalMux
    port map (
            O => \N__44448\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__10251\ : LocalMux
    port map (
            O => \N__44445\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__10250\ : InMux
    port map (
            O => \N__44438\,
            I => \bfn_18_16_0_\
        );

    \I__10249\ : InMux
    port map (
            O => \N__44435\,
            I => \N__44432\
        );

    \I__10248\ : LocalMux
    port map (
            O => \N__44432\,
            I => \N__44427\
        );

    \I__10247\ : InMux
    port map (
            O => \N__44431\,
            I => \N__44424\
        );

    \I__10246\ : InMux
    port map (
            O => \N__44430\,
            I => \N__44421\
        );

    \I__10245\ : Odrv4
    port map (
            O => \N__44427\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__10244\ : LocalMux
    port map (
            O => \N__44424\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__10243\ : LocalMux
    port map (
            O => \N__44421\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__10242\ : InMux
    port map (
            O => \N__44414\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__10241\ : CascadeMux
    port map (
            O => \N__44411\,
            I => \N__44407\
        );

    \I__10240\ : InMux
    port map (
            O => \N__44410\,
            I => \N__44404\
        );

    \I__10239\ : InMux
    port map (
            O => \N__44407\,
            I => \N__44401\
        );

    \I__10238\ : LocalMux
    port map (
            O => \N__44404\,
            I => \N__44395\
        );

    \I__10237\ : LocalMux
    port map (
            O => \N__44401\,
            I => \N__44395\
        );

    \I__10236\ : InMux
    port map (
            O => \N__44400\,
            I => \N__44392\
        );

    \I__10235\ : Span4Mux_v
    port map (
            O => \N__44395\,
            I => \N__44389\
        );

    \I__10234\ : LocalMux
    port map (
            O => \N__44392\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__10233\ : Odrv4
    port map (
            O => \N__44389\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__10232\ : InMux
    port map (
            O => \N__44384\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__10231\ : InMux
    port map (
            O => \N__44381\,
            I => \N__44378\
        );

    \I__10230\ : LocalMux
    port map (
            O => \N__44378\,
            I => \N__44375\
        );

    \I__10229\ : Span4Mux_h
    port map (
            O => \N__44375\,
            I => \N__44370\
        );

    \I__10228\ : InMux
    port map (
            O => \N__44374\,
            I => \N__44367\
        );

    \I__10227\ : InMux
    port map (
            O => \N__44373\,
            I => \N__44364\
        );

    \I__10226\ : Odrv4
    port map (
            O => \N__44370\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__10225\ : LocalMux
    port map (
            O => \N__44367\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__10224\ : LocalMux
    port map (
            O => \N__44364\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__10223\ : InMux
    port map (
            O => \N__44357\,
            I => \N__44352\
        );

    \I__10222\ : InMux
    port map (
            O => \N__44356\,
            I => \N__44349\
        );

    \I__10221\ : InMux
    port map (
            O => \N__44355\,
            I => \N__44346\
        );

    \I__10220\ : LocalMux
    port map (
            O => \N__44352\,
            I => \N__44341\
        );

    \I__10219\ : LocalMux
    port map (
            O => \N__44349\,
            I => \N__44341\
        );

    \I__10218\ : LocalMux
    port map (
            O => \N__44346\,
            I => \N__44336\
        );

    \I__10217\ : Span4Mux_v
    port map (
            O => \N__44341\,
            I => \N__44336\
        );

    \I__10216\ : Odrv4
    port map (
            O => \N__44336\,
            I => \delay_measurement_inst.elapsed_time_hc_2\
        );

    \I__10215\ : CEMux
    port map (
            O => \N__44333\,
            I => \N__44315\
        );

    \I__10214\ : CEMux
    port map (
            O => \N__44332\,
            I => \N__44315\
        );

    \I__10213\ : CEMux
    port map (
            O => \N__44331\,
            I => \N__44315\
        );

    \I__10212\ : CEMux
    port map (
            O => \N__44330\,
            I => \N__44315\
        );

    \I__10211\ : CEMux
    port map (
            O => \N__44329\,
            I => \N__44315\
        );

    \I__10210\ : CEMux
    port map (
            O => \N__44328\,
            I => \N__44315\
        );

    \I__10209\ : GlobalMux
    port map (
            O => \N__44315\,
            I => \N__44312\
        );

    \I__10208\ : gio2CtrlBuf
    port map (
            O => \N__44312\,
            I => \delay_measurement_inst.delay_hc_timer.N_335_i_g\
        );

    \I__10207\ : InMux
    port map (
            O => \N__44309\,
            I => \N__44306\
        );

    \I__10206\ : LocalMux
    port map (
            O => \N__44306\,
            I => \N__44302\
        );

    \I__10205\ : InMux
    port map (
            O => \N__44305\,
            I => \N__44299\
        );

    \I__10204\ : Span4Mux_v
    port map (
            O => \N__44302\,
            I => \N__44293\
        );

    \I__10203\ : LocalMux
    port map (
            O => \N__44299\,
            I => \N__44293\
        );

    \I__10202\ : InMux
    port map (
            O => \N__44298\,
            I => \N__44290\
        );

    \I__10201\ : Odrv4
    port map (
            O => \N__44293\,
            I => \delay_measurement_inst.elapsed_time_hc_18\
        );

    \I__10200\ : LocalMux
    port map (
            O => \N__44290\,
            I => \delay_measurement_inst.elapsed_time_hc_18\
        );

    \I__10199\ : InMux
    port map (
            O => \N__44285\,
            I => \N__44281\
        );

    \I__10198\ : InMux
    port map (
            O => \N__44284\,
            I => \N__44278\
        );

    \I__10197\ : LocalMux
    port map (
            O => \N__44281\,
            I => \N__44274\
        );

    \I__10196\ : LocalMux
    port map (
            O => \N__44278\,
            I => \N__44271\
        );

    \I__10195\ : InMux
    port map (
            O => \N__44277\,
            I => \N__44268\
        );

    \I__10194\ : Odrv12
    port map (
            O => \N__44274\,
            I => \delay_measurement_inst.elapsed_time_hc_17\
        );

    \I__10193\ : Odrv4
    port map (
            O => \N__44271\,
            I => \delay_measurement_inst.elapsed_time_hc_17\
        );

    \I__10192\ : LocalMux
    port map (
            O => \N__44268\,
            I => \delay_measurement_inst.elapsed_time_hc_17\
        );

    \I__10191\ : CascadeMux
    port map (
            O => \N__44261\,
            I => \N__44258\
        );

    \I__10190\ : InMux
    port map (
            O => \N__44258\,
            I => \N__44254\
        );

    \I__10189\ : InMux
    port map (
            O => \N__44257\,
            I => \N__44251\
        );

    \I__10188\ : LocalMux
    port map (
            O => \N__44254\,
            I => \N__44247\
        );

    \I__10187\ : LocalMux
    port map (
            O => \N__44251\,
            I => \N__44244\
        );

    \I__10186\ : CascadeMux
    port map (
            O => \N__44250\,
            I => \N__44241\
        );

    \I__10185\ : Span4Mux_v
    port map (
            O => \N__44247\,
            I => \N__44236\
        );

    \I__10184\ : Span4Mux_v
    port map (
            O => \N__44244\,
            I => \N__44236\
        );

    \I__10183\ : InMux
    port map (
            O => \N__44241\,
            I => \N__44233\
        );

    \I__10182\ : Odrv4
    port map (
            O => \N__44236\,
            I => \delay_measurement_inst.elapsed_time_hc_19\
        );

    \I__10181\ : LocalMux
    port map (
            O => \N__44233\,
            I => \delay_measurement_inst.elapsed_time_hc_19\
        );

    \I__10180\ : InMux
    port map (
            O => \N__44228\,
            I => \N__44224\
        );

    \I__10179\ : InMux
    port map (
            O => \N__44227\,
            I => \N__44221\
        );

    \I__10178\ : LocalMux
    port map (
            O => \N__44224\,
            I => \N__44217\
        );

    \I__10177\ : LocalMux
    port map (
            O => \N__44221\,
            I => \N__44214\
        );

    \I__10176\ : InMux
    port map (
            O => \N__44220\,
            I => \N__44211\
        );

    \I__10175\ : Odrv12
    port map (
            O => \N__44217\,
            I => \delay_measurement_inst.elapsed_time_hc_16\
        );

    \I__10174\ : Odrv4
    port map (
            O => \N__44214\,
            I => \delay_measurement_inst.elapsed_time_hc_16\
        );

    \I__10173\ : LocalMux
    port map (
            O => \N__44211\,
            I => \delay_measurement_inst.elapsed_time_hc_16\
        );

    \I__10172\ : InMux
    port map (
            O => \N__44204\,
            I => \N__44201\
        );

    \I__10171\ : LocalMux
    port map (
            O => \N__44201\,
            I => \N__44197\
        );

    \I__10170\ : InMux
    port map (
            O => \N__44200\,
            I => \N__44194\
        );

    \I__10169\ : Span4Mux_v
    port map (
            O => \N__44197\,
            I => \N__44189\
        );

    \I__10168\ : LocalMux
    port map (
            O => \N__44194\,
            I => \N__44189\
        );

    \I__10167\ : Span4Mux_v
    port map (
            O => \N__44189\,
            I => \N__44186\
        );

    \I__10166\ : Sp12to4
    port map (
            O => \N__44186\,
            I => \N__44178\
        );

    \I__10165\ : InMux
    port map (
            O => \N__44185\,
            I => \N__44175\
        );

    \I__10164\ : InMux
    port map (
            O => \N__44184\,
            I => \N__44168\
        );

    \I__10163\ : InMux
    port map (
            O => \N__44183\,
            I => \N__44168\
        );

    \I__10162\ : InMux
    port map (
            O => \N__44182\,
            I => \N__44168\
        );

    \I__10161\ : InMux
    port map (
            O => \N__44181\,
            I => \N__44165\
        );

    \I__10160\ : Odrv12
    port map (
            O => \N__44178\,
            I => \delay_measurement_inst.elapsed_time_hc_31\
        );

    \I__10159\ : LocalMux
    port map (
            O => \N__44175\,
            I => \delay_measurement_inst.elapsed_time_hc_31\
        );

    \I__10158\ : LocalMux
    port map (
            O => \N__44168\,
            I => \delay_measurement_inst.elapsed_time_hc_31\
        );

    \I__10157\ : LocalMux
    port map (
            O => \N__44165\,
            I => \delay_measurement_inst.elapsed_time_hc_31\
        );

    \I__10156\ : InMux
    port map (
            O => \N__44156\,
            I => \N__44153\
        );

    \I__10155\ : LocalMux
    port map (
            O => \N__44153\,
            I => \N__44150\
        );

    \I__10154\ : Span4Mux_h
    port map (
            O => \N__44150\,
            I => \N__44146\
        );

    \I__10153\ : InMux
    port map (
            O => \N__44149\,
            I => \N__44142\
        );

    \I__10152\ : Span4Mux_h
    port map (
            O => \N__44146\,
            I => \N__44139\
        );

    \I__10151\ : InMux
    port map (
            O => \N__44145\,
            I => \N__44135\
        );

    \I__10150\ : LocalMux
    port map (
            O => \N__44142\,
            I => \N__44130\
        );

    \I__10149\ : Span4Mux_v
    port map (
            O => \N__44139\,
            I => \N__44127\
        );

    \I__10148\ : InMux
    port map (
            O => \N__44138\,
            I => \N__44124\
        );

    \I__10147\ : LocalMux
    port map (
            O => \N__44135\,
            I => \N__44121\
        );

    \I__10146\ : InMux
    port map (
            O => \N__44134\,
            I => \N__44118\
        );

    \I__10145\ : InMux
    port map (
            O => \N__44133\,
            I => \N__44115\
        );

    \I__10144\ : Span4Mux_h
    port map (
            O => \N__44130\,
            I => \N__44112\
        );

    \I__10143\ : Span4Mux_v
    port map (
            O => \N__44127\,
            I => \N__44107\
        );

    \I__10142\ : LocalMux
    port map (
            O => \N__44124\,
            I => \N__44107\
        );

    \I__10141\ : Span4Mux_v
    port map (
            O => \N__44121\,
            I => \N__44102\
        );

    \I__10140\ : LocalMux
    port map (
            O => \N__44118\,
            I => \N__44102\
        );

    \I__10139\ : LocalMux
    port map (
            O => \N__44115\,
            I => \N__44099\
        );

    \I__10138\ : Odrv4
    port map (
            O => \N__44112\,
            I => \delay_measurement_inst.delay_hc_reg3lto14\
        );

    \I__10137\ : Odrv4
    port map (
            O => \N__44107\,
            I => \delay_measurement_inst.delay_hc_reg3lto14\
        );

    \I__10136\ : Odrv4
    port map (
            O => \N__44102\,
            I => \delay_measurement_inst.delay_hc_reg3lto14\
        );

    \I__10135\ : Odrv4
    port map (
            O => \N__44099\,
            I => \delay_measurement_inst.delay_hc_reg3lto14\
        );

    \I__10134\ : InMux
    port map (
            O => \N__44090\,
            I => \N__44087\
        );

    \I__10133\ : LocalMux
    port map (
            O => \N__44087\,
            I => \N__44084\
        );

    \I__10132\ : Odrv4
    port map (
            O => \N__44084\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_a0_1\
        );

    \I__10131\ : InMux
    port map (
            O => \N__44081\,
            I => \N__44075\
        );

    \I__10130\ : InMux
    port map (
            O => \N__44080\,
            I => \N__44072\
        );

    \I__10129\ : InMux
    port map (
            O => \N__44079\,
            I => \N__44068\
        );

    \I__10128\ : InMux
    port map (
            O => \N__44078\,
            I => \N__44064\
        );

    \I__10127\ : LocalMux
    port map (
            O => \N__44075\,
            I => \N__44061\
        );

    \I__10126\ : LocalMux
    port map (
            O => \N__44072\,
            I => \N__44058\
        );

    \I__10125\ : InMux
    port map (
            O => \N__44071\,
            I => \N__44055\
        );

    \I__10124\ : LocalMux
    port map (
            O => \N__44068\,
            I => \N__44052\
        );

    \I__10123\ : InMux
    port map (
            O => \N__44067\,
            I => \N__44049\
        );

    \I__10122\ : LocalMux
    port map (
            O => \N__44064\,
            I => \N__44046\
        );

    \I__10121\ : Span4Mux_h
    port map (
            O => \N__44061\,
            I => \N__44043\
        );

    \I__10120\ : Span4Mux_h
    port map (
            O => \N__44058\,
            I => \N__44040\
        );

    \I__10119\ : LocalMux
    port map (
            O => \N__44055\,
            I => \N__44037\
        );

    \I__10118\ : Span4Mux_h
    port map (
            O => \N__44052\,
            I => \N__44032\
        );

    \I__10117\ : LocalMux
    port map (
            O => \N__44049\,
            I => \N__44032\
        );

    \I__10116\ : Odrv4
    port map (
            O => \N__44046\,
            I => \delay_measurement_inst.delay_hc_reg3lto9\
        );

    \I__10115\ : Odrv4
    port map (
            O => \N__44043\,
            I => \delay_measurement_inst.delay_hc_reg3lto9\
        );

    \I__10114\ : Odrv4
    port map (
            O => \N__44040\,
            I => \delay_measurement_inst.delay_hc_reg3lto9\
        );

    \I__10113\ : Odrv4
    port map (
            O => \N__44037\,
            I => \delay_measurement_inst.delay_hc_reg3lto9\
        );

    \I__10112\ : Odrv4
    port map (
            O => \N__44032\,
            I => \delay_measurement_inst.delay_hc_reg3lto9\
        );

    \I__10111\ : CascadeMux
    port map (
            O => \N__44021\,
            I => \N__44017\
        );

    \I__10110\ : InMux
    port map (
            O => \N__44020\,
            I => \N__44010\
        );

    \I__10109\ : InMux
    port map (
            O => \N__44017\,
            I => \N__44007\
        );

    \I__10108\ : InMux
    port map (
            O => \N__44016\,
            I => \N__44000\
        );

    \I__10107\ : InMux
    port map (
            O => \N__44015\,
            I => \N__44000\
        );

    \I__10106\ : InMux
    port map (
            O => \N__44014\,
            I => \N__44000\
        );

    \I__10105\ : InMux
    port map (
            O => \N__44013\,
            I => \N__43997\
        );

    \I__10104\ : LocalMux
    port map (
            O => \N__44010\,
            I => \N__43994\
        );

    \I__10103\ : LocalMux
    port map (
            O => \N__44007\,
            I => \N__43991\
        );

    \I__10102\ : LocalMux
    port map (
            O => \N__44000\,
            I => \N__43988\
        );

    \I__10101\ : LocalMux
    port map (
            O => \N__43997\,
            I => \N__43985\
        );

    \I__10100\ : Span4Mux_h
    port map (
            O => \N__43994\,
            I => \N__43982\
        );

    \I__10099\ : Span4Mux_h
    port map (
            O => \N__43991\,
            I => \N__43977\
        );

    \I__10098\ : Span4Mux_h
    port map (
            O => \N__43988\,
            I => \N__43977\
        );

    \I__10097\ : Odrv4
    port map (
            O => \N__43985\,
            I => \delay_measurement_inst.delay_hc_reg3lto6\
        );

    \I__10096\ : Odrv4
    port map (
            O => \N__43982\,
            I => \delay_measurement_inst.delay_hc_reg3lto6\
        );

    \I__10095\ : Odrv4
    port map (
            O => \N__43977\,
            I => \delay_measurement_inst.delay_hc_reg3lto6\
        );

    \I__10094\ : CascadeMux
    port map (
            O => \N__43970\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_a0_1_cascade_\
        );

    \I__10093\ : InMux
    port map (
            O => \N__43967\,
            I => \N__43964\
        );

    \I__10092\ : LocalMux
    port map (
            O => \N__43964\,
            I => \N__43960\
        );

    \I__10091\ : InMux
    port map (
            O => \N__43963\,
            I => \N__43957\
        );

    \I__10090\ : Span4Mux_v
    port map (
            O => \N__43960\,
            I => \N__43951\
        );

    \I__10089\ : LocalMux
    port map (
            O => \N__43957\,
            I => \N__43951\
        );

    \I__10088\ : InMux
    port map (
            O => \N__43956\,
            I => \N__43947\
        );

    \I__10087\ : Span4Mux_v
    port map (
            O => \N__43951\,
            I => \N__43944\
        );

    \I__10086\ : InMux
    port map (
            O => \N__43950\,
            I => \N__43940\
        );

    \I__10085\ : LocalMux
    port map (
            O => \N__43947\,
            I => \N__43935\
        );

    \I__10084\ : Span4Mux_h
    port map (
            O => \N__43944\,
            I => \N__43935\
        );

    \I__10083\ : InMux
    port map (
            O => \N__43943\,
            I => \N__43932\
        );

    \I__10082\ : LocalMux
    port map (
            O => \N__43940\,
            I => \N__43929\
        );

    \I__10081\ : Span4Mux_h
    port map (
            O => \N__43935\,
            I => \N__43925\
        );

    \I__10080\ : LocalMux
    port map (
            O => \N__43932\,
            I => \N__43922\
        );

    \I__10079\ : Span4Mux_h
    port map (
            O => \N__43929\,
            I => \N__43919\
        );

    \I__10078\ : InMux
    port map (
            O => \N__43928\,
            I => \N__43916\
        );

    \I__10077\ : Odrv4
    port map (
            O => \N__43925\,
            I => \delay_measurement_inst.delay_hc_reg3lto19_1\
        );

    \I__10076\ : Odrv4
    port map (
            O => \N__43922\,
            I => \delay_measurement_inst.delay_hc_reg3lto19_1\
        );

    \I__10075\ : Odrv4
    port map (
            O => \N__43919\,
            I => \delay_measurement_inst.delay_hc_reg3lto19_1\
        );

    \I__10074\ : LocalMux
    port map (
            O => \N__43916\,
            I => \delay_measurement_inst.delay_hc_reg3lto19_1\
        );

    \I__10073\ : InMux
    port map (
            O => \N__43907\,
            I => \N__43904\
        );

    \I__10072\ : LocalMux
    port map (
            O => \N__43904\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_a0_2\
        );

    \I__10071\ : InMux
    port map (
            O => \N__43901\,
            I => \N__43897\
        );

    \I__10070\ : InMux
    port map (
            O => \N__43900\,
            I => \N__43893\
        );

    \I__10069\ : LocalMux
    port map (
            O => \N__43897\,
            I => \N__43890\
        );

    \I__10068\ : InMux
    port map (
            O => \N__43896\,
            I => \N__43887\
        );

    \I__10067\ : LocalMux
    port map (
            O => \N__43893\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__10066\ : Odrv4
    port map (
            O => \N__43890\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__10065\ : LocalMux
    port map (
            O => \N__43887\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__10064\ : InMux
    port map (
            O => \N__43880\,
            I => \N__43876\
        );

    \I__10063\ : InMux
    port map (
            O => \N__43879\,
            I => \N__43872\
        );

    \I__10062\ : LocalMux
    port map (
            O => \N__43876\,
            I => \N__43869\
        );

    \I__10061\ : InMux
    port map (
            O => \N__43875\,
            I => \N__43866\
        );

    \I__10060\ : LocalMux
    port map (
            O => \N__43872\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__10059\ : Odrv4
    port map (
            O => \N__43869\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__10058\ : LocalMux
    port map (
            O => \N__43866\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__10057\ : InMux
    port map (
            O => \N__43859\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__10056\ : CascadeMux
    port map (
            O => \N__43856\,
            I => \N__43849\
        );

    \I__10055\ : CascadeMux
    port map (
            O => \N__43855\,
            I => \N__43846\
        );

    \I__10054\ : InMux
    port map (
            O => \N__43854\,
            I => \N__43836\
        );

    \I__10053\ : InMux
    port map (
            O => \N__43853\,
            I => \N__43830\
        );

    \I__10052\ : InMux
    port map (
            O => \N__43852\,
            I => \N__43819\
        );

    \I__10051\ : InMux
    port map (
            O => \N__43849\,
            I => \N__43816\
        );

    \I__10050\ : InMux
    port map (
            O => \N__43846\,
            I => \N__43799\
        );

    \I__10049\ : InMux
    port map (
            O => \N__43845\,
            I => \N__43799\
        );

    \I__10048\ : InMux
    port map (
            O => \N__43844\,
            I => \N__43799\
        );

    \I__10047\ : InMux
    port map (
            O => \N__43843\,
            I => \N__43799\
        );

    \I__10046\ : InMux
    port map (
            O => \N__43842\,
            I => \N__43799\
        );

    \I__10045\ : InMux
    port map (
            O => \N__43841\,
            I => \N__43799\
        );

    \I__10044\ : InMux
    port map (
            O => \N__43840\,
            I => \N__43799\
        );

    \I__10043\ : InMux
    port map (
            O => \N__43839\,
            I => \N__43799\
        );

    \I__10042\ : LocalMux
    port map (
            O => \N__43836\,
            I => \N__43796\
        );

    \I__10041\ : InMux
    port map (
            O => \N__43835\,
            I => \N__43791\
        );

    \I__10040\ : InMux
    port map (
            O => \N__43834\,
            I => \N__43791\
        );

    \I__10039\ : CascadeMux
    port map (
            O => \N__43833\,
            I => \N__43787\
        );

    \I__10038\ : LocalMux
    port map (
            O => \N__43830\,
            I => \N__43784\
        );

    \I__10037\ : InMux
    port map (
            O => \N__43829\,
            I => \N__43767\
        );

    \I__10036\ : InMux
    port map (
            O => \N__43828\,
            I => \N__43767\
        );

    \I__10035\ : InMux
    port map (
            O => \N__43827\,
            I => \N__43767\
        );

    \I__10034\ : InMux
    port map (
            O => \N__43826\,
            I => \N__43767\
        );

    \I__10033\ : InMux
    port map (
            O => \N__43825\,
            I => \N__43767\
        );

    \I__10032\ : InMux
    port map (
            O => \N__43824\,
            I => \N__43767\
        );

    \I__10031\ : InMux
    port map (
            O => \N__43823\,
            I => \N__43767\
        );

    \I__10030\ : InMux
    port map (
            O => \N__43822\,
            I => \N__43767\
        );

    \I__10029\ : LocalMux
    port map (
            O => \N__43819\,
            I => \N__43764\
        );

    \I__10028\ : LocalMux
    port map (
            O => \N__43816\,
            I => \N__43755\
        );

    \I__10027\ : LocalMux
    port map (
            O => \N__43799\,
            I => \N__43755\
        );

    \I__10026\ : Span4Mux_v
    port map (
            O => \N__43796\,
            I => \N__43755\
        );

    \I__10025\ : LocalMux
    port map (
            O => \N__43791\,
            I => \N__43755\
        );

    \I__10024\ : InMux
    port map (
            O => \N__43790\,
            I => \N__43750\
        );

    \I__10023\ : InMux
    port map (
            O => \N__43787\,
            I => \N__43750\
        );

    \I__10022\ : Span4Mux_v
    port map (
            O => \N__43784\,
            I => \N__43747\
        );

    \I__10021\ : LocalMux
    port map (
            O => \N__43767\,
            I => \N__43740\
        );

    \I__10020\ : Span4Mux_v
    port map (
            O => \N__43764\,
            I => \N__43740\
        );

    \I__10019\ : Span4Mux_v
    port map (
            O => \N__43755\,
            I => \N__43740\
        );

    \I__10018\ : LocalMux
    port map (
            O => \N__43750\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__10017\ : Odrv4
    port map (
            O => \N__43747\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__10016\ : Odrv4
    port map (
            O => \N__43740\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__10015\ : CascadeMux
    port map (
            O => \N__43733\,
            I => \N__43729\
        );

    \I__10014\ : CascadeMux
    port map (
            O => \N__43732\,
            I => \N__43725\
        );

    \I__10013\ : InMux
    port map (
            O => \N__43729\,
            I => \N__43715\
        );

    \I__10012\ : InMux
    port map (
            O => \N__43728\,
            I => \N__43715\
        );

    \I__10011\ : InMux
    port map (
            O => \N__43725\,
            I => \N__43707\
        );

    \I__10010\ : CascadeMux
    port map (
            O => \N__43724\,
            I => \N__43704\
        );

    \I__10009\ : CascadeMux
    port map (
            O => \N__43723\,
            I => \N__43697\
        );

    \I__10008\ : CascadeMux
    port map (
            O => \N__43722\,
            I => \N__43694\
        );

    \I__10007\ : CascadeMux
    port map (
            O => \N__43721\,
            I => \N__43691\
        );

    \I__10006\ : CascadeMux
    port map (
            O => \N__43720\,
            I => \N__43688\
        );

    \I__10005\ : LocalMux
    port map (
            O => \N__43715\,
            I => \N__43685\
        );

    \I__10004\ : InMux
    port map (
            O => \N__43714\,
            I => \N__43682\
        );

    \I__10003\ : CascadeMux
    port map (
            O => \N__43713\,
            I => \N__43678\
        );

    \I__10002\ : CascadeMux
    port map (
            O => \N__43712\,
            I => \N__43675\
        );

    \I__10001\ : CascadeMux
    port map (
            O => \N__43711\,
            I => \N__43672\
        );

    \I__10000\ : CascadeMux
    port map (
            O => \N__43710\,
            I => \N__43669\
        );

    \I__9999\ : LocalMux
    port map (
            O => \N__43707\,
            I => \N__43661\
        );

    \I__9998\ : InMux
    port map (
            O => \N__43704\,
            I => \N__43657\
        );

    \I__9997\ : InMux
    port map (
            O => \N__43703\,
            I => \N__43640\
        );

    \I__9996\ : InMux
    port map (
            O => \N__43702\,
            I => \N__43640\
        );

    \I__9995\ : InMux
    port map (
            O => \N__43701\,
            I => \N__43640\
        );

    \I__9994\ : InMux
    port map (
            O => \N__43700\,
            I => \N__43640\
        );

    \I__9993\ : InMux
    port map (
            O => \N__43697\,
            I => \N__43640\
        );

    \I__9992\ : InMux
    port map (
            O => \N__43694\,
            I => \N__43640\
        );

    \I__9991\ : InMux
    port map (
            O => \N__43691\,
            I => \N__43640\
        );

    \I__9990\ : InMux
    port map (
            O => \N__43688\,
            I => \N__43640\
        );

    \I__9989\ : Span4Mux_v
    port map (
            O => \N__43685\,
            I => \N__43635\
        );

    \I__9988\ : LocalMux
    port map (
            O => \N__43682\,
            I => \N__43635\
        );

    \I__9987\ : InMux
    port map (
            O => \N__43681\,
            I => \N__43618\
        );

    \I__9986\ : InMux
    port map (
            O => \N__43678\,
            I => \N__43618\
        );

    \I__9985\ : InMux
    port map (
            O => \N__43675\,
            I => \N__43618\
        );

    \I__9984\ : InMux
    port map (
            O => \N__43672\,
            I => \N__43618\
        );

    \I__9983\ : InMux
    port map (
            O => \N__43669\,
            I => \N__43618\
        );

    \I__9982\ : InMux
    port map (
            O => \N__43668\,
            I => \N__43618\
        );

    \I__9981\ : InMux
    port map (
            O => \N__43667\,
            I => \N__43618\
        );

    \I__9980\ : InMux
    port map (
            O => \N__43666\,
            I => \N__43618\
        );

    \I__9979\ : InMux
    port map (
            O => \N__43665\,
            I => \N__43613\
        );

    \I__9978\ : InMux
    port map (
            O => \N__43664\,
            I => \N__43613\
        );

    \I__9977\ : Span4Mux_v
    port map (
            O => \N__43661\,
            I => \N__43610\
        );

    \I__9976\ : InMux
    port map (
            O => \N__43660\,
            I => \N__43607\
        );

    \I__9975\ : LocalMux
    port map (
            O => \N__43657\,
            I => \N__43600\
        );

    \I__9974\ : LocalMux
    port map (
            O => \N__43640\,
            I => \N__43600\
        );

    \I__9973\ : Span4Mux_h
    port map (
            O => \N__43635\,
            I => \N__43600\
        );

    \I__9972\ : LocalMux
    port map (
            O => \N__43618\,
            I => \phase_controller_slave.start_timer_hcZ0\
        );

    \I__9971\ : LocalMux
    port map (
            O => \N__43613\,
            I => \phase_controller_slave.start_timer_hcZ0\
        );

    \I__9970\ : Odrv4
    port map (
            O => \N__43610\,
            I => \phase_controller_slave.start_timer_hcZ0\
        );

    \I__9969\ : LocalMux
    port map (
            O => \N__43607\,
            I => \phase_controller_slave.start_timer_hcZ0\
        );

    \I__9968\ : Odrv4
    port map (
            O => \N__43600\,
            I => \phase_controller_slave.start_timer_hcZ0\
        );

    \I__9967\ : CascadeMux
    port map (
            O => \N__43589\,
            I => \N__43580\
        );

    \I__9966\ : CascadeMux
    port map (
            O => \N__43588\,
            I => \N__43577\
        );

    \I__9965\ : CascadeMux
    port map (
            O => \N__43587\,
            I => \N__43574\
        );

    \I__9964\ : CascadeMux
    port map (
            O => \N__43586\,
            I => \N__43565\
        );

    \I__9963\ : InMux
    port map (
            O => \N__43585\,
            I => \N__43561\
        );

    \I__9962\ : InMux
    port map (
            O => \N__43584\,
            I => \N__43550\
        );

    \I__9961\ : InMux
    port map (
            O => \N__43583\,
            I => \N__43547\
        );

    \I__9960\ : InMux
    port map (
            O => \N__43580\,
            I => \N__43540\
        );

    \I__9959\ : InMux
    port map (
            O => \N__43577\,
            I => \N__43540\
        );

    \I__9958\ : InMux
    port map (
            O => \N__43574\,
            I => \N__43540\
        );

    \I__9957\ : InMux
    port map (
            O => \N__43573\,
            I => \N__43529\
        );

    \I__9956\ : InMux
    port map (
            O => \N__43572\,
            I => \N__43529\
        );

    \I__9955\ : InMux
    port map (
            O => \N__43571\,
            I => \N__43529\
        );

    \I__9954\ : InMux
    port map (
            O => \N__43570\,
            I => \N__43529\
        );

    \I__9953\ : InMux
    port map (
            O => \N__43569\,
            I => \N__43529\
        );

    \I__9952\ : InMux
    port map (
            O => \N__43568\,
            I => \N__43526\
        );

    \I__9951\ : InMux
    port map (
            O => \N__43565\,
            I => \N__43521\
        );

    \I__9950\ : InMux
    port map (
            O => \N__43564\,
            I => \N__43521\
        );

    \I__9949\ : LocalMux
    port map (
            O => \N__43561\,
            I => \N__43516\
        );

    \I__9948\ : InMux
    port map (
            O => \N__43560\,
            I => \N__43499\
        );

    \I__9947\ : InMux
    port map (
            O => \N__43559\,
            I => \N__43499\
        );

    \I__9946\ : InMux
    port map (
            O => \N__43558\,
            I => \N__43499\
        );

    \I__9945\ : InMux
    port map (
            O => \N__43557\,
            I => \N__43499\
        );

    \I__9944\ : InMux
    port map (
            O => \N__43556\,
            I => \N__43499\
        );

    \I__9943\ : InMux
    port map (
            O => \N__43555\,
            I => \N__43499\
        );

    \I__9942\ : InMux
    port map (
            O => \N__43554\,
            I => \N__43499\
        );

    \I__9941\ : InMux
    port map (
            O => \N__43553\,
            I => \N__43499\
        );

    \I__9940\ : LocalMux
    port map (
            O => \N__43550\,
            I => \N__43494\
        );

    \I__9939\ : LocalMux
    port map (
            O => \N__43547\,
            I => \N__43494\
        );

    \I__9938\ : LocalMux
    port map (
            O => \N__43540\,
            I => \N__43485\
        );

    \I__9937\ : LocalMux
    port map (
            O => \N__43529\,
            I => \N__43485\
        );

    \I__9936\ : LocalMux
    port map (
            O => \N__43526\,
            I => \N__43485\
        );

    \I__9935\ : LocalMux
    port map (
            O => \N__43521\,
            I => \N__43485\
        );

    \I__9934\ : InMux
    port map (
            O => \N__43520\,
            I => \N__43480\
        );

    \I__9933\ : InMux
    port map (
            O => \N__43519\,
            I => \N__43480\
        );

    \I__9932\ : Span4Mux_v
    port map (
            O => \N__43516\,
            I => \N__43477\
        );

    \I__9931\ : LocalMux
    port map (
            O => \N__43499\,
            I => \N__43470\
        );

    \I__9930\ : Span4Mux_v
    port map (
            O => \N__43494\,
            I => \N__43470\
        );

    \I__9929\ : Span4Mux_v
    port map (
            O => \N__43485\,
            I => \N__43470\
        );

    \I__9928\ : LocalMux
    port map (
            O => \N__43480\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__9927\ : Odrv4
    port map (
            O => \N__43477\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__9926\ : Odrv4
    port map (
            O => \N__43470\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__9925\ : CascadeMux
    port map (
            O => \N__43463\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4Z0Z_3_cascade_\
        );

    \I__9924\ : CascadeMux
    port map (
            O => \N__43460\,
            I => \N__43457\
        );

    \I__9923\ : InMux
    port map (
            O => \N__43457\,
            I => \N__43453\
        );

    \I__9922\ : InMux
    port map (
            O => \N__43456\,
            I => \N__43450\
        );

    \I__9921\ : LocalMux
    port map (
            O => \N__43453\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9\
        );

    \I__9920\ : LocalMux
    port map (
            O => \N__43450\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9\
        );

    \I__9919\ : InMux
    port map (
            O => \N__43445\,
            I => \N__43442\
        );

    \I__9918\ : LocalMux
    port map (
            O => \N__43442\,
            I => \N__43431\
        );

    \I__9917\ : InMux
    port map (
            O => \N__43441\,
            I => \N__43424\
        );

    \I__9916\ : InMux
    port map (
            O => \N__43440\,
            I => \N__43424\
        );

    \I__9915\ : InMux
    port map (
            O => \N__43439\,
            I => \N__43424\
        );

    \I__9914\ : InMux
    port map (
            O => \N__43438\,
            I => \N__43413\
        );

    \I__9913\ : InMux
    port map (
            O => \N__43437\,
            I => \N__43413\
        );

    \I__9912\ : InMux
    port map (
            O => \N__43436\,
            I => \N__43413\
        );

    \I__9911\ : InMux
    port map (
            O => \N__43435\,
            I => \N__43413\
        );

    \I__9910\ : InMux
    port map (
            O => \N__43434\,
            I => \N__43413\
        );

    \I__9909\ : Span4Mux_h
    port map (
            O => \N__43431\,
            I => \N__43403\
        );

    \I__9908\ : LocalMux
    port map (
            O => \N__43424\,
            I => \N__43400\
        );

    \I__9907\ : LocalMux
    port map (
            O => \N__43413\,
            I => \N__43397\
        );

    \I__9906\ : InMux
    port map (
            O => \N__43412\,
            I => \N__43382\
        );

    \I__9905\ : InMux
    port map (
            O => \N__43411\,
            I => \N__43382\
        );

    \I__9904\ : InMux
    port map (
            O => \N__43410\,
            I => \N__43382\
        );

    \I__9903\ : InMux
    port map (
            O => \N__43409\,
            I => \N__43382\
        );

    \I__9902\ : InMux
    port map (
            O => \N__43408\,
            I => \N__43382\
        );

    \I__9901\ : InMux
    port map (
            O => \N__43407\,
            I => \N__43382\
        );

    \I__9900\ : InMux
    port map (
            O => \N__43406\,
            I => \N__43382\
        );

    \I__9899\ : Odrv4
    port map (
            O => \N__43403\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6\
        );

    \I__9898\ : Odrv4
    port map (
            O => \N__43400\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6\
        );

    \I__9897\ : Odrv4
    port map (
            O => \N__43397\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6\
        );

    \I__9896\ : LocalMux
    port map (
            O => \N__43382\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6\
        );

    \I__9895\ : CascadeMux
    port map (
            O => \N__43373\,
            I => \N__43370\
        );

    \I__9894\ : InMux
    port map (
            O => \N__43370\,
            I => \N__43367\
        );

    \I__9893\ : LocalMux
    port map (
            O => \N__43367\,
            I => \N__43364\
        );

    \I__9892\ : Span4Mux_h
    port map (
            O => \N__43364\,
            I => \N__43361\
        );

    \I__9891\ : Odrv4
    port map (
            O => \N__43361\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_14\
        );

    \I__9890\ : CEMux
    port map (
            O => \N__43358\,
            I => \N__43355\
        );

    \I__9889\ : LocalMux
    port map (
            O => \N__43355\,
            I => \N__43349\
        );

    \I__9888\ : CEMux
    port map (
            O => \N__43354\,
            I => \N__43345\
        );

    \I__9887\ : CEMux
    port map (
            O => \N__43353\,
            I => \N__43342\
        );

    \I__9886\ : CEMux
    port map (
            O => \N__43352\,
            I => \N__43339\
        );

    \I__9885\ : Span4Mux_h
    port map (
            O => \N__43349\,
            I => \N__43336\
        );

    \I__9884\ : CEMux
    port map (
            O => \N__43348\,
            I => \N__43333\
        );

    \I__9883\ : LocalMux
    port map (
            O => \N__43345\,
            I => \N__43330\
        );

    \I__9882\ : LocalMux
    port map (
            O => \N__43342\,
            I => \N__43325\
        );

    \I__9881\ : LocalMux
    port map (
            O => \N__43339\,
            I => \N__43325\
        );

    \I__9880\ : Span4Mux_v
    port map (
            O => \N__43336\,
            I => \N__43318\
        );

    \I__9879\ : LocalMux
    port map (
            O => \N__43333\,
            I => \N__43318\
        );

    \I__9878\ : Span4Mux_h
    port map (
            O => \N__43330\,
            I => \N__43318\
        );

    \I__9877\ : Span4Mux_v
    port map (
            O => \N__43325\,
            I => \N__43315\
        );

    \I__9876\ : Odrv4
    port map (
            O => \N__43318\,
            I => \phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__9875\ : Odrv4
    port map (
            O => \N__43315\,
            I => \phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__9874\ : InMux
    port map (
            O => \N__43310\,
            I => \N__43304\
        );

    \I__9873\ : InMux
    port map (
            O => \N__43309\,
            I => \N__43304\
        );

    \I__9872\ : LocalMux
    port map (
            O => \N__43304\,
            I => \N__43293\
        );

    \I__9871\ : InMux
    port map (
            O => \N__43303\,
            I => \N__43290\
        );

    \I__9870\ : InMux
    port map (
            O => \N__43302\,
            I => \N__43281\
        );

    \I__9869\ : InMux
    port map (
            O => \N__43301\,
            I => \N__43281\
        );

    \I__9868\ : InMux
    port map (
            O => \N__43300\,
            I => \N__43281\
        );

    \I__9867\ : InMux
    port map (
            O => \N__43299\,
            I => \N__43281\
        );

    \I__9866\ : InMux
    port map (
            O => \N__43298\,
            I => \N__43274\
        );

    \I__9865\ : InMux
    port map (
            O => \N__43297\,
            I => \N__43274\
        );

    \I__9864\ : InMux
    port map (
            O => \N__43296\,
            I => \N__43274\
        );

    \I__9863\ : Odrv4
    port map (
            O => \N__43293\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9\
        );

    \I__9862\ : LocalMux
    port map (
            O => \N__43290\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9\
        );

    \I__9861\ : LocalMux
    port map (
            O => \N__43281\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9\
        );

    \I__9860\ : LocalMux
    port map (
            O => \N__43274\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9\
        );

    \I__9859\ : InMux
    port map (
            O => \N__43265\,
            I => \N__43260\
        );

    \I__9858\ : InMux
    port map (
            O => \N__43264\,
            I => \N__43257\
        );

    \I__9857\ : InMux
    port map (
            O => \N__43263\,
            I => \N__43254\
        );

    \I__9856\ : LocalMux
    port map (
            O => \N__43260\,
            I => \N__43249\
        );

    \I__9855\ : LocalMux
    port map (
            O => \N__43257\,
            I => \N__43249\
        );

    \I__9854\ : LocalMux
    port map (
            O => \N__43254\,
            I => \phase_controller_inst1.stoper_tr.N_279\
        );

    \I__9853\ : Odrv4
    port map (
            O => \N__43249\,
            I => \phase_controller_inst1.stoper_tr.N_279\
        );

    \I__9852\ : InMux
    port map (
            O => \N__43244\,
            I => \N__43238\
        );

    \I__9851\ : InMux
    port map (
            O => \N__43243\,
            I => \N__43238\
        );

    \I__9850\ : LocalMux
    port map (
            O => \N__43238\,
            I => \N__43233\
        );

    \I__9849\ : InMux
    port map (
            O => \N__43237\,
            I => \N__43228\
        );

    \I__9848\ : InMux
    port map (
            O => \N__43236\,
            I => \N__43228\
        );

    \I__9847\ : Odrv4
    port map (
            O => \N__43233\,
            I => \phase_controller_inst1.stoper_tr.N_262\
        );

    \I__9846\ : LocalMux
    port map (
            O => \N__43228\,
            I => \phase_controller_inst1.stoper_tr.N_262\
        );

    \I__9845\ : CascadeMux
    port map (
            O => \N__43223\,
            I => \N__43219\
        );

    \I__9844\ : InMux
    port map (
            O => \N__43222\,
            I => \N__43215\
        );

    \I__9843\ : InMux
    port map (
            O => \N__43219\,
            I => \N__43212\
        );

    \I__9842\ : InMux
    port map (
            O => \N__43218\,
            I => \N__43209\
        );

    \I__9841\ : LocalMux
    port map (
            O => \N__43215\,
            I => \N__43206\
        );

    \I__9840\ : LocalMux
    port map (
            O => \N__43212\,
            I => \N__43203\
        );

    \I__9839\ : LocalMux
    port map (
            O => \N__43209\,
            I => \N__43200\
        );

    \I__9838\ : Span4Mux_v
    port map (
            O => \N__43206\,
            I => \N__43197\
        );

    \I__9837\ : Odrv12
    port map (
            O => \N__43203\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6\
        );

    \I__9836\ : Odrv4
    port map (
            O => \N__43200\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6\
        );

    \I__9835\ : Odrv4
    port map (
            O => \N__43197\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6\
        );

    \I__9834\ : InMux
    port map (
            O => \N__43190\,
            I => \N__43176\
        );

    \I__9833\ : InMux
    port map (
            O => \N__43189\,
            I => \N__43176\
        );

    \I__9832\ : InMux
    port map (
            O => \N__43188\,
            I => \N__43176\
        );

    \I__9831\ : InMux
    port map (
            O => \N__43187\,
            I => \N__43176\
        );

    \I__9830\ : InMux
    port map (
            O => \N__43186\,
            I => \N__43171\
        );

    \I__9829\ : InMux
    port map (
            O => \N__43185\,
            I => \N__43171\
        );

    \I__9828\ : LocalMux
    port map (
            O => \N__43176\,
            I => \N__43166\
        );

    \I__9827\ : LocalMux
    port map (
            O => \N__43171\,
            I => \N__43166\
        );

    \I__9826\ : Span4Mux_h
    port map (
            O => \N__43166\,
            I => \N__43157\
        );

    \I__9825\ : InMux
    port map (
            O => \N__43165\,
            I => \N__43154\
        );

    \I__9824\ : InMux
    port map (
            O => \N__43164\,
            I => \N__43143\
        );

    \I__9823\ : InMux
    port map (
            O => \N__43163\,
            I => \N__43143\
        );

    \I__9822\ : InMux
    port map (
            O => \N__43162\,
            I => \N__43143\
        );

    \I__9821\ : InMux
    port map (
            O => \N__43161\,
            I => \N__43143\
        );

    \I__9820\ : InMux
    port map (
            O => \N__43160\,
            I => \N__43143\
        );

    \I__9819\ : Odrv4
    port map (
            O => \N__43157\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6\
        );

    \I__9818\ : LocalMux
    port map (
            O => \N__43154\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6\
        );

    \I__9817\ : LocalMux
    port map (
            O => \N__43143\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6\
        );

    \I__9816\ : InMux
    port map (
            O => \N__43136\,
            I => \N__43133\
        );

    \I__9815\ : LocalMux
    port map (
            O => \N__43133\,
            I => \N__43130\
        );

    \I__9814\ : Span4Mux_h
    port map (
            O => \N__43130\,
            I => \N__43127\
        );

    \I__9813\ : Odrv4
    port map (
            O => \N__43127\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\
        );

    \I__9812\ : CEMux
    port map (
            O => \N__43124\,
            I => \N__43120\
        );

    \I__9811\ : CEMux
    port map (
            O => \N__43123\,
            I => \N__43117\
        );

    \I__9810\ : LocalMux
    port map (
            O => \N__43120\,
            I => \N__43112\
        );

    \I__9809\ : LocalMux
    port map (
            O => \N__43117\,
            I => \N__43112\
        );

    \I__9808\ : Span4Mux_v
    port map (
            O => \N__43112\,
            I => \N__43107\
        );

    \I__9807\ : CEMux
    port map (
            O => \N__43111\,
            I => \N__43104\
        );

    \I__9806\ : CEMux
    port map (
            O => \N__43110\,
            I => \N__43100\
        );

    \I__9805\ : Span4Mux_h
    port map (
            O => \N__43107\,
            I => \N__43095\
        );

    \I__9804\ : LocalMux
    port map (
            O => \N__43104\,
            I => \N__43095\
        );

    \I__9803\ : CEMux
    port map (
            O => \N__43103\,
            I => \N__43091\
        );

    \I__9802\ : LocalMux
    port map (
            O => \N__43100\,
            I => \N__43088\
        );

    \I__9801\ : Span4Mux_v
    port map (
            O => \N__43095\,
            I => \N__43085\
        );

    \I__9800\ : CEMux
    port map (
            O => \N__43094\,
            I => \N__43082\
        );

    \I__9799\ : LocalMux
    port map (
            O => \N__43091\,
            I => \N__43079\
        );

    \I__9798\ : Span4Mux_h
    port map (
            O => \N__43088\,
            I => \N__43076\
        );

    \I__9797\ : Sp12to4
    port map (
            O => \N__43085\,
            I => \N__43071\
        );

    \I__9796\ : LocalMux
    port map (
            O => \N__43082\,
            I => \N__43071\
        );

    \I__9795\ : Odrv4
    port map (
            O => \N__43079\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__9794\ : Odrv4
    port map (
            O => \N__43076\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__9793\ : Odrv12
    port map (
            O => \N__43071\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__9792\ : InMux
    port map (
            O => \N__43064\,
            I => \N__43058\
        );

    \I__9791\ : InMux
    port map (
            O => \N__43063\,
            I => \N__43055\
        );

    \I__9790\ : InMux
    port map (
            O => \N__43062\,
            I => \N__43050\
        );

    \I__9789\ : InMux
    port map (
            O => \N__43061\,
            I => \N__43050\
        );

    \I__9788\ : LocalMux
    port map (
            O => \N__43058\,
            I => \phase_controller_slave.stoper_hc.time_passed11\
        );

    \I__9787\ : LocalMux
    port map (
            O => \N__43055\,
            I => \phase_controller_slave.stoper_hc.time_passed11\
        );

    \I__9786\ : LocalMux
    port map (
            O => \N__43050\,
            I => \phase_controller_slave.stoper_hc.time_passed11\
        );

    \I__9785\ : CascadeMux
    port map (
            O => \N__43043\,
            I => \N__43040\
        );

    \I__9784\ : InMux
    port map (
            O => \N__43040\,
            I => \N__43037\
        );

    \I__9783\ : LocalMux
    port map (
            O => \N__43037\,
            I => \phase_controller_slave.stoper_hc.time_passed_1_sqmuxa\
        );

    \I__9782\ : InMux
    port map (
            O => \N__43034\,
            I => \N__43029\
        );

    \I__9781\ : InMux
    port map (
            O => \N__43033\,
            I => \N__43024\
        );

    \I__9780\ : InMux
    port map (
            O => \N__43032\,
            I => \N__43024\
        );

    \I__9779\ : LocalMux
    port map (
            O => \N__43029\,
            I => \N__43019\
        );

    \I__9778\ : LocalMux
    port map (
            O => \N__43024\,
            I => \N__43016\
        );

    \I__9777\ : InMux
    port map (
            O => \N__43023\,
            I => \N__43010\
        );

    \I__9776\ : InMux
    port map (
            O => \N__43022\,
            I => \N__43010\
        );

    \I__9775\ : Span4Mux_v
    port map (
            O => \N__43019\,
            I => \N__43007\
        );

    \I__9774\ : Span4Mux_h
    port map (
            O => \N__43016\,
            I => \N__43004\
        );

    \I__9773\ : InMux
    port map (
            O => \N__43015\,
            I => \N__43001\
        );

    \I__9772\ : LocalMux
    port map (
            O => \N__43010\,
            I => \N__42998\
        );

    \I__9771\ : Odrv4
    port map (
            O => \N__43007\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__9770\ : Odrv4
    port map (
            O => \N__43004\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__9769\ : LocalMux
    port map (
            O => \N__43001\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__9768\ : Odrv4
    port map (
            O => \N__42998\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__9767\ : InMux
    port map (
            O => \N__42989\,
            I => \N__42985\
        );

    \I__9766\ : InMux
    port map (
            O => \N__42988\,
            I => \N__42982\
        );

    \I__9765\ : LocalMux
    port map (
            O => \N__42985\,
            I => \N__42977\
        );

    \I__9764\ : LocalMux
    port map (
            O => \N__42982\,
            I => \N__42974\
        );

    \I__9763\ : InMux
    port map (
            O => \N__42981\,
            I => \N__42971\
        );

    \I__9762\ : InMux
    port map (
            O => \N__42980\,
            I => \N__42968\
        );

    \I__9761\ : Span12Mux_h
    port map (
            O => \N__42977\,
            I => \N__42965\
        );

    \I__9760\ : Odrv12
    port map (
            O => \N__42974\,
            I => \phase_controller_slave.hc_time_passed\
        );

    \I__9759\ : LocalMux
    port map (
            O => \N__42971\,
            I => \phase_controller_slave.hc_time_passed\
        );

    \I__9758\ : LocalMux
    port map (
            O => \N__42968\,
            I => \phase_controller_slave.hc_time_passed\
        );

    \I__9757\ : Odrv12
    port map (
            O => \N__42965\,
            I => \phase_controller_slave.hc_time_passed\
        );

    \I__9756\ : InMux
    port map (
            O => \N__42956\,
            I => \N__42953\
        );

    \I__9755\ : LocalMux
    port map (
            O => \N__42953\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19\
        );

    \I__9754\ : CascadeMux
    port map (
            O => \N__42950\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19_cascade_\
        );

    \I__9753\ : InMux
    port map (
            O => \N__42947\,
            I => \N__42944\
        );

    \I__9752\ : LocalMux
    port map (
            O => \N__42944\,
            I => \delay_measurement_inst.delay_tr_timer.N_293\
        );

    \I__9751\ : CascadeMux
    port map (
            O => \N__42941\,
            I => \delay_measurement_inst.N_358_cascade_\
        );

    \I__9750\ : InMux
    port map (
            O => \N__42938\,
            I => \N__42935\
        );

    \I__9749\ : LocalMux
    port map (
            O => \N__42935\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19\
        );

    \I__9748\ : InMux
    port map (
            O => \N__42932\,
            I => \N__42929\
        );

    \I__9747\ : LocalMux
    port map (
            O => \N__42929\,
            I => \N__42926\
        );

    \I__9746\ : Odrv4
    port map (
            O => \N__42926\,
            I => \delay_measurement_inst.N_307\
        );

    \I__9745\ : InMux
    port map (
            O => \N__42923\,
            I => \N__42920\
        );

    \I__9744\ : LocalMux
    port map (
            O => \N__42920\,
            I => \N__42917\
        );

    \I__9743\ : Span12Mux_h
    port map (
            O => \N__42917\,
            I => \N__42914\
        );

    \I__9742\ : Odrv12
    port map (
            O => \N__42914\,
            I => \phase_controller_slave.start_timer_hc_RNO_0_0\
        );

    \I__9741\ : CascadeMux
    port map (
            O => \N__42911\,
            I => \phase_controller_slave.start_timer_hc_0_sqmuxa_cascade_\
        );

    \I__9740\ : InMux
    port map (
            O => \N__42908\,
            I => \N__42905\
        );

    \I__9739\ : LocalMux
    port map (
            O => \N__42905\,
            I => \N__42900\
        );

    \I__9738\ : InMux
    port map (
            O => \N__42904\,
            I => \N__42897\
        );

    \I__9737\ : InMux
    port map (
            O => \N__42903\,
            I => \N__42894\
        );

    \I__9736\ : Span4Mux_v
    port map (
            O => \N__42900\,
            I => \N__42888\
        );

    \I__9735\ : LocalMux
    port map (
            O => \N__42897\,
            I => \N__42885\
        );

    \I__9734\ : LocalMux
    port map (
            O => \N__42894\,
            I => \N__42882\
        );

    \I__9733\ : InMux
    port map (
            O => \N__42893\,
            I => \N__42877\
        );

    \I__9732\ : InMux
    port map (
            O => \N__42892\,
            I => \N__42877\
        );

    \I__9731\ : InMux
    port map (
            O => \N__42891\,
            I => \N__42874\
        );

    \I__9730\ : Odrv4
    port map (
            O => \N__42888\,
            I => phase_controller_inst1_state_4
        );

    \I__9729\ : Odrv4
    port map (
            O => \N__42885\,
            I => phase_controller_inst1_state_4
        );

    \I__9728\ : Odrv12
    port map (
            O => \N__42882\,
            I => phase_controller_inst1_state_4
        );

    \I__9727\ : LocalMux
    port map (
            O => \N__42877\,
            I => phase_controller_inst1_state_4
        );

    \I__9726\ : LocalMux
    port map (
            O => \N__42874\,
            I => phase_controller_inst1_state_4
        );

    \I__9725\ : InMux
    port map (
            O => \N__42863\,
            I => \N__42856\
        );

    \I__9724\ : InMux
    port map (
            O => \N__42862\,
            I => \N__42856\
        );

    \I__9723\ : InMux
    port map (
            O => \N__42861\,
            I => \N__42853\
        );

    \I__9722\ : LocalMux
    port map (
            O => \N__42856\,
            I => \N__42850\
        );

    \I__9721\ : LocalMux
    port map (
            O => \N__42853\,
            I => \N__42847\
        );

    \I__9720\ : Span4Mux_v
    port map (
            O => \N__42850\,
            I => \N__42844\
        );

    \I__9719\ : Span4Mux_v
    port map (
            O => \N__42847\,
            I => \N__42841\
        );

    \I__9718\ : Span4Mux_v
    port map (
            O => \N__42844\,
            I => \N__42838\
        );

    \I__9717\ : Span4Mux_v
    port map (
            O => \N__42841\,
            I => \N__42835\
        );

    \I__9716\ : Span4Mux_v
    port map (
            O => \N__42838\,
            I => \N__42832\
        );

    \I__9715\ : Odrv4
    port map (
            O => \N__42835\,
            I => \il_max_comp2_D2\
        );

    \I__9714\ : Odrv4
    port map (
            O => \N__42832\,
            I => \il_max_comp2_D2\
        );

    \I__9713\ : CascadeMux
    port map (
            O => \N__42827\,
            I => \N__42824\
        );

    \I__9712\ : InMux
    port map (
            O => \N__42824\,
            I => \N__42818\
        );

    \I__9711\ : InMux
    port map (
            O => \N__42823\,
            I => \N__42818\
        );

    \I__9710\ : LocalMux
    port map (
            O => \N__42818\,
            I => \N__42814\
        );

    \I__9709\ : InMux
    port map (
            O => \N__42817\,
            I => \N__42809\
        );

    \I__9708\ : Span4Mux_h
    port map (
            O => \N__42814\,
            I => \N__42806\
        );

    \I__9707\ : InMux
    port map (
            O => \N__42813\,
            I => \N__42803\
        );

    \I__9706\ : InMux
    port map (
            O => \N__42812\,
            I => \N__42800\
        );

    \I__9705\ : LocalMux
    port map (
            O => \N__42809\,
            I => \N__42797\
        );

    \I__9704\ : Span4Mux_h
    port map (
            O => \N__42806\,
            I => \N__42794\
        );

    \I__9703\ : LocalMux
    port map (
            O => \N__42803\,
            I => \phase_controller_slave.stateZ0Z_3\
        );

    \I__9702\ : LocalMux
    port map (
            O => \N__42800\,
            I => \phase_controller_slave.stateZ0Z_3\
        );

    \I__9701\ : Odrv4
    port map (
            O => \N__42797\,
            I => \phase_controller_slave.stateZ0Z_3\
        );

    \I__9700\ : Odrv4
    port map (
            O => \N__42794\,
            I => \phase_controller_slave.stateZ0Z_3\
        );

    \I__9699\ : InMux
    port map (
            O => \N__42785\,
            I => \N__42782\
        );

    \I__9698\ : LocalMux
    port map (
            O => \N__42782\,
            I => \N__42778\
        );

    \I__9697\ : InMux
    port map (
            O => \N__42781\,
            I => \N__42775\
        );

    \I__9696\ : Span4Mux_h
    port map (
            O => \N__42778\,
            I => \N__42771\
        );

    \I__9695\ : LocalMux
    port map (
            O => \N__42775\,
            I => \N__42768\
        );

    \I__9694\ : InMux
    port map (
            O => \N__42774\,
            I => \N__42765\
        );

    \I__9693\ : Span4Mux_v
    port map (
            O => \N__42771\,
            I => \N__42762\
        );

    \I__9692\ : Odrv12
    port map (
            O => \N__42768\,
            I => \phase_controller_slave.stateZ0Z_2\
        );

    \I__9691\ : LocalMux
    port map (
            O => \N__42765\,
            I => \phase_controller_slave.stateZ0Z_2\
        );

    \I__9690\ : Odrv4
    port map (
            O => \N__42762\,
            I => \phase_controller_slave.stateZ0Z_2\
        );

    \I__9689\ : InMux
    port map (
            O => \N__42755\,
            I => \bfn_17_16_0_\
        );

    \I__9688\ : InMux
    port map (
            O => \N__42752\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_24\
        );

    \I__9687\ : InMux
    port map (
            O => \N__42749\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_25\
        );

    \I__9686\ : InMux
    port map (
            O => \N__42746\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_26\
        );

    \I__9685\ : InMux
    port map (
            O => \N__42743\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_27\
        );

    \I__9684\ : InMux
    port map (
            O => \N__42740\,
            I => \N__42724\
        );

    \I__9683\ : InMux
    port map (
            O => \N__42739\,
            I => \N__42724\
        );

    \I__9682\ : InMux
    port map (
            O => \N__42738\,
            I => \N__42724\
        );

    \I__9681\ : InMux
    port map (
            O => \N__42737\,
            I => \N__42724\
        );

    \I__9680\ : InMux
    port map (
            O => \N__42736\,
            I => \N__42693\
        );

    \I__9679\ : InMux
    port map (
            O => \N__42735\,
            I => \N__42693\
        );

    \I__9678\ : InMux
    port map (
            O => \N__42734\,
            I => \N__42693\
        );

    \I__9677\ : InMux
    port map (
            O => \N__42733\,
            I => \N__42693\
        );

    \I__9676\ : LocalMux
    port map (
            O => \N__42724\,
            I => \N__42690\
        );

    \I__9675\ : InMux
    port map (
            O => \N__42723\,
            I => \N__42681\
        );

    \I__9674\ : InMux
    port map (
            O => \N__42722\,
            I => \N__42681\
        );

    \I__9673\ : InMux
    port map (
            O => \N__42721\,
            I => \N__42681\
        );

    \I__9672\ : InMux
    port map (
            O => \N__42720\,
            I => \N__42681\
        );

    \I__9671\ : InMux
    port map (
            O => \N__42719\,
            I => \N__42672\
        );

    \I__9670\ : InMux
    port map (
            O => \N__42718\,
            I => \N__42672\
        );

    \I__9669\ : InMux
    port map (
            O => \N__42717\,
            I => \N__42672\
        );

    \I__9668\ : InMux
    port map (
            O => \N__42716\,
            I => \N__42672\
        );

    \I__9667\ : InMux
    port map (
            O => \N__42715\,
            I => \N__42663\
        );

    \I__9666\ : InMux
    port map (
            O => \N__42714\,
            I => \N__42663\
        );

    \I__9665\ : InMux
    port map (
            O => \N__42713\,
            I => \N__42663\
        );

    \I__9664\ : InMux
    port map (
            O => \N__42712\,
            I => \N__42663\
        );

    \I__9663\ : InMux
    port map (
            O => \N__42711\,
            I => \N__42654\
        );

    \I__9662\ : InMux
    port map (
            O => \N__42710\,
            I => \N__42654\
        );

    \I__9661\ : InMux
    port map (
            O => \N__42709\,
            I => \N__42654\
        );

    \I__9660\ : InMux
    port map (
            O => \N__42708\,
            I => \N__42654\
        );

    \I__9659\ : InMux
    port map (
            O => \N__42707\,
            I => \N__42649\
        );

    \I__9658\ : InMux
    port map (
            O => \N__42706\,
            I => \N__42649\
        );

    \I__9657\ : InMux
    port map (
            O => \N__42705\,
            I => \N__42640\
        );

    \I__9656\ : InMux
    port map (
            O => \N__42704\,
            I => \N__42640\
        );

    \I__9655\ : InMux
    port map (
            O => \N__42703\,
            I => \N__42640\
        );

    \I__9654\ : InMux
    port map (
            O => \N__42702\,
            I => \N__42640\
        );

    \I__9653\ : LocalMux
    port map (
            O => \N__42693\,
            I => \N__42633\
        );

    \I__9652\ : Span4Mux_h
    port map (
            O => \N__42690\,
            I => \N__42633\
        );

    \I__9651\ : LocalMux
    port map (
            O => \N__42681\,
            I => \N__42633\
        );

    \I__9650\ : LocalMux
    port map (
            O => \N__42672\,
            I => \N__42626\
        );

    \I__9649\ : LocalMux
    port map (
            O => \N__42663\,
            I => \N__42626\
        );

    \I__9648\ : LocalMux
    port map (
            O => \N__42654\,
            I => \N__42626\
        );

    \I__9647\ : LocalMux
    port map (
            O => \N__42649\,
            I => \N__42621\
        );

    \I__9646\ : LocalMux
    port map (
            O => \N__42640\,
            I => \N__42621\
        );

    \I__9645\ : Span4Mux_v
    port map (
            O => \N__42633\,
            I => \N__42616\
        );

    \I__9644\ : Span4Mux_v
    port map (
            O => \N__42626\,
            I => \N__42616\
        );

    \I__9643\ : Span4Mux_h
    port map (
            O => \N__42621\,
            I => \N__42613\
        );

    \I__9642\ : Span4Mux_h
    port map (
            O => \N__42616\,
            I => \N__42610\
        );

    \I__9641\ : Span4Mux_v
    port map (
            O => \N__42613\,
            I => \N__42607\
        );

    \I__9640\ : Odrv4
    port map (
            O => \N__42610\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__9639\ : Odrv4
    port map (
            O => \N__42607\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__9638\ : InMux
    port map (
            O => \N__42602\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_28\
        );

    \I__9637\ : CEMux
    port map (
            O => \N__42599\,
            I => \N__42596\
        );

    \I__9636\ : LocalMux
    port map (
            O => \N__42596\,
            I => \N__42592\
        );

    \I__9635\ : CEMux
    port map (
            O => \N__42595\,
            I => \N__42587\
        );

    \I__9634\ : Span4Mux_h
    port map (
            O => \N__42592\,
            I => \N__42584\
        );

    \I__9633\ : CEMux
    port map (
            O => \N__42591\,
            I => \N__42581\
        );

    \I__9632\ : CEMux
    port map (
            O => \N__42590\,
            I => \N__42578\
        );

    \I__9631\ : LocalMux
    port map (
            O => \N__42587\,
            I => \N__42575\
        );

    \I__9630\ : Span4Mux_h
    port map (
            O => \N__42584\,
            I => \N__42572\
        );

    \I__9629\ : LocalMux
    port map (
            O => \N__42581\,
            I => \N__42569\
        );

    \I__9628\ : LocalMux
    port map (
            O => \N__42578\,
            I => \N__42566\
        );

    \I__9627\ : Span4Mux_v
    port map (
            O => \N__42575\,
            I => \N__42563\
        );

    \I__9626\ : Sp12to4
    port map (
            O => \N__42572\,
            I => \N__42560\
        );

    \I__9625\ : Span4Mux_h
    port map (
            O => \N__42569\,
            I => \N__42557\
        );

    \I__9624\ : Span4Mux_h
    port map (
            O => \N__42566\,
            I => \N__42554\
        );

    \I__9623\ : Span4Mux_v
    port map (
            O => \N__42563\,
            I => \N__42551\
        );

    \I__9622\ : Span12Mux_v
    port map (
            O => \N__42560\,
            I => \N__42548\
        );

    \I__9621\ : Span4Mux_v
    port map (
            O => \N__42557\,
            I => \N__42545\
        );

    \I__9620\ : Span4Mux_v
    port map (
            O => \N__42554\,
            I => \N__42542\
        );

    \I__9619\ : Odrv4
    port map (
            O => \N__42551\,
            I => \delay_measurement_inst.delay_tr_timer.N_338_i\
        );

    \I__9618\ : Odrv12
    port map (
            O => \N__42548\,
            I => \delay_measurement_inst.delay_tr_timer.N_338_i\
        );

    \I__9617\ : Odrv4
    port map (
            O => \N__42545\,
            I => \delay_measurement_inst.delay_tr_timer.N_338_i\
        );

    \I__9616\ : Odrv4
    port map (
            O => \N__42542\,
            I => \delay_measurement_inst.delay_tr_timer.N_338_i\
        );

    \I__9615\ : InMux
    port map (
            O => \N__42533\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_14\
        );

    \I__9614\ : InMux
    port map (
            O => \N__42530\,
            I => \bfn_17_15_0_\
        );

    \I__9613\ : InMux
    port map (
            O => \N__42527\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_16\
        );

    \I__9612\ : InMux
    port map (
            O => \N__42524\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_17\
        );

    \I__9611\ : InMux
    port map (
            O => \N__42521\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_18\
        );

    \I__9610\ : InMux
    port map (
            O => \N__42518\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_19\
        );

    \I__9609\ : InMux
    port map (
            O => \N__42515\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_20\
        );

    \I__9608\ : InMux
    port map (
            O => \N__42512\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_21\
        );

    \I__9607\ : InMux
    port map (
            O => \N__42509\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_22\
        );

    \I__9606\ : InMux
    port map (
            O => \N__42506\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_5\
        );

    \I__9605\ : InMux
    port map (
            O => \N__42503\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_6\
        );

    \I__9604\ : InMux
    port map (
            O => \N__42500\,
            I => \bfn_17_14_0_\
        );

    \I__9603\ : InMux
    port map (
            O => \N__42497\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_8\
        );

    \I__9602\ : InMux
    port map (
            O => \N__42494\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_9\
        );

    \I__9601\ : InMux
    port map (
            O => \N__42491\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_10\
        );

    \I__9600\ : InMux
    port map (
            O => \N__42488\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_11\
        );

    \I__9599\ : InMux
    port map (
            O => \N__42485\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_12\
        );

    \I__9598\ : InMux
    port map (
            O => \N__42482\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_13\
        );

    \I__9597\ : InMux
    port map (
            O => \N__42479\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__9596\ : InMux
    port map (
            O => \N__42476\,
            I => \N__42471\
        );

    \I__9595\ : InMux
    port map (
            O => \N__42475\,
            I => \N__42467\
        );

    \I__9594\ : InMux
    port map (
            O => \N__42474\,
            I => \N__42464\
        );

    \I__9593\ : LocalMux
    port map (
            O => \N__42471\,
            I => \N__42461\
        );

    \I__9592\ : InMux
    port map (
            O => \N__42470\,
            I => \N__42458\
        );

    \I__9591\ : LocalMux
    port map (
            O => \N__42467\,
            I => \N__42455\
        );

    \I__9590\ : LocalMux
    port map (
            O => \N__42464\,
            I => \N__42448\
        );

    \I__9589\ : Span4Mux_h
    port map (
            O => \N__42461\,
            I => \N__42448\
        );

    \I__9588\ : LocalMux
    port map (
            O => \N__42458\,
            I => \N__42448\
        );

    \I__9587\ : Span4Mux_h
    port map (
            O => \N__42455\,
            I => \N__42445\
        );

    \I__9586\ : Span4Mux_v
    port map (
            O => \N__42448\,
            I => \N__42442\
        );

    \I__9585\ : Odrv4
    port map (
            O => \N__42445\,
            I => \delay_measurement_inst.elapsed_time_hc_4\
        );

    \I__9584\ : Odrv4
    port map (
            O => \N__42442\,
            I => \delay_measurement_inst.elapsed_time_hc_4\
        );

    \I__9583\ : InMux
    port map (
            O => \N__42437\,
            I => \N__42433\
        );

    \I__9582\ : InMux
    port map (
            O => \N__42436\,
            I => \N__42428\
        );

    \I__9581\ : LocalMux
    port map (
            O => \N__42433\,
            I => \N__42425\
        );

    \I__9580\ : InMux
    port map (
            O => \N__42432\,
            I => \N__42422\
        );

    \I__9579\ : InMux
    port map (
            O => \N__42431\,
            I => \N__42419\
        );

    \I__9578\ : LocalMux
    port map (
            O => \N__42428\,
            I => \N__42416\
        );

    \I__9577\ : Span4Mux_h
    port map (
            O => \N__42425\,
            I => \N__42409\
        );

    \I__9576\ : LocalMux
    port map (
            O => \N__42422\,
            I => \N__42409\
        );

    \I__9575\ : LocalMux
    port map (
            O => \N__42419\,
            I => \N__42409\
        );

    \I__9574\ : Span4Mux_h
    port map (
            O => \N__42416\,
            I => \N__42404\
        );

    \I__9573\ : Span4Mux_v
    port map (
            O => \N__42409\,
            I => \N__42404\
        );

    \I__9572\ : Odrv4
    port map (
            O => \N__42404\,
            I => \delay_measurement_inst.elapsed_time_hc_3\
        );

    \I__9571\ : CascadeMux
    port map (
            O => \N__42401\,
            I => \N__42398\
        );

    \I__9570\ : InMux
    port map (
            O => \N__42398\,
            I => \N__42395\
        );

    \I__9569\ : LocalMux
    port map (
            O => \N__42395\,
            I => \N__42392\
        );

    \I__9568\ : Span4Mux_h
    port map (
            O => \N__42392\,
            I => \N__42388\
        );

    \I__9567\ : InMux
    port map (
            O => \N__42391\,
            I => \N__42385\
        );

    \I__9566\ : Odrv4
    port map (
            O => \N__42388\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto5_2\
        );

    \I__9565\ : LocalMux
    port map (
            O => \N__42385\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto5_2\
        );

    \I__9564\ : CascadeMux
    port map (
            O => \N__42380\,
            I => \N__42376\
        );

    \I__9563\ : InMux
    port map (
            O => \N__42379\,
            I => \N__42373\
        );

    \I__9562\ : InMux
    port map (
            O => \N__42376\,
            I => \N__42370\
        );

    \I__9561\ : LocalMux
    port map (
            O => \N__42373\,
            I => \N__42366\
        );

    \I__9560\ : LocalMux
    port map (
            O => \N__42370\,
            I => \N__42363\
        );

    \I__9559\ : InMux
    port map (
            O => \N__42369\,
            I => \N__42360\
        );

    \I__9558\ : Span4Mux_h
    port map (
            O => \N__42366\,
            I => \N__42357\
        );

    \I__9557\ : Span12Mux_v
    port map (
            O => \N__42363\,
            I => \N__42354\
        );

    \I__9556\ : LocalMux
    port map (
            O => \N__42360\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1\
        );

    \I__9555\ : Odrv4
    port map (
            O => \N__42357\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1\
        );

    \I__9554\ : Odrv12
    port map (
            O => \N__42354\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1\
        );

    \I__9553\ : CascadeMux
    port map (
            O => \N__42347\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIB3GH4Z0Z_3_cascade_\
        );

    \I__9552\ : InMux
    port map (
            O => \N__42344\,
            I => \N__42341\
        );

    \I__9551\ : LocalMux
    port map (
            O => \N__42341\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_7_0\
        );

    \I__9550\ : InMux
    port map (
            O => \N__42338\,
            I => \bfn_17_13_0_\
        );

    \I__9549\ : InMux
    port map (
            O => \N__42335\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_0\
        );

    \I__9548\ : InMux
    port map (
            O => \N__42332\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_1\
        );

    \I__9547\ : InMux
    port map (
            O => \N__42329\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_2\
        );

    \I__9546\ : InMux
    port map (
            O => \N__42326\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_3\
        );

    \I__9545\ : InMux
    port map (
            O => \N__42323\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_4\
        );

    \I__9544\ : CascadeMux
    port map (
            O => \N__42320\,
            I => \N__42315\
        );

    \I__9543\ : InMux
    port map (
            O => \N__42319\,
            I => \N__42312\
        );

    \I__9542\ : InMux
    port map (
            O => \N__42318\,
            I => \N__42309\
        );

    \I__9541\ : InMux
    port map (
            O => \N__42315\,
            I => \N__42306\
        );

    \I__9540\ : LocalMux
    port map (
            O => \N__42312\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__9539\ : LocalMux
    port map (
            O => \N__42309\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__9538\ : LocalMux
    port map (
            O => \N__42306\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__9537\ : InMux
    port map (
            O => \N__42299\,
            I => \N__42296\
        );

    \I__9536\ : LocalMux
    port map (
            O => \N__42296\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__9535\ : InMux
    port map (
            O => \N__42293\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__9534\ : CascadeMux
    port map (
            O => \N__42290\,
            I => \N__42285\
        );

    \I__9533\ : InMux
    port map (
            O => \N__42289\,
            I => \N__42282\
        );

    \I__9532\ : InMux
    port map (
            O => \N__42288\,
            I => \N__42279\
        );

    \I__9531\ : InMux
    port map (
            O => \N__42285\,
            I => \N__42276\
        );

    \I__9530\ : LocalMux
    port map (
            O => \N__42282\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__9529\ : LocalMux
    port map (
            O => \N__42279\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__9528\ : LocalMux
    port map (
            O => \N__42276\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__9527\ : InMux
    port map (
            O => \N__42269\,
            I => \N__42266\
        );

    \I__9526\ : LocalMux
    port map (
            O => \N__42266\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__9525\ : InMux
    port map (
            O => \N__42263\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__9524\ : CascadeMux
    port map (
            O => \N__42260\,
            I => \N__42255\
        );

    \I__9523\ : InMux
    port map (
            O => \N__42259\,
            I => \N__42252\
        );

    \I__9522\ : InMux
    port map (
            O => \N__42258\,
            I => \N__42249\
        );

    \I__9521\ : InMux
    port map (
            O => \N__42255\,
            I => \N__42246\
        );

    \I__9520\ : LocalMux
    port map (
            O => \N__42252\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__9519\ : LocalMux
    port map (
            O => \N__42249\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__9518\ : LocalMux
    port map (
            O => \N__42246\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__9517\ : InMux
    port map (
            O => \N__42239\,
            I => \N__42236\
        );

    \I__9516\ : LocalMux
    port map (
            O => \N__42236\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__9515\ : InMux
    port map (
            O => \N__42233\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__9514\ : CascadeMux
    port map (
            O => \N__42230\,
            I => \N__42225\
        );

    \I__9513\ : InMux
    port map (
            O => \N__42229\,
            I => \N__42222\
        );

    \I__9512\ : InMux
    port map (
            O => \N__42228\,
            I => \N__42219\
        );

    \I__9511\ : InMux
    port map (
            O => \N__42225\,
            I => \N__42216\
        );

    \I__9510\ : LocalMux
    port map (
            O => \N__42222\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__9509\ : LocalMux
    port map (
            O => \N__42219\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__9508\ : LocalMux
    port map (
            O => \N__42216\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__9507\ : InMux
    port map (
            O => \N__42209\,
            I => \N__42206\
        );

    \I__9506\ : LocalMux
    port map (
            O => \N__42206\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__9505\ : InMux
    port map (
            O => \N__42203\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__9504\ : CascadeMux
    port map (
            O => \N__42200\,
            I => \N__42195\
        );

    \I__9503\ : InMux
    port map (
            O => \N__42199\,
            I => \N__42192\
        );

    \I__9502\ : InMux
    port map (
            O => \N__42198\,
            I => \N__42189\
        );

    \I__9501\ : InMux
    port map (
            O => \N__42195\,
            I => \N__42186\
        );

    \I__9500\ : LocalMux
    port map (
            O => \N__42192\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__9499\ : LocalMux
    port map (
            O => \N__42189\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__9498\ : LocalMux
    port map (
            O => \N__42186\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__9497\ : InMux
    port map (
            O => \N__42179\,
            I => \N__42176\
        );

    \I__9496\ : LocalMux
    port map (
            O => \N__42176\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__9495\ : InMux
    port map (
            O => \N__42173\,
            I => \bfn_17_11_0_\
        );

    \I__9494\ : CascadeMux
    port map (
            O => \N__42170\,
            I => \N__42165\
        );

    \I__9493\ : InMux
    port map (
            O => \N__42169\,
            I => \N__42162\
        );

    \I__9492\ : InMux
    port map (
            O => \N__42168\,
            I => \N__42159\
        );

    \I__9491\ : InMux
    port map (
            O => \N__42165\,
            I => \N__42156\
        );

    \I__9490\ : LocalMux
    port map (
            O => \N__42162\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__9489\ : LocalMux
    port map (
            O => \N__42159\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__9488\ : LocalMux
    port map (
            O => \N__42156\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__9487\ : InMux
    port map (
            O => \N__42149\,
            I => \N__42146\
        );

    \I__9486\ : LocalMux
    port map (
            O => \N__42146\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__9485\ : InMux
    port map (
            O => \N__42143\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__9484\ : CascadeMux
    port map (
            O => \N__42140\,
            I => \N__42135\
        );

    \I__9483\ : InMux
    port map (
            O => \N__42139\,
            I => \N__42132\
        );

    \I__9482\ : InMux
    port map (
            O => \N__42138\,
            I => \N__42129\
        );

    \I__9481\ : InMux
    port map (
            O => \N__42135\,
            I => \N__42126\
        );

    \I__9480\ : LocalMux
    port map (
            O => \N__42132\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__9479\ : LocalMux
    port map (
            O => \N__42129\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__9478\ : LocalMux
    port map (
            O => \N__42126\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__9477\ : CascadeMux
    port map (
            O => \N__42119\,
            I => \N__42115\
        );

    \I__9476\ : InMux
    port map (
            O => \N__42118\,
            I => \N__42112\
        );

    \I__9475\ : InMux
    port map (
            O => \N__42115\,
            I => \N__42109\
        );

    \I__9474\ : LocalMux
    port map (
            O => \N__42112\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__9473\ : LocalMux
    port map (
            O => \N__42109\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__9472\ : InMux
    port map (
            O => \N__42104\,
            I => \N__42101\
        );

    \I__9471\ : LocalMux
    port map (
            O => \N__42101\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__9470\ : InMux
    port map (
            O => \N__42098\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__9469\ : CascadeMux
    port map (
            O => \N__42095\,
            I => \N__42090\
        );

    \I__9468\ : InMux
    port map (
            O => \N__42094\,
            I => \N__42087\
        );

    \I__9467\ : InMux
    port map (
            O => \N__42093\,
            I => \N__42084\
        );

    \I__9466\ : InMux
    port map (
            O => \N__42090\,
            I => \N__42081\
        );

    \I__9465\ : LocalMux
    port map (
            O => \N__42087\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__9464\ : LocalMux
    port map (
            O => \N__42084\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__9463\ : LocalMux
    port map (
            O => \N__42081\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__9462\ : CascadeMux
    port map (
            O => \N__42074\,
            I => \N__42070\
        );

    \I__9461\ : InMux
    port map (
            O => \N__42073\,
            I => \N__42067\
        );

    \I__9460\ : InMux
    port map (
            O => \N__42070\,
            I => \N__42064\
        );

    \I__9459\ : LocalMux
    port map (
            O => \N__42067\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__9458\ : LocalMux
    port map (
            O => \N__42064\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__9457\ : CascadeMux
    port map (
            O => \N__42059\,
            I => \N__42056\
        );

    \I__9456\ : InMux
    port map (
            O => \N__42056\,
            I => \N__42053\
        );

    \I__9455\ : LocalMux
    port map (
            O => \N__42053\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_30\
        );

    \I__9454\ : InMux
    port map (
            O => \N__42050\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__9453\ : CascadeMux
    port map (
            O => \N__42047\,
            I => \N__42042\
        );

    \I__9452\ : InMux
    port map (
            O => \N__42046\,
            I => \N__42039\
        );

    \I__9451\ : InMux
    port map (
            O => \N__42045\,
            I => \N__42036\
        );

    \I__9450\ : InMux
    port map (
            O => \N__42042\,
            I => \N__42033\
        );

    \I__9449\ : LocalMux
    port map (
            O => \N__42039\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__9448\ : LocalMux
    port map (
            O => \N__42036\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__9447\ : LocalMux
    port map (
            O => \N__42033\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__9446\ : InMux
    port map (
            O => \N__42026\,
            I => \N__42023\
        );

    \I__9445\ : LocalMux
    port map (
            O => \N__42023\,
            I => \N__42020\
        );

    \I__9444\ : Span4Mux_h
    port map (
            O => \N__42020\,
            I => \N__42017\
        );

    \I__9443\ : Span4Mux_h
    port map (
            O => \N__42017\,
            I => \N__42013\
        );

    \I__9442\ : CascadeMux
    port map (
            O => \N__42016\,
            I => \N__42007\
        );

    \I__9441\ : Span4Mux_v
    port map (
            O => \N__42013\,
            I => \N__42004\
        );

    \I__9440\ : InMux
    port map (
            O => \N__42012\,
            I => \N__42001\
        );

    \I__9439\ : InMux
    port map (
            O => \N__42011\,
            I => \N__41998\
        );

    \I__9438\ : CascadeMux
    port map (
            O => \N__42010\,
            I => \N__41995\
        );

    \I__9437\ : InMux
    port map (
            O => \N__42007\,
            I => \N__41992\
        );

    \I__9436\ : Span4Mux_h
    port map (
            O => \N__42004\,
            I => \N__41987\
        );

    \I__9435\ : LocalMux
    port map (
            O => \N__42001\,
            I => \N__41987\
        );

    \I__9434\ : LocalMux
    port map (
            O => \N__41998\,
            I => \N__41984\
        );

    \I__9433\ : InMux
    port map (
            O => \N__41995\,
            I => \N__41981\
        );

    \I__9432\ : LocalMux
    port map (
            O => \N__41992\,
            I => \N__41978\
        );

    \I__9431\ : Span4Mux_v
    port map (
            O => \N__41987\,
            I => \N__41975\
        );

    \I__9430\ : Span4Mux_v
    port map (
            O => \N__41984\,
            I => \N__41970\
        );

    \I__9429\ : LocalMux
    port map (
            O => \N__41981\,
            I => \N__41970\
        );

    \I__9428\ : Odrv12
    port map (
            O => \N__41978\,
            I => \delay_measurement_inst.delay_hc_reg3lto15\
        );

    \I__9427\ : Odrv4
    port map (
            O => \N__41975\,
            I => \delay_measurement_inst.delay_hc_reg3lto15\
        );

    \I__9426\ : Odrv4
    port map (
            O => \N__41970\,
            I => \delay_measurement_inst.delay_hc_reg3lto15\
        );

    \I__9425\ : InMux
    port map (
            O => \N__41963\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__9424\ : CascadeMux
    port map (
            O => \N__41960\,
            I => \N__41955\
        );

    \I__9423\ : InMux
    port map (
            O => \N__41959\,
            I => \N__41952\
        );

    \I__9422\ : InMux
    port map (
            O => \N__41958\,
            I => \N__41949\
        );

    \I__9421\ : InMux
    port map (
            O => \N__41955\,
            I => \N__41946\
        );

    \I__9420\ : LocalMux
    port map (
            O => \N__41952\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__9419\ : LocalMux
    port map (
            O => \N__41949\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__9418\ : LocalMux
    port map (
            O => \N__41946\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__9417\ : InMux
    port map (
            O => \N__41939\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__9416\ : CascadeMux
    port map (
            O => \N__41936\,
            I => \N__41931\
        );

    \I__9415\ : InMux
    port map (
            O => \N__41935\,
            I => \N__41928\
        );

    \I__9414\ : InMux
    port map (
            O => \N__41934\,
            I => \N__41925\
        );

    \I__9413\ : InMux
    port map (
            O => \N__41931\,
            I => \N__41922\
        );

    \I__9412\ : LocalMux
    port map (
            O => \N__41928\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__9411\ : LocalMux
    port map (
            O => \N__41925\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__9410\ : LocalMux
    port map (
            O => \N__41922\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__9409\ : InMux
    port map (
            O => \N__41915\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__9408\ : CascadeMux
    port map (
            O => \N__41912\,
            I => \N__41907\
        );

    \I__9407\ : InMux
    port map (
            O => \N__41911\,
            I => \N__41904\
        );

    \I__9406\ : InMux
    port map (
            O => \N__41910\,
            I => \N__41901\
        );

    \I__9405\ : InMux
    port map (
            O => \N__41907\,
            I => \N__41898\
        );

    \I__9404\ : LocalMux
    port map (
            O => \N__41904\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__9403\ : LocalMux
    port map (
            O => \N__41901\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__9402\ : LocalMux
    port map (
            O => \N__41898\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__9401\ : InMux
    port map (
            O => \N__41891\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__9400\ : CascadeMux
    port map (
            O => \N__41888\,
            I => \N__41883\
        );

    \I__9399\ : InMux
    port map (
            O => \N__41887\,
            I => \N__41880\
        );

    \I__9398\ : InMux
    port map (
            O => \N__41886\,
            I => \N__41877\
        );

    \I__9397\ : InMux
    port map (
            O => \N__41883\,
            I => \N__41874\
        );

    \I__9396\ : LocalMux
    port map (
            O => \N__41880\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__9395\ : LocalMux
    port map (
            O => \N__41877\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__9394\ : LocalMux
    port map (
            O => \N__41874\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__9393\ : InMux
    port map (
            O => \N__41867\,
            I => \bfn_17_10_0_\
        );

    \I__9392\ : CascadeMux
    port map (
            O => \N__41864\,
            I => \N__41859\
        );

    \I__9391\ : InMux
    port map (
            O => \N__41863\,
            I => \N__41856\
        );

    \I__9390\ : InMux
    port map (
            O => \N__41862\,
            I => \N__41853\
        );

    \I__9389\ : InMux
    port map (
            O => \N__41859\,
            I => \N__41850\
        );

    \I__9388\ : LocalMux
    port map (
            O => \N__41856\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__9387\ : LocalMux
    port map (
            O => \N__41853\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__9386\ : LocalMux
    port map (
            O => \N__41850\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__9385\ : CascadeMux
    port map (
            O => \N__41843\,
            I => \N__41840\
        );

    \I__9384\ : InMux
    port map (
            O => \N__41840\,
            I => \N__41837\
        );

    \I__9383\ : LocalMux
    port map (
            O => \N__41837\,
            I => \N__41833\
        );

    \I__9382\ : InMux
    port map (
            O => \N__41836\,
            I => \N__41830\
        );

    \I__9381\ : Odrv4
    port map (
            O => \N__41833\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__9380\ : LocalMux
    port map (
            O => \N__41830\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__9379\ : InMux
    port map (
            O => \N__41825\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__9378\ : CascadeMux
    port map (
            O => \N__41822\,
            I => \N__41817\
        );

    \I__9377\ : InMux
    port map (
            O => \N__41821\,
            I => \N__41814\
        );

    \I__9376\ : InMux
    port map (
            O => \N__41820\,
            I => \N__41811\
        );

    \I__9375\ : InMux
    port map (
            O => \N__41817\,
            I => \N__41808\
        );

    \I__9374\ : LocalMux
    port map (
            O => \N__41814\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__9373\ : LocalMux
    port map (
            O => \N__41811\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__9372\ : LocalMux
    port map (
            O => \N__41808\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__9371\ : InMux
    port map (
            O => \N__41801\,
            I => \N__41798\
        );

    \I__9370\ : LocalMux
    port map (
            O => \N__41798\,
            I => \N__41794\
        );

    \I__9369\ : InMux
    port map (
            O => \N__41797\,
            I => \N__41791\
        );

    \I__9368\ : Span4Mux_v
    port map (
            O => \N__41794\,
            I => \N__41788\
        );

    \I__9367\ : LocalMux
    port map (
            O => \N__41791\,
            I => \N__41785\
        );

    \I__9366\ : Odrv4
    port map (
            O => \N__41788\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__9365\ : Odrv4
    port map (
            O => \N__41785\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__9364\ : InMux
    port map (
            O => \N__41780\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__9363\ : CascadeMux
    port map (
            O => \N__41777\,
            I => \N__41772\
        );

    \I__9362\ : InMux
    port map (
            O => \N__41776\,
            I => \N__41769\
        );

    \I__9361\ : InMux
    port map (
            O => \N__41775\,
            I => \N__41766\
        );

    \I__9360\ : InMux
    port map (
            O => \N__41772\,
            I => \N__41763\
        );

    \I__9359\ : LocalMux
    port map (
            O => \N__41769\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__9358\ : LocalMux
    port map (
            O => \N__41766\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__9357\ : LocalMux
    port map (
            O => \N__41763\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__9356\ : InMux
    port map (
            O => \N__41756\,
            I => \N__41753\
        );

    \I__9355\ : LocalMux
    port map (
            O => \N__41753\,
            I => \N__41749\
        );

    \I__9354\ : CascadeMux
    port map (
            O => \N__41752\,
            I => \N__41746\
        );

    \I__9353\ : Span4Mux_v
    port map (
            O => \N__41749\,
            I => \N__41743\
        );

    \I__9352\ : InMux
    port map (
            O => \N__41746\,
            I => \N__41740\
        );

    \I__9351\ : Odrv4
    port map (
            O => \N__41743\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__9350\ : LocalMux
    port map (
            O => \N__41740\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__9349\ : InMux
    port map (
            O => \N__41735\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__9348\ : CascadeMux
    port map (
            O => \N__41732\,
            I => \N__41727\
        );

    \I__9347\ : InMux
    port map (
            O => \N__41731\,
            I => \N__41724\
        );

    \I__9346\ : InMux
    port map (
            O => \N__41730\,
            I => \N__41721\
        );

    \I__9345\ : InMux
    port map (
            O => \N__41727\,
            I => \N__41718\
        );

    \I__9344\ : LocalMux
    port map (
            O => \N__41724\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__9343\ : LocalMux
    port map (
            O => \N__41721\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__9342\ : LocalMux
    port map (
            O => \N__41718\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__9341\ : CascadeMux
    port map (
            O => \N__41711\,
            I => \N__41708\
        );

    \I__9340\ : InMux
    port map (
            O => \N__41708\,
            I => \N__41702\
        );

    \I__9339\ : InMux
    port map (
            O => \N__41707\,
            I => \N__41699\
        );

    \I__9338\ : InMux
    port map (
            O => \N__41706\,
            I => \N__41693\
        );

    \I__9337\ : InMux
    port map (
            O => \N__41705\,
            I => \N__41693\
        );

    \I__9336\ : LocalMux
    port map (
            O => \N__41702\,
            I => \N__41688\
        );

    \I__9335\ : LocalMux
    port map (
            O => \N__41699\,
            I => \N__41688\
        );

    \I__9334\ : InMux
    port map (
            O => \N__41698\,
            I => \N__41685\
        );

    \I__9333\ : LocalMux
    port map (
            O => \N__41693\,
            I => \N__41682\
        );

    \I__9332\ : Span4Mux_v
    port map (
            O => \N__41688\,
            I => \N__41679\
        );

    \I__9331\ : LocalMux
    port map (
            O => \N__41685\,
            I => \N__41674\
        );

    \I__9330\ : Span4Mux_h
    port map (
            O => \N__41682\,
            I => \N__41674\
        );

    \I__9329\ : Odrv4
    port map (
            O => \N__41679\,
            I => \delay_measurement_inst.elapsed_time_hc_7\
        );

    \I__9328\ : Odrv4
    port map (
            O => \N__41674\,
            I => \delay_measurement_inst.elapsed_time_hc_7\
        );

    \I__9327\ : InMux
    port map (
            O => \N__41669\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__9326\ : CascadeMux
    port map (
            O => \N__41666\,
            I => \N__41661\
        );

    \I__9325\ : InMux
    port map (
            O => \N__41665\,
            I => \N__41658\
        );

    \I__9324\ : InMux
    port map (
            O => \N__41664\,
            I => \N__41655\
        );

    \I__9323\ : InMux
    port map (
            O => \N__41661\,
            I => \N__41652\
        );

    \I__9322\ : LocalMux
    port map (
            O => \N__41658\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__9321\ : LocalMux
    port map (
            O => \N__41655\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__9320\ : LocalMux
    port map (
            O => \N__41652\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__9319\ : CascadeMux
    port map (
            O => \N__41645\,
            I => \N__41639\
        );

    \I__9318\ : InMux
    port map (
            O => \N__41644\,
            I => \N__41635\
        );

    \I__9317\ : InMux
    port map (
            O => \N__41643\,
            I => \N__41632\
        );

    \I__9316\ : InMux
    port map (
            O => \N__41642\,
            I => \N__41629\
        );

    \I__9315\ : InMux
    port map (
            O => \N__41639\,
            I => \N__41624\
        );

    \I__9314\ : InMux
    port map (
            O => \N__41638\,
            I => \N__41624\
        );

    \I__9313\ : LocalMux
    port map (
            O => \N__41635\,
            I => \N__41619\
        );

    \I__9312\ : LocalMux
    port map (
            O => \N__41632\,
            I => \N__41619\
        );

    \I__9311\ : LocalMux
    port map (
            O => \N__41629\,
            I => \N__41614\
        );

    \I__9310\ : LocalMux
    port map (
            O => \N__41624\,
            I => \N__41614\
        );

    \I__9309\ : Span4Mux_v
    port map (
            O => \N__41619\,
            I => \N__41611\
        );

    \I__9308\ : Span4Mux_h
    port map (
            O => \N__41614\,
            I => \N__41608\
        );

    \I__9307\ : Odrv4
    port map (
            O => \N__41611\,
            I => \delay_measurement_inst.elapsed_time_hc_8\
        );

    \I__9306\ : Odrv4
    port map (
            O => \N__41608\,
            I => \delay_measurement_inst.elapsed_time_hc_8\
        );

    \I__9305\ : InMux
    port map (
            O => \N__41603\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__9304\ : CascadeMux
    port map (
            O => \N__41600\,
            I => \N__41595\
        );

    \I__9303\ : InMux
    port map (
            O => \N__41599\,
            I => \N__41592\
        );

    \I__9302\ : InMux
    port map (
            O => \N__41598\,
            I => \N__41589\
        );

    \I__9301\ : InMux
    port map (
            O => \N__41595\,
            I => \N__41586\
        );

    \I__9300\ : LocalMux
    port map (
            O => \N__41592\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__9299\ : LocalMux
    port map (
            O => \N__41589\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__9298\ : LocalMux
    port map (
            O => \N__41586\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__9297\ : InMux
    port map (
            O => \N__41579\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__9296\ : CascadeMux
    port map (
            O => \N__41576\,
            I => \N__41571\
        );

    \I__9295\ : InMux
    port map (
            O => \N__41575\,
            I => \N__41568\
        );

    \I__9294\ : InMux
    port map (
            O => \N__41574\,
            I => \N__41565\
        );

    \I__9293\ : InMux
    port map (
            O => \N__41571\,
            I => \N__41562\
        );

    \I__9292\ : LocalMux
    port map (
            O => \N__41568\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__9291\ : LocalMux
    port map (
            O => \N__41565\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__9290\ : LocalMux
    port map (
            O => \N__41562\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__9289\ : CascadeMux
    port map (
            O => \N__41555\,
            I => \N__41551\
        );

    \I__9288\ : CascadeMux
    port map (
            O => \N__41554\,
            I => \N__41547\
        );

    \I__9287\ : InMux
    port map (
            O => \N__41551\,
            I => \N__41544\
        );

    \I__9286\ : InMux
    port map (
            O => \N__41550\,
            I => \N__41541\
        );

    \I__9285\ : InMux
    port map (
            O => \N__41547\,
            I => \N__41538\
        );

    \I__9284\ : LocalMux
    port map (
            O => \N__41544\,
            I => \N__41535\
        );

    \I__9283\ : LocalMux
    port map (
            O => \N__41541\,
            I => \N__41530\
        );

    \I__9282\ : LocalMux
    port map (
            O => \N__41538\,
            I => \N__41530\
        );

    \I__9281\ : Span4Mux_h
    port map (
            O => \N__41535\,
            I => \N__41527\
        );

    \I__9280\ : Span4Mux_h
    port map (
            O => \N__41530\,
            I => \N__41524\
        );

    \I__9279\ : Odrv4
    port map (
            O => \N__41527\,
            I => \delay_measurement_inst.elapsed_time_hc_10\
        );

    \I__9278\ : Odrv4
    port map (
            O => \N__41524\,
            I => \delay_measurement_inst.elapsed_time_hc_10\
        );

    \I__9277\ : InMux
    port map (
            O => \N__41519\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__9276\ : CascadeMux
    port map (
            O => \N__41516\,
            I => \N__41511\
        );

    \I__9275\ : InMux
    port map (
            O => \N__41515\,
            I => \N__41508\
        );

    \I__9274\ : InMux
    port map (
            O => \N__41514\,
            I => \N__41505\
        );

    \I__9273\ : InMux
    port map (
            O => \N__41511\,
            I => \N__41502\
        );

    \I__9272\ : LocalMux
    port map (
            O => \N__41508\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__9271\ : LocalMux
    port map (
            O => \N__41505\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__9270\ : LocalMux
    port map (
            O => \N__41502\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__9269\ : CascadeMux
    port map (
            O => \N__41495\,
            I => \N__41492\
        );

    \I__9268\ : InMux
    port map (
            O => \N__41492\,
            I => \N__41489\
        );

    \I__9267\ : LocalMux
    port map (
            O => \N__41489\,
            I => \N__41484\
        );

    \I__9266\ : InMux
    port map (
            O => \N__41488\,
            I => \N__41479\
        );

    \I__9265\ : InMux
    port map (
            O => \N__41487\,
            I => \N__41479\
        );

    \I__9264\ : Span12Mux_v
    port map (
            O => \N__41484\,
            I => \N__41474\
        );

    \I__9263\ : LocalMux
    port map (
            O => \N__41479\,
            I => \N__41474\
        );

    \I__9262\ : Odrv12
    port map (
            O => \N__41474\,
            I => \delay_measurement_inst.elapsed_time_hc_11\
        );

    \I__9261\ : InMux
    port map (
            O => \N__41471\,
            I => \bfn_17_9_0_\
        );

    \I__9260\ : CascadeMux
    port map (
            O => \N__41468\,
            I => \N__41463\
        );

    \I__9259\ : InMux
    port map (
            O => \N__41467\,
            I => \N__41460\
        );

    \I__9258\ : InMux
    port map (
            O => \N__41466\,
            I => \N__41457\
        );

    \I__9257\ : InMux
    port map (
            O => \N__41463\,
            I => \N__41454\
        );

    \I__9256\ : LocalMux
    port map (
            O => \N__41460\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__9255\ : LocalMux
    port map (
            O => \N__41457\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__9254\ : LocalMux
    port map (
            O => \N__41454\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__9253\ : InMux
    port map (
            O => \N__41447\,
            I => \N__41443\
        );

    \I__9252\ : CascadeMux
    port map (
            O => \N__41446\,
            I => \N__41439\
        );

    \I__9251\ : LocalMux
    port map (
            O => \N__41443\,
            I => \N__41436\
        );

    \I__9250\ : InMux
    port map (
            O => \N__41442\,
            I => \N__41431\
        );

    \I__9249\ : InMux
    port map (
            O => \N__41439\,
            I => \N__41431\
        );

    \I__9248\ : Span4Mux_v
    port map (
            O => \N__41436\,
            I => \N__41428\
        );

    \I__9247\ : LocalMux
    port map (
            O => \N__41431\,
            I => \N__41425\
        );

    \I__9246\ : Odrv4
    port map (
            O => \N__41428\,
            I => \delay_measurement_inst.elapsed_time_hc_12\
        );

    \I__9245\ : Odrv12
    port map (
            O => \N__41425\,
            I => \delay_measurement_inst.elapsed_time_hc_12\
        );

    \I__9244\ : InMux
    port map (
            O => \N__41420\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__9243\ : CascadeMux
    port map (
            O => \N__41417\,
            I => \N__41412\
        );

    \I__9242\ : InMux
    port map (
            O => \N__41416\,
            I => \N__41409\
        );

    \I__9241\ : InMux
    port map (
            O => \N__41415\,
            I => \N__41406\
        );

    \I__9240\ : InMux
    port map (
            O => \N__41412\,
            I => \N__41403\
        );

    \I__9239\ : LocalMux
    port map (
            O => \N__41409\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__9238\ : LocalMux
    port map (
            O => \N__41406\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__9237\ : LocalMux
    port map (
            O => \N__41403\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__9236\ : CascadeMux
    port map (
            O => \N__41396\,
            I => \N__41392\
        );

    \I__9235\ : CascadeMux
    port map (
            O => \N__41395\,
            I => \N__41388\
        );

    \I__9234\ : InMux
    port map (
            O => \N__41392\,
            I => \N__41385\
        );

    \I__9233\ : InMux
    port map (
            O => \N__41391\,
            I => \N__41380\
        );

    \I__9232\ : InMux
    port map (
            O => \N__41388\,
            I => \N__41380\
        );

    \I__9231\ : LocalMux
    port map (
            O => \N__41385\,
            I => \N__41377\
        );

    \I__9230\ : LocalMux
    port map (
            O => \N__41380\,
            I => \N__41374\
        );

    \I__9229\ : Span4Mux_h
    port map (
            O => \N__41377\,
            I => \N__41369\
        );

    \I__9228\ : Span4Mux_h
    port map (
            O => \N__41374\,
            I => \N__41369\
        );

    \I__9227\ : Odrv4
    port map (
            O => \N__41369\,
            I => \delay_measurement_inst.elapsed_time_hc_13\
        );

    \I__9226\ : InMux
    port map (
            O => \N__41366\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__9225\ : CascadeMux
    port map (
            O => \N__41363\,
            I => \N__41358\
        );

    \I__9224\ : InMux
    port map (
            O => \N__41362\,
            I => \N__41355\
        );

    \I__9223\ : InMux
    port map (
            O => \N__41361\,
            I => \N__41352\
        );

    \I__9222\ : InMux
    port map (
            O => \N__41358\,
            I => \N__41349\
        );

    \I__9221\ : LocalMux
    port map (
            O => \N__41355\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__9220\ : LocalMux
    port map (
            O => \N__41352\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__9219\ : LocalMux
    port map (
            O => \N__41349\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__9218\ : InMux
    port map (
            O => \N__41342\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__9217\ : CascadeMux
    port map (
            O => \N__41339\,
            I => \N__41336\
        );

    \I__9216\ : InMux
    port map (
            O => \N__41336\,
            I => \N__41333\
        );

    \I__9215\ : LocalMux
    port map (
            O => \N__41333\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\
        );

    \I__9214\ : CascadeMux
    port map (
            O => \N__41330\,
            I => \N__41327\
        );

    \I__9213\ : InMux
    port map (
            O => \N__41327\,
            I => \N__41324\
        );

    \I__9212\ : LocalMux
    port map (
            O => \N__41324\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\
        );

    \I__9211\ : CascadeMux
    port map (
            O => \N__41321\,
            I => \N__41318\
        );

    \I__9210\ : InMux
    port map (
            O => \N__41318\,
            I => \N__41315\
        );

    \I__9209\ : LocalMux
    port map (
            O => \N__41315\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\
        );

    \I__9208\ : InMux
    port map (
            O => \N__41312\,
            I => \N__41308\
        );

    \I__9207\ : InMux
    port map (
            O => \N__41311\,
            I => \N__41305\
        );

    \I__9206\ : LocalMux
    port map (
            O => \N__41308\,
            I => \N__41301\
        );

    \I__9205\ : LocalMux
    port map (
            O => \N__41305\,
            I => \N__41298\
        );

    \I__9204\ : InMux
    port map (
            O => \N__41304\,
            I => \N__41295\
        );

    \I__9203\ : Odrv12
    port map (
            O => \N__41301\,
            I => measured_delay_tr_12
        );

    \I__9202\ : Odrv4
    port map (
            O => \N__41298\,
            I => measured_delay_tr_12
        );

    \I__9201\ : LocalMux
    port map (
            O => \N__41295\,
            I => measured_delay_tr_12
        );

    \I__9200\ : CascadeMux
    port map (
            O => \N__41288\,
            I => \N__41285\
        );

    \I__9199\ : InMux
    port map (
            O => \N__41285\,
            I => \N__41282\
        );

    \I__9198\ : LocalMux
    port map (
            O => \N__41282\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\
        );

    \I__9197\ : InMux
    port map (
            O => \N__41279\,
            I => \N__41276\
        );

    \I__9196\ : LocalMux
    port map (
            O => \N__41276\,
            I => \N__41273\
        );

    \I__9195\ : Span4Mux_v
    port map (
            O => \N__41273\,
            I => \N__41269\
        );

    \I__9194\ : InMux
    port map (
            O => \N__41272\,
            I => \N__41266\
        );

    \I__9193\ : Span4Mux_h
    port map (
            O => \N__41269\,
            I => \N__41263\
        );

    \I__9192\ : LocalMux
    port map (
            O => \N__41266\,
            I => \N__41260\
        );

    \I__9191\ : Span4Mux_h
    port map (
            O => \N__41263\,
            I => \N__41257\
        );

    \I__9190\ : Span4Mux_v
    port map (
            O => \N__41260\,
            I => \N__41254\
        );

    \I__9189\ : Odrv4
    port map (
            O => \N__41257\,
            I => \delay_measurement_inst.elapsed_time_hc_1\
        );

    \I__9188\ : Odrv4
    port map (
            O => \N__41254\,
            I => \delay_measurement_inst.elapsed_time_hc_1\
        );

    \I__9187\ : InMux
    port map (
            O => \N__41249\,
            I => \N__41244\
        );

    \I__9186\ : InMux
    port map (
            O => \N__41248\,
            I => \N__41241\
        );

    \I__9185\ : InMux
    port map (
            O => \N__41247\,
            I => \N__41238\
        );

    \I__9184\ : LocalMux
    port map (
            O => \N__41244\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__9183\ : LocalMux
    port map (
            O => \N__41241\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__9182\ : LocalMux
    port map (
            O => \N__41238\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__9181\ : InMux
    port map (
            O => \N__41231\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__9180\ : CascadeMux
    port map (
            O => \N__41228\,
            I => \N__41223\
        );

    \I__9179\ : InMux
    port map (
            O => \N__41227\,
            I => \N__41220\
        );

    \I__9178\ : InMux
    port map (
            O => \N__41226\,
            I => \N__41217\
        );

    \I__9177\ : InMux
    port map (
            O => \N__41223\,
            I => \N__41214\
        );

    \I__9176\ : LocalMux
    port map (
            O => \N__41220\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__9175\ : LocalMux
    port map (
            O => \N__41217\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__9174\ : LocalMux
    port map (
            O => \N__41214\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__9173\ : InMux
    port map (
            O => \N__41207\,
            I => \N__41202\
        );

    \I__9172\ : InMux
    port map (
            O => \N__41206\,
            I => \N__41199\
        );

    \I__9171\ : InMux
    port map (
            O => \N__41205\,
            I => \N__41196\
        );

    \I__9170\ : LocalMux
    port map (
            O => \N__41202\,
            I => \N__41193\
        );

    \I__9169\ : LocalMux
    port map (
            O => \N__41199\,
            I => \N__41190\
        );

    \I__9168\ : LocalMux
    port map (
            O => \N__41196\,
            I => \N__41187\
        );

    \I__9167\ : Span4Mux_h
    port map (
            O => \N__41193\,
            I => \N__41184\
        );

    \I__9166\ : Span4Mux_h
    port map (
            O => \N__41190\,
            I => \N__41181\
        );

    \I__9165\ : Odrv4
    port map (
            O => \N__41187\,
            I => \delay_measurement_inst.elapsed_time_hc_5\
        );

    \I__9164\ : Odrv4
    port map (
            O => \N__41184\,
            I => \delay_measurement_inst.elapsed_time_hc_5\
        );

    \I__9163\ : Odrv4
    port map (
            O => \N__41181\,
            I => \delay_measurement_inst.elapsed_time_hc_5\
        );

    \I__9162\ : InMux
    port map (
            O => \N__41174\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__9161\ : CascadeMux
    port map (
            O => \N__41171\,
            I => \N__41166\
        );

    \I__9160\ : InMux
    port map (
            O => \N__41170\,
            I => \N__41163\
        );

    \I__9159\ : InMux
    port map (
            O => \N__41169\,
            I => \N__41160\
        );

    \I__9158\ : InMux
    port map (
            O => \N__41166\,
            I => \N__41157\
        );

    \I__9157\ : LocalMux
    port map (
            O => \N__41163\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__9156\ : LocalMux
    port map (
            O => \N__41160\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__9155\ : LocalMux
    port map (
            O => \N__41157\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__9154\ : InMux
    port map (
            O => \N__41150\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__9153\ : InMux
    port map (
            O => \N__41147\,
            I => \N__41144\
        );

    \I__9152\ : LocalMux
    port map (
            O => \N__41144\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\
        );

    \I__9151\ : CascadeMux
    port map (
            O => \N__41141\,
            I => \N__41138\
        );

    \I__9150\ : InMux
    port map (
            O => \N__41138\,
            I => \N__41135\
        );

    \I__9149\ : LocalMux
    port map (
            O => \N__41135\,
            I => \N__41132\
        );

    \I__9148\ : Odrv4
    port map (
            O => \N__41132\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\
        );

    \I__9147\ : CascadeMux
    port map (
            O => \N__41129\,
            I => \N__41126\
        );

    \I__9146\ : InMux
    port map (
            O => \N__41126\,
            I => \N__41123\
        );

    \I__9145\ : LocalMux
    port map (
            O => \N__41123\,
            I => \N__41120\
        );

    \I__9144\ : Span4Mux_h
    port map (
            O => \N__41120\,
            I => \N__41117\
        );

    \I__9143\ : Odrv4
    port map (
            O => \N__41117\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\
        );

    \I__9142\ : CascadeMux
    port map (
            O => \N__41114\,
            I => \N__41111\
        );

    \I__9141\ : InMux
    port map (
            O => \N__41111\,
            I => \N__41108\
        );

    \I__9140\ : LocalMux
    port map (
            O => \N__41108\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\
        );

    \I__9139\ : CascadeMux
    port map (
            O => \N__41105\,
            I => \N__41102\
        );

    \I__9138\ : InMux
    port map (
            O => \N__41102\,
            I => \N__41099\
        );

    \I__9137\ : LocalMux
    port map (
            O => \N__41099\,
            I => \N__41096\
        );

    \I__9136\ : Span4Mux_v
    port map (
            O => \N__41096\,
            I => \N__41093\
        );

    \I__9135\ : Odrv4
    port map (
            O => \N__41093\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\
        );

    \I__9134\ : CascadeMux
    port map (
            O => \N__41090\,
            I => \N__41087\
        );

    \I__9133\ : InMux
    port map (
            O => \N__41087\,
            I => \N__41084\
        );

    \I__9132\ : LocalMux
    port map (
            O => \N__41084\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\
        );

    \I__9131\ : InMux
    port map (
            O => \N__41081\,
            I => \N__41077\
        );

    \I__9130\ : InMux
    port map (
            O => \N__41080\,
            I => \N__41074\
        );

    \I__9129\ : LocalMux
    port map (
            O => \N__41077\,
            I => \N__41070\
        );

    \I__9128\ : LocalMux
    port map (
            O => \N__41074\,
            I => \N__41067\
        );

    \I__9127\ : InMux
    port map (
            O => \N__41073\,
            I => \N__41064\
        );

    \I__9126\ : Odrv12
    port map (
            O => \N__41070\,
            I => measured_delay_tr_10
        );

    \I__9125\ : Odrv4
    port map (
            O => \N__41067\,
            I => measured_delay_tr_10
        );

    \I__9124\ : LocalMux
    port map (
            O => \N__41064\,
            I => measured_delay_tr_10
        );

    \I__9123\ : CascadeMux
    port map (
            O => \N__41057\,
            I => \N__41054\
        );

    \I__9122\ : InMux
    port map (
            O => \N__41054\,
            I => \N__41051\
        );

    \I__9121\ : LocalMux
    port map (
            O => \N__41051\,
            I => \N__41048\
        );

    \I__9120\ : Odrv4
    port map (
            O => \N__41048\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\
        );

    \I__9119\ : CascadeMux
    port map (
            O => \N__41045\,
            I => \N__41042\
        );

    \I__9118\ : InMux
    port map (
            O => \N__41042\,
            I => \N__41039\
        );

    \I__9117\ : LocalMux
    port map (
            O => \N__41039\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\
        );

    \I__9116\ : CascadeMux
    port map (
            O => \N__41036\,
            I => \N__41033\
        );

    \I__9115\ : InMux
    port map (
            O => \N__41033\,
            I => \N__41030\
        );

    \I__9114\ : LocalMux
    port map (
            O => \N__41030\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\
        );

    \I__9113\ : InMux
    port map (
            O => \N__41027\,
            I => \N__41023\
        );

    \I__9112\ : InMux
    port map (
            O => \N__41026\,
            I => \N__41020\
        );

    \I__9111\ : LocalMux
    port map (
            O => \N__41023\,
            I => \N__41014\
        );

    \I__9110\ : LocalMux
    port map (
            O => \N__41020\,
            I => \N__41014\
        );

    \I__9109\ : InMux
    port map (
            O => \N__41019\,
            I => \N__41011\
        );

    \I__9108\ : Odrv12
    port map (
            O => \N__41014\,
            I => measured_delay_tr_9
        );

    \I__9107\ : LocalMux
    port map (
            O => \N__41011\,
            I => measured_delay_tr_9
        );

    \I__9106\ : CascadeMux
    port map (
            O => \N__41006\,
            I => \N__41003\
        );

    \I__9105\ : InMux
    port map (
            O => \N__41003\,
            I => \N__41000\
        );

    \I__9104\ : LocalMux
    port map (
            O => \N__41000\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_3\
        );

    \I__9103\ : CascadeMux
    port map (
            O => \N__40997\,
            I => \N__40994\
        );

    \I__9102\ : InMux
    port map (
            O => \N__40994\,
            I => \N__40991\
        );

    \I__9101\ : LocalMux
    port map (
            O => \N__40991\,
            I => \N__40988\
        );

    \I__9100\ : Odrv4
    port map (
            O => \N__40988\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_5\
        );

    \I__9099\ : CascadeMux
    port map (
            O => \N__40985\,
            I => \N__40982\
        );

    \I__9098\ : InMux
    port map (
            O => \N__40982\,
            I => \N__40979\
        );

    \I__9097\ : LocalMux
    port map (
            O => \N__40979\,
            I => \N__40976\
        );

    \I__9096\ : Odrv4
    port map (
            O => \N__40976\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_10\
        );

    \I__9095\ : CascadeMux
    port map (
            O => \N__40973\,
            I => \N__40970\
        );

    \I__9094\ : InMux
    port map (
            O => \N__40970\,
            I => \N__40967\
        );

    \I__9093\ : LocalMux
    port map (
            O => \N__40967\,
            I => \N__40964\
        );

    \I__9092\ : Span4Mux_h
    port map (
            O => \N__40964\,
            I => \N__40961\
        );

    \I__9091\ : Odrv4
    port map (
            O => \N__40961\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_11\
        );

    \I__9090\ : CascadeMux
    port map (
            O => \N__40958\,
            I => \N__40955\
        );

    \I__9089\ : InMux
    port map (
            O => \N__40955\,
            I => \N__40952\
        );

    \I__9088\ : LocalMux
    port map (
            O => \N__40952\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_13\
        );

    \I__9087\ : CascadeMux
    port map (
            O => \N__40949\,
            I => \N__40946\
        );

    \I__9086\ : InMux
    port map (
            O => \N__40946\,
            I => \N__40943\
        );

    \I__9085\ : LocalMux
    port map (
            O => \N__40943\,
            I => \N__40940\
        );

    \I__9084\ : Odrv4
    port map (
            O => \N__40940\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_12\
        );

    \I__9083\ : CascadeMux
    port map (
            O => \N__40937\,
            I => \N__40934\
        );

    \I__9082\ : InMux
    port map (
            O => \N__40934\,
            I => \N__40931\
        );

    \I__9081\ : LocalMux
    port map (
            O => \N__40931\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_9\
        );

    \I__9080\ : CascadeMux
    port map (
            O => \N__40928\,
            I => \N__40925\
        );

    \I__9079\ : InMux
    port map (
            O => \N__40925\,
            I => \N__40922\
        );

    \I__9078\ : LocalMux
    port map (
            O => \N__40922\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_19\
        );

    \I__9077\ : InMux
    port map (
            O => \N__40919\,
            I => \N__40916\
        );

    \I__9076\ : LocalMux
    port map (
            O => \N__40916\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\
        );

    \I__9075\ : CascadeMux
    port map (
            O => \N__40913\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6_cascade_\
        );

    \I__9074\ : CascadeMux
    port map (
            O => \N__40910\,
            I => \N__40907\
        );

    \I__9073\ : InMux
    port map (
            O => \N__40907\,
            I => \N__40904\
        );

    \I__9072\ : LocalMux
    port map (
            O => \N__40904\,
            I => \N__40901\
        );

    \I__9071\ : Odrv4
    port map (
            O => \N__40901\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_2\
        );

    \I__9070\ : InMux
    port map (
            O => \N__40898\,
            I => \N__40895\
        );

    \I__9069\ : LocalMux
    port map (
            O => \N__40895\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_15\
        );

    \I__9068\ : CascadeMux
    port map (
            O => \N__40892\,
            I => \N__40889\
        );

    \I__9067\ : InMux
    port map (
            O => \N__40889\,
            I => \N__40886\
        );

    \I__9066\ : LocalMux
    port map (
            O => \N__40886\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_1\
        );

    \I__9065\ : CascadeMux
    port map (
            O => \N__40883\,
            I => \N__40880\
        );

    \I__9064\ : InMux
    port map (
            O => \N__40880\,
            I => \N__40877\
        );

    \I__9063\ : LocalMux
    port map (
            O => \N__40877\,
            I => \N__40874\
        );

    \I__9062\ : Odrv4
    port map (
            O => \N__40874\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_6\
        );

    \I__9061\ : CascadeMux
    port map (
            O => \N__40871\,
            I => \N__40868\
        );

    \I__9060\ : InMux
    port map (
            O => \N__40868\,
            I => \N__40865\
        );

    \I__9059\ : LocalMux
    port map (
            O => \N__40865\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_7\
        );

    \I__9058\ : CascadeMux
    port map (
            O => \N__40862\,
            I => \N__40859\
        );

    \I__9057\ : InMux
    port map (
            O => \N__40859\,
            I => \N__40856\
        );

    \I__9056\ : LocalMux
    port map (
            O => \N__40856\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_4\
        );

    \I__9055\ : InMux
    port map (
            O => \N__40853\,
            I => \N__40839\
        );

    \I__9054\ : InMux
    port map (
            O => \N__40852\,
            I => \N__40832\
        );

    \I__9053\ : InMux
    port map (
            O => \N__40851\,
            I => \N__40832\
        );

    \I__9052\ : InMux
    port map (
            O => \N__40850\,
            I => \N__40832\
        );

    \I__9051\ : InMux
    port map (
            O => \N__40849\,
            I => \N__40822\
        );

    \I__9050\ : InMux
    port map (
            O => \N__40848\,
            I => \N__40822\
        );

    \I__9049\ : InMux
    port map (
            O => \N__40847\,
            I => \N__40822\
        );

    \I__9048\ : InMux
    port map (
            O => \N__40846\,
            I => \N__40822\
        );

    \I__9047\ : InMux
    port map (
            O => \N__40845\,
            I => \N__40817\
        );

    \I__9046\ : InMux
    port map (
            O => \N__40844\,
            I => \N__40817\
        );

    \I__9045\ : InMux
    port map (
            O => \N__40843\,
            I => \N__40812\
        );

    \I__9044\ : InMux
    port map (
            O => \N__40842\,
            I => \N__40812\
        );

    \I__9043\ : LocalMux
    port map (
            O => \N__40839\,
            I => \N__40809\
        );

    \I__9042\ : LocalMux
    port map (
            O => \N__40832\,
            I => \N__40806\
        );

    \I__9041\ : InMux
    port map (
            O => \N__40831\,
            I => \N__40803\
        );

    \I__9040\ : LocalMux
    port map (
            O => \N__40822\,
            I => \N__40800\
        );

    \I__9039\ : LocalMux
    port map (
            O => \N__40817\,
            I => \N__40795\
        );

    \I__9038\ : LocalMux
    port map (
            O => \N__40812\,
            I => \N__40795\
        );

    \I__9037\ : Span4Mux_v
    port map (
            O => \N__40809\,
            I => \N__40781\
        );

    \I__9036\ : Span4Mux_h
    port map (
            O => \N__40806\,
            I => \N__40778\
        );

    \I__9035\ : LocalMux
    port map (
            O => \N__40803\,
            I => \N__40775\
        );

    \I__9034\ : Span4Mux_h
    port map (
            O => \N__40800\,
            I => \N__40772\
        );

    \I__9033\ : Span4Mux_h
    port map (
            O => \N__40795\,
            I => \N__40769\
        );

    \I__9032\ : InMux
    port map (
            O => \N__40794\,
            I => \N__40762\
        );

    \I__9031\ : InMux
    port map (
            O => \N__40793\,
            I => \N__40762\
        );

    \I__9030\ : InMux
    port map (
            O => \N__40792\,
            I => \N__40762\
        );

    \I__9029\ : InMux
    port map (
            O => \N__40791\,
            I => \N__40745\
        );

    \I__9028\ : InMux
    port map (
            O => \N__40790\,
            I => \N__40745\
        );

    \I__9027\ : InMux
    port map (
            O => \N__40789\,
            I => \N__40745\
        );

    \I__9026\ : InMux
    port map (
            O => \N__40788\,
            I => \N__40745\
        );

    \I__9025\ : InMux
    port map (
            O => \N__40787\,
            I => \N__40745\
        );

    \I__9024\ : InMux
    port map (
            O => \N__40786\,
            I => \N__40745\
        );

    \I__9023\ : InMux
    port map (
            O => \N__40785\,
            I => \N__40745\
        );

    \I__9022\ : InMux
    port map (
            O => \N__40784\,
            I => \N__40745\
        );

    \I__9021\ : Odrv4
    port map (
            O => \N__40781\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__9020\ : Odrv4
    port map (
            O => \N__40778\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__9019\ : Odrv12
    port map (
            O => \N__40775\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__9018\ : Odrv4
    port map (
            O => \N__40772\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__9017\ : Odrv4
    port map (
            O => \N__40769\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__9016\ : LocalMux
    port map (
            O => \N__40762\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__9015\ : LocalMux
    port map (
            O => \N__40745\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__9014\ : CascadeMux
    port map (
            O => \N__40730\,
            I => \N__40725\
        );

    \I__9013\ : CascadeMux
    port map (
            O => \N__40729\,
            I => \N__40713\
        );

    \I__9012\ : CascadeMux
    port map (
            O => \N__40728\,
            I => \N__40710\
        );

    \I__9011\ : InMux
    port map (
            O => \N__40725\,
            I => \N__40706\
        );

    \I__9010\ : InMux
    port map (
            O => \N__40724\,
            I => \N__40703\
        );

    \I__9009\ : InMux
    port map (
            O => \N__40723\,
            I => \N__40688\
        );

    \I__9008\ : InMux
    port map (
            O => \N__40722\,
            I => \N__40688\
        );

    \I__9007\ : CascadeMux
    port map (
            O => \N__40721\,
            I => \N__40685\
        );

    \I__9006\ : InMux
    port map (
            O => \N__40720\,
            I => \N__40672\
        );

    \I__9005\ : InMux
    port map (
            O => \N__40719\,
            I => \N__40672\
        );

    \I__9004\ : InMux
    port map (
            O => \N__40718\,
            I => \N__40672\
        );

    \I__9003\ : InMux
    port map (
            O => \N__40717\,
            I => \N__40672\
        );

    \I__9002\ : CascadeMux
    port map (
            O => \N__40716\,
            I => \N__40667\
        );

    \I__9001\ : InMux
    port map (
            O => \N__40713\,
            I => \N__40659\
        );

    \I__9000\ : InMux
    port map (
            O => \N__40710\,
            I => \N__40659\
        );

    \I__8999\ : InMux
    port map (
            O => \N__40709\,
            I => \N__40659\
        );

    \I__8998\ : LocalMux
    port map (
            O => \N__40706\,
            I => \N__40654\
        );

    \I__8997\ : LocalMux
    port map (
            O => \N__40703\,
            I => \N__40654\
        );

    \I__8996\ : InMux
    port map (
            O => \N__40702\,
            I => \N__40649\
        );

    \I__8995\ : InMux
    port map (
            O => \N__40701\,
            I => \N__40632\
        );

    \I__8994\ : InMux
    port map (
            O => \N__40700\,
            I => \N__40632\
        );

    \I__8993\ : InMux
    port map (
            O => \N__40699\,
            I => \N__40632\
        );

    \I__8992\ : InMux
    port map (
            O => \N__40698\,
            I => \N__40632\
        );

    \I__8991\ : InMux
    port map (
            O => \N__40697\,
            I => \N__40632\
        );

    \I__8990\ : InMux
    port map (
            O => \N__40696\,
            I => \N__40632\
        );

    \I__8989\ : InMux
    port map (
            O => \N__40695\,
            I => \N__40632\
        );

    \I__8988\ : InMux
    port map (
            O => \N__40694\,
            I => \N__40632\
        );

    \I__8987\ : InMux
    port map (
            O => \N__40693\,
            I => \N__40629\
        );

    \I__8986\ : LocalMux
    port map (
            O => \N__40688\,
            I => \N__40626\
        );

    \I__8985\ : InMux
    port map (
            O => \N__40685\,
            I => \N__40615\
        );

    \I__8984\ : InMux
    port map (
            O => \N__40684\,
            I => \N__40615\
        );

    \I__8983\ : InMux
    port map (
            O => \N__40683\,
            I => \N__40615\
        );

    \I__8982\ : InMux
    port map (
            O => \N__40682\,
            I => \N__40615\
        );

    \I__8981\ : InMux
    port map (
            O => \N__40681\,
            I => \N__40615\
        );

    \I__8980\ : LocalMux
    port map (
            O => \N__40672\,
            I => \N__40612\
        );

    \I__8979\ : InMux
    port map (
            O => \N__40671\,
            I => \N__40603\
        );

    \I__8978\ : InMux
    port map (
            O => \N__40670\,
            I => \N__40603\
        );

    \I__8977\ : InMux
    port map (
            O => \N__40667\,
            I => \N__40603\
        );

    \I__8976\ : InMux
    port map (
            O => \N__40666\,
            I => \N__40603\
        );

    \I__8975\ : LocalMux
    port map (
            O => \N__40659\,
            I => \N__40600\
        );

    \I__8974\ : Span4Mux_h
    port map (
            O => \N__40654\,
            I => \N__40597\
        );

    \I__8973\ : InMux
    port map (
            O => \N__40653\,
            I => \N__40592\
        );

    \I__8972\ : InMux
    port map (
            O => \N__40652\,
            I => \N__40592\
        );

    \I__8971\ : LocalMux
    port map (
            O => \N__40649\,
            I => \N__40587\
        );

    \I__8970\ : LocalMux
    port map (
            O => \N__40632\,
            I => \N__40587\
        );

    \I__8969\ : LocalMux
    port map (
            O => \N__40629\,
            I => \N__40582\
        );

    \I__8968\ : Span4Mux_h
    port map (
            O => \N__40626\,
            I => \N__40582\
        );

    \I__8967\ : LocalMux
    port map (
            O => \N__40615\,
            I => \N__40577\
        );

    \I__8966\ : Span4Mux_h
    port map (
            O => \N__40612\,
            I => \N__40577\
        );

    \I__8965\ : LocalMux
    port map (
            O => \N__40603\,
            I => \N__40570\
        );

    \I__8964\ : Span4Mux_h
    port map (
            O => \N__40600\,
            I => \N__40570\
        );

    \I__8963\ : Span4Mux_h
    port map (
            O => \N__40597\,
            I => \N__40570\
        );

    \I__8962\ : LocalMux
    port map (
            O => \N__40592\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__8961\ : Odrv4
    port map (
            O => \N__40587\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__8960\ : Odrv4
    port map (
            O => \N__40582\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__8959\ : Odrv4
    port map (
            O => \N__40577\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__8958\ : Odrv4
    port map (
            O => \N__40570\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__8957\ : CascadeMux
    port map (
            O => \N__40559\,
            I => \N__40555\
        );

    \I__8956\ : CascadeMux
    port map (
            O => \N__40558\,
            I => \N__40548\
        );

    \I__8955\ : InMux
    port map (
            O => \N__40555\,
            I => \N__40541\
        );

    \I__8954\ : InMux
    port map (
            O => \N__40554\,
            I => \N__40541\
        );

    \I__8953\ : CascadeMux
    port map (
            O => \N__40553\,
            I => \N__40538\
        );

    \I__8952\ : CascadeMux
    port map (
            O => \N__40552\,
            I => \N__40526\
        );

    \I__8951\ : CascadeMux
    port map (
            O => \N__40551\,
            I => \N__40521\
        );

    \I__8950\ : InMux
    port map (
            O => \N__40548\,
            I => \N__40512\
        );

    \I__8949\ : InMux
    port map (
            O => \N__40547\,
            I => \N__40512\
        );

    \I__8948\ : InMux
    port map (
            O => \N__40546\,
            I => \N__40512\
        );

    \I__8947\ : LocalMux
    port map (
            O => \N__40541\,
            I => \N__40506\
        );

    \I__8946\ : InMux
    port map (
            O => \N__40538\,
            I => \N__40503\
        );

    \I__8945\ : CascadeMux
    port map (
            O => \N__40537\,
            I => \N__40499\
        );

    \I__8944\ : CascadeMux
    port map (
            O => \N__40536\,
            I => \N__40493\
        );

    \I__8943\ : CascadeMux
    port map (
            O => \N__40535\,
            I => \N__40490\
        );

    \I__8942\ : CascadeMux
    port map (
            O => \N__40534\,
            I => \N__40482\
        );

    \I__8941\ : CascadeMux
    port map (
            O => \N__40533\,
            I => \N__40479\
        );

    \I__8940\ : CascadeMux
    port map (
            O => \N__40532\,
            I => \N__40472\
        );

    \I__8939\ : CascadeMux
    port map (
            O => \N__40531\,
            I => \N__40468\
        );

    \I__8938\ : CascadeMux
    port map (
            O => \N__40530\,
            I => \N__40465\
        );

    \I__8937\ : InMux
    port map (
            O => \N__40529\,
            I => \N__40458\
        );

    \I__8936\ : InMux
    port map (
            O => \N__40526\,
            I => \N__40445\
        );

    \I__8935\ : InMux
    port map (
            O => \N__40525\,
            I => \N__40445\
        );

    \I__8934\ : InMux
    port map (
            O => \N__40524\,
            I => \N__40445\
        );

    \I__8933\ : InMux
    port map (
            O => \N__40521\,
            I => \N__40445\
        );

    \I__8932\ : InMux
    port map (
            O => \N__40520\,
            I => \N__40445\
        );

    \I__8931\ : InMux
    port map (
            O => \N__40519\,
            I => \N__40445\
        );

    \I__8930\ : LocalMux
    port map (
            O => \N__40512\,
            I => \N__40442\
        );

    \I__8929\ : InMux
    port map (
            O => \N__40511\,
            I => \N__40437\
        );

    \I__8928\ : InMux
    port map (
            O => \N__40510\,
            I => \N__40437\
        );

    \I__8927\ : CascadeMux
    port map (
            O => \N__40509\,
            I => \N__40434\
        );

    \I__8926\ : Sp12to4
    port map (
            O => \N__40506\,
            I => \N__40429\
        );

    \I__8925\ : LocalMux
    port map (
            O => \N__40503\,
            I => \N__40429\
        );

    \I__8924\ : InMux
    port map (
            O => \N__40502\,
            I => \N__40418\
        );

    \I__8923\ : InMux
    port map (
            O => \N__40499\,
            I => \N__40418\
        );

    \I__8922\ : InMux
    port map (
            O => \N__40498\,
            I => \N__40418\
        );

    \I__8921\ : InMux
    port map (
            O => \N__40497\,
            I => \N__40418\
        );

    \I__8920\ : InMux
    port map (
            O => \N__40496\,
            I => \N__40418\
        );

    \I__8919\ : InMux
    port map (
            O => \N__40493\,
            I => \N__40407\
        );

    \I__8918\ : InMux
    port map (
            O => \N__40490\,
            I => \N__40407\
        );

    \I__8917\ : InMux
    port map (
            O => \N__40489\,
            I => \N__40407\
        );

    \I__8916\ : InMux
    port map (
            O => \N__40488\,
            I => \N__40407\
        );

    \I__8915\ : InMux
    port map (
            O => \N__40487\,
            I => \N__40407\
        );

    \I__8914\ : InMux
    port map (
            O => \N__40486\,
            I => \N__40390\
        );

    \I__8913\ : InMux
    port map (
            O => \N__40485\,
            I => \N__40390\
        );

    \I__8912\ : InMux
    port map (
            O => \N__40482\,
            I => \N__40390\
        );

    \I__8911\ : InMux
    port map (
            O => \N__40479\,
            I => \N__40390\
        );

    \I__8910\ : InMux
    port map (
            O => \N__40478\,
            I => \N__40390\
        );

    \I__8909\ : InMux
    port map (
            O => \N__40477\,
            I => \N__40390\
        );

    \I__8908\ : InMux
    port map (
            O => \N__40476\,
            I => \N__40390\
        );

    \I__8907\ : InMux
    port map (
            O => \N__40475\,
            I => \N__40390\
        );

    \I__8906\ : InMux
    port map (
            O => \N__40472\,
            I => \N__40385\
        );

    \I__8905\ : InMux
    port map (
            O => \N__40471\,
            I => \N__40385\
        );

    \I__8904\ : InMux
    port map (
            O => \N__40468\,
            I => \N__40374\
        );

    \I__8903\ : InMux
    port map (
            O => \N__40465\,
            I => \N__40374\
        );

    \I__8902\ : InMux
    port map (
            O => \N__40464\,
            I => \N__40374\
        );

    \I__8901\ : InMux
    port map (
            O => \N__40463\,
            I => \N__40374\
        );

    \I__8900\ : InMux
    port map (
            O => \N__40462\,
            I => \N__40374\
        );

    \I__8899\ : InMux
    port map (
            O => \N__40461\,
            I => \N__40371\
        );

    \I__8898\ : LocalMux
    port map (
            O => \N__40458\,
            I => \N__40362\
        );

    \I__8897\ : LocalMux
    port map (
            O => \N__40445\,
            I => \N__40362\
        );

    \I__8896\ : Span4Mux_v
    port map (
            O => \N__40442\,
            I => \N__40362\
        );

    \I__8895\ : LocalMux
    port map (
            O => \N__40437\,
            I => \N__40362\
        );

    \I__8894\ : InMux
    port map (
            O => \N__40434\,
            I => \N__40359\
        );

    \I__8893\ : Span12Mux_s4_h
    port map (
            O => \N__40429\,
            I => \N__40355\
        );

    \I__8892\ : LocalMux
    port map (
            O => \N__40418\,
            I => \N__40346\
        );

    \I__8891\ : LocalMux
    port map (
            O => \N__40407\,
            I => \N__40346\
        );

    \I__8890\ : LocalMux
    port map (
            O => \N__40390\,
            I => \N__40346\
        );

    \I__8889\ : LocalMux
    port map (
            O => \N__40385\,
            I => \N__40346\
        );

    \I__8888\ : LocalMux
    port map (
            O => \N__40374\,
            I => \N__40343\
        );

    \I__8887\ : LocalMux
    port map (
            O => \N__40371\,
            I => \N__40340\
        );

    \I__8886\ : Span4Mux_v
    port map (
            O => \N__40362\,
            I => \N__40335\
        );

    \I__8885\ : LocalMux
    port map (
            O => \N__40359\,
            I => \N__40335\
        );

    \I__8884\ : InMux
    port map (
            O => \N__40358\,
            I => \N__40332\
        );

    \I__8883\ : Span12Mux_h
    port map (
            O => \N__40355\,
            I => \N__40329\
        );

    \I__8882\ : Span4Mux_v
    port map (
            O => \N__40346\,
            I => \N__40326\
        );

    \I__8881\ : Span4Mux_h
    port map (
            O => \N__40343\,
            I => \N__40323\
        );

    \I__8880\ : Span4Mux_h
    port map (
            O => \N__40340\,
            I => \N__40318\
        );

    \I__8879\ : Span4Mux_h
    port map (
            O => \N__40335\,
            I => \N__40318\
        );

    \I__8878\ : LocalMux
    port map (
            O => \N__40332\,
            I => measured_delay_hc_31
        );

    \I__8877\ : Odrv12
    port map (
            O => \N__40329\,
            I => measured_delay_hc_31
        );

    \I__8876\ : Odrv4
    port map (
            O => \N__40326\,
            I => measured_delay_hc_31
        );

    \I__8875\ : Odrv4
    port map (
            O => \N__40323\,
            I => measured_delay_hc_31
        );

    \I__8874\ : Odrv4
    port map (
            O => \N__40318\,
            I => measured_delay_hc_31
        );

    \I__8873\ : InMux
    port map (
            O => \N__40307\,
            I => \N__40304\
        );

    \I__8872\ : LocalMux
    port map (
            O => \N__40304\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10\
        );

    \I__8871\ : InMux
    port map (
            O => \N__40301\,
            I => \N__40297\
        );

    \I__8870\ : InMux
    port map (
            O => \N__40300\,
            I => \N__40294\
        );

    \I__8869\ : LocalMux
    port map (
            O => \N__40297\,
            I => \N__40291\
        );

    \I__8868\ : LocalMux
    port map (
            O => \N__40294\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__8867\ : Odrv12
    port map (
            O => \N__40291\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__8866\ : InMux
    port map (
            O => \N__40286\,
            I => \N__40283\
        );

    \I__8865\ : LocalMux
    port map (
            O => \N__40283\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13\
        );

    \I__8864\ : InMux
    port map (
            O => \N__40280\,
            I => \N__40276\
        );

    \I__8863\ : InMux
    port map (
            O => \N__40279\,
            I => \N__40273\
        );

    \I__8862\ : LocalMux
    port map (
            O => \N__40276\,
            I => \N__40270\
        );

    \I__8861\ : LocalMux
    port map (
            O => \N__40273\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__8860\ : Odrv4
    port map (
            O => \N__40270\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__8859\ : InMux
    port map (
            O => \N__40265\,
            I => \N__40262\
        );

    \I__8858\ : LocalMux
    port map (
            O => \N__40262\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15\
        );

    \I__8857\ : InMux
    port map (
            O => \N__40259\,
            I => \N__40255\
        );

    \I__8856\ : InMux
    port map (
            O => \N__40258\,
            I => \N__40252\
        );

    \I__8855\ : LocalMux
    port map (
            O => \N__40255\,
            I => \N__40249\
        );

    \I__8854\ : LocalMux
    port map (
            O => \N__40252\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__8853\ : Odrv12
    port map (
            O => \N__40249\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__8852\ : InMux
    port map (
            O => \N__40244\,
            I => \N__40220\
        );

    \I__8851\ : InMux
    port map (
            O => \N__40243\,
            I => \N__40220\
        );

    \I__8850\ : InMux
    port map (
            O => \N__40242\,
            I => \N__40220\
        );

    \I__8849\ : InMux
    port map (
            O => \N__40241\,
            I => \N__40220\
        );

    \I__8848\ : InMux
    port map (
            O => \N__40240\,
            I => \N__40203\
        );

    \I__8847\ : InMux
    port map (
            O => \N__40239\,
            I => \N__40203\
        );

    \I__8846\ : InMux
    port map (
            O => \N__40238\,
            I => \N__40203\
        );

    \I__8845\ : InMux
    port map (
            O => \N__40237\,
            I => \N__40203\
        );

    \I__8844\ : InMux
    port map (
            O => \N__40236\,
            I => \N__40203\
        );

    \I__8843\ : InMux
    port map (
            O => \N__40235\,
            I => \N__40203\
        );

    \I__8842\ : InMux
    port map (
            O => \N__40234\,
            I => \N__40203\
        );

    \I__8841\ : InMux
    port map (
            O => \N__40233\,
            I => \N__40203\
        );

    \I__8840\ : InMux
    port map (
            O => \N__40232\,
            I => \N__40194\
        );

    \I__8839\ : InMux
    port map (
            O => \N__40231\,
            I => \N__40188\
        );

    \I__8838\ : InMux
    port map (
            O => \N__40230\,
            I => \N__40188\
        );

    \I__8837\ : CascadeMux
    port map (
            O => \N__40229\,
            I => \N__40185\
        );

    \I__8836\ : LocalMux
    port map (
            O => \N__40220\,
            I => \N__40179\
        );

    \I__8835\ : LocalMux
    port map (
            O => \N__40203\,
            I => \N__40179\
        );

    \I__8834\ : InMux
    port map (
            O => \N__40202\,
            I => \N__40176\
        );

    \I__8833\ : InMux
    port map (
            O => \N__40201\,
            I => \N__40165\
        );

    \I__8832\ : InMux
    port map (
            O => \N__40200\,
            I => \N__40165\
        );

    \I__8831\ : InMux
    port map (
            O => \N__40199\,
            I => \N__40165\
        );

    \I__8830\ : InMux
    port map (
            O => \N__40198\,
            I => \N__40165\
        );

    \I__8829\ : InMux
    port map (
            O => \N__40197\,
            I => \N__40165\
        );

    \I__8828\ : LocalMux
    port map (
            O => \N__40194\,
            I => \N__40162\
        );

    \I__8827\ : InMux
    port map (
            O => \N__40193\,
            I => \N__40159\
        );

    \I__8826\ : LocalMux
    port map (
            O => \N__40188\,
            I => \N__40156\
        );

    \I__8825\ : InMux
    port map (
            O => \N__40185\,
            I => \N__40151\
        );

    \I__8824\ : InMux
    port map (
            O => \N__40184\,
            I => \N__40151\
        );

    \I__8823\ : Span4Mux_h
    port map (
            O => \N__40179\,
            I => \N__40148\
        );

    \I__8822\ : LocalMux
    port map (
            O => \N__40176\,
            I => \N__40145\
        );

    \I__8821\ : LocalMux
    port map (
            O => \N__40165\,
            I => \N__40136\
        );

    \I__8820\ : Span4Mux_v
    port map (
            O => \N__40162\,
            I => \N__40136\
        );

    \I__8819\ : LocalMux
    port map (
            O => \N__40159\,
            I => \N__40136\
        );

    \I__8818\ : Span4Mux_h
    port map (
            O => \N__40156\,
            I => \N__40136\
        );

    \I__8817\ : LocalMux
    port map (
            O => \N__40151\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__8816\ : Odrv4
    port map (
            O => \N__40148\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__8815\ : Odrv12
    port map (
            O => \N__40145\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__8814\ : Odrv4
    port map (
            O => \N__40136\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__8813\ : CascadeMux
    port map (
            O => \N__40127\,
            I => \N__40117\
        );

    \I__8812\ : CascadeMux
    port map (
            O => \N__40126\,
            I => \N__40110\
        );

    \I__8811\ : CascadeMux
    port map (
            O => \N__40125\,
            I => \N__40107\
        );

    \I__8810\ : CascadeMux
    port map (
            O => \N__40124\,
            I => \N__40104\
        );

    \I__8809\ : CascadeMux
    port map (
            O => \N__40123\,
            I => \N__40101\
        );

    \I__8808\ : CascadeMux
    port map (
            O => \N__40122\,
            I => \N__40097\
        );

    \I__8807\ : CascadeMux
    port map (
            O => \N__40121\,
            I => \N__40094\
        );

    \I__8806\ : CascadeMux
    port map (
            O => \N__40120\,
            I => \N__40091\
        );

    \I__8805\ : InMux
    port map (
            O => \N__40117\,
            I => \N__40087\
        );

    \I__8804\ : InMux
    port map (
            O => \N__40116\,
            I => \N__40070\
        );

    \I__8803\ : InMux
    port map (
            O => \N__40115\,
            I => \N__40070\
        );

    \I__8802\ : InMux
    port map (
            O => \N__40114\,
            I => \N__40070\
        );

    \I__8801\ : InMux
    port map (
            O => \N__40113\,
            I => \N__40070\
        );

    \I__8800\ : InMux
    port map (
            O => \N__40110\,
            I => \N__40070\
        );

    \I__8799\ : InMux
    port map (
            O => \N__40107\,
            I => \N__40070\
        );

    \I__8798\ : InMux
    port map (
            O => \N__40104\,
            I => \N__40070\
        );

    \I__8797\ : InMux
    port map (
            O => \N__40101\,
            I => \N__40070\
        );

    \I__8796\ : CascadeMux
    port map (
            O => \N__40100\,
            I => \N__40067\
        );

    \I__8795\ : InMux
    port map (
            O => \N__40097\,
            I => \N__40051\
        );

    \I__8794\ : InMux
    port map (
            O => \N__40094\,
            I => \N__40051\
        );

    \I__8793\ : InMux
    port map (
            O => \N__40091\,
            I => \N__40051\
        );

    \I__8792\ : InMux
    port map (
            O => \N__40090\,
            I => \N__40051\
        );

    \I__8791\ : LocalMux
    port map (
            O => \N__40087\,
            I => \N__40048\
        );

    \I__8790\ : LocalMux
    port map (
            O => \N__40070\,
            I => \N__40045\
        );

    \I__8789\ : InMux
    port map (
            O => \N__40067\,
            I => \N__40040\
        );

    \I__8788\ : InMux
    port map (
            O => \N__40066\,
            I => \N__40040\
        );

    \I__8787\ : InMux
    port map (
            O => \N__40065\,
            I => \N__40029\
        );

    \I__8786\ : InMux
    port map (
            O => \N__40064\,
            I => \N__40029\
        );

    \I__8785\ : InMux
    port map (
            O => \N__40063\,
            I => \N__40029\
        );

    \I__8784\ : InMux
    port map (
            O => \N__40062\,
            I => \N__40029\
        );

    \I__8783\ : InMux
    port map (
            O => \N__40061\,
            I => \N__40029\
        );

    \I__8782\ : InMux
    port map (
            O => \N__40060\,
            I => \N__40026\
        );

    \I__8781\ : LocalMux
    port map (
            O => \N__40051\,
            I => \N__40021\
        );

    \I__8780\ : Span4Mux_v
    port map (
            O => \N__40048\,
            I => \N__40018\
        );

    \I__8779\ : Span4Mux_h
    port map (
            O => \N__40045\,
            I => \N__40013\
        );

    \I__8778\ : LocalMux
    port map (
            O => \N__40040\,
            I => \N__40013\
        );

    \I__8777\ : LocalMux
    port map (
            O => \N__40029\,
            I => \N__40010\
        );

    \I__8776\ : LocalMux
    port map (
            O => \N__40026\,
            I => \N__40007\
        );

    \I__8775\ : InMux
    port map (
            O => \N__40025\,
            I => \N__40001\
        );

    \I__8774\ : InMux
    port map (
            O => \N__40024\,
            I => \N__40001\
        );

    \I__8773\ : Span4Mux_v
    port map (
            O => \N__40021\,
            I => \N__39996\
        );

    \I__8772\ : Span4Mux_h
    port map (
            O => \N__40018\,
            I => \N__39996\
        );

    \I__8771\ : Span4Mux_v
    port map (
            O => \N__40013\,
            I => \N__39991\
        );

    \I__8770\ : Span4Mux_h
    port map (
            O => \N__40010\,
            I => \N__39991\
        );

    \I__8769\ : Span4Mux_h
    port map (
            O => \N__40007\,
            I => \N__39988\
        );

    \I__8768\ : InMux
    port map (
            O => \N__40006\,
            I => \N__39985\
        );

    \I__8767\ : LocalMux
    port map (
            O => \N__40001\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__8766\ : Odrv4
    port map (
            O => \N__39996\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__8765\ : Odrv4
    port map (
            O => \N__39991\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__8764\ : Odrv4
    port map (
            O => \N__39988\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__8763\ : LocalMux
    port map (
            O => \N__39985\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__8762\ : CascadeMux
    port map (
            O => \N__39974\,
            I => \N__39971\
        );

    \I__8761\ : InMux
    port map (
            O => \N__39971\,
            I => \N__39968\
        );

    \I__8760\ : LocalMux
    port map (
            O => \N__39968\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19\
        );

    \I__8759\ : InMux
    port map (
            O => \N__39965\,
            I => \N__39939\
        );

    \I__8758\ : InMux
    port map (
            O => \N__39964\,
            I => \N__39939\
        );

    \I__8757\ : InMux
    port map (
            O => \N__39963\,
            I => \N__39939\
        );

    \I__8756\ : InMux
    port map (
            O => \N__39962\,
            I => \N__39939\
        );

    \I__8755\ : CascadeMux
    port map (
            O => \N__39961\,
            I => \N__39933\
        );

    \I__8754\ : CascadeMux
    port map (
            O => \N__39960\,
            I => \N__39930\
        );

    \I__8753\ : CascadeMux
    port map (
            O => \N__39959\,
            I => \N__39927\
        );

    \I__8752\ : InMux
    port map (
            O => \N__39958\,
            I => \N__39924\
        );

    \I__8751\ : InMux
    port map (
            O => \N__39957\,
            I => \N__39920\
        );

    \I__8750\ : InMux
    port map (
            O => \N__39956\,
            I => \N__39917\
        );

    \I__8749\ : InMux
    port map (
            O => \N__39955\,
            I => \N__39898\
        );

    \I__8748\ : InMux
    port map (
            O => \N__39954\,
            I => \N__39898\
        );

    \I__8747\ : InMux
    port map (
            O => \N__39953\,
            I => \N__39898\
        );

    \I__8746\ : InMux
    port map (
            O => \N__39952\,
            I => \N__39898\
        );

    \I__8745\ : InMux
    port map (
            O => \N__39951\,
            I => \N__39898\
        );

    \I__8744\ : InMux
    port map (
            O => \N__39950\,
            I => \N__39898\
        );

    \I__8743\ : InMux
    port map (
            O => \N__39949\,
            I => \N__39898\
        );

    \I__8742\ : InMux
    port map (
            O => \N__39948\,
            I => \N__39898\
        );

    \I__8741\ : LocalMux
    port map (
            O => \N__39939\,
            I => \N__39895\
        );

    \I__8740\ : InMux
    port map (
            O => \N__39938\,
            I => \N__39892\
        );

    \I__8739\ : InMux
    port map (
            O => \N__39937\,
            I => \N__39881\
        );

    \I__8738\ : InMux
    port map (
            O => \N__39936\,
            I => \N__39881\
        );

    \I__8737\ : InMux
    port map (
            O => \N__39933\,
            I => \N__39881\
        );

    \I__8736\ : InMux
    port map (
            O => \N__39930\,
            I => \N__39881\
        );

    \I__8735\ : InMux
    port map (
            O => \N__39927\,
            I => \N__39881\
        );

    \I__8734\ : LocalMux
    port map (
            O => \N__39924\,
            I => \N__39878\
        );

    \I__8733\ : InMux
    port map (
            O => \N__39923\,
            I => \N__39875\
        );

    \I__8732\ : LocalMux
    port map (
            O => \N__39920\,
            I => \N__39870\
        );

    \I__8731\ : LocalMux
    port map (
            O => \N__39917\,
            I => \N__39870\
        );

    \I__8730\ : InMux
    port map (
            O => \N__39916\,
            I => \N__39865\
        );

    \I__8729\ : InMux
    port map (
            O => \N__39915\,
            I => \N__39865\
        );

    \I__8728\ : LocalMux
    port map (
            O => \N__39898\,
            I => \N__39862\
        );

    \I__8727\ : Span4Mux_h
    port map (
            O => \N__39895\,
            I => \N__39859\
        );

    \I__8726\ : LocalMux
    port map (
            O => \N__39892\,
            I => \N__39856\
        );

    \I__8725\ : LocalMux
    port map (
            O => \N__39881\,
            I => \N__39847\
        );

    \I__8724\ : Span4Mux_v
    port map (
            O => \N__39878\,
            I => \N__39847\
        );

    \I__8723\ : LocalMux
    port map (
            O => \N__39875\,
            I => \N__39847\
        );

    \I__8722\ : Span4Mux_h
    port map (
            O => \N__39870\,
            I => \N__39847\
        );

    \I__8721\ : LocalMux
    port map (
            O => \N__39865\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__8720\ : Odrv4
    port map (
            O => \N__39862\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__8719\ : Odrv4
    port map (
            O => \N__39859\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__8718\ : Odrv12
    port map (
            O => \N__39856\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__8717\ : Odrv4
    port map (
            O => \N__39847\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__8716\ : InMux
    port map (
            O => \N__39836\,
            I => \N__39833\
        );

    \I__8715\ : LocalMux
    port map (
            O => \N__39833\,
            I => \N__39829\
        );

    \I__8714\ : InMux
    port map (
            O => \N__39832\,
            I => \N__39826\
        );

    \I__8713\ : Span4Mux_h
    port map (
            O => \N__39829\,
            I => \N__39823\
        );

    \I__8712\ : LocalMux
    port map (
            O => \N__39826\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__8711\ : Odrv4
    port map (
            O => \N__39823\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__8710\ : CEMux
    port map (
            O => \N__39818\,
            I => \N__39814\
        );

    \I__8709\ : CEMux
    port map (
            O => \N__39817\,
            I => \N__39811\
        );

    \I__8708\ : LocalMux
    port map (
            O => \N__39814\,
            I => \N__39808\
        );

    \I__8707\ : LocalMux
    port map (
            O => \N__39811\,
            I => \N__39805\
        );

    \I__8706\ : Span4Mux_v
    port map (
            O => \N__39808\,
            I => \N__39802\
        );

    \I__8705\ : Span4Mux_h
    port map (
            O => \N__39805\,
            I => \N__39798\
        );

    \I__8704\ : Span4Mux_h
    port map (
            O => \N__39802\,
            I => \N__39795\
        );

    \I__8703\ : CEMux
    port map (
            O => \N__39801\,
            I => \N__39792\
        );

    \I__8702\ : Span4Mux_h
    port map (
            O => \N__39798\,
            I => \N__39789\
        );

    \I__8701\ : Sp12to4
    port map (
            O => \N__39795\,
            I => \N__39784\
        );

    \I__8700\ : LocalMux
    port map (
            O => \N__39792\,
            I => \N__39784\
        );

    \I__8699\ : Odrv4
    port map (
            O => \N__39789\,
            I => \phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__8698\ : Odrv12
    port map (
            O => \N__39784\,
            I => \phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__8697\ : InMux
    port map (
            O => \N__39779\,
            I => \N__39776\
        );

    \I__8696\ : LocalMux
    port map (
            O => \N__39776\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_0\
        );

    \I__8695\ : CascadeMux
    port map (
            O => \N__39773\,
            I => \delay_measurement_inst.delay_hc_reg3lto30_2_cascade_\
        );

    \I__8694\ : CascadeMux
    port map (
            O => \N__39770\,
            I => \delay_measurement_inst.delay_hc_reg3_cascade_\
        );

    \I__8693\ : InMux
    port map (
            O => \N__39767\,
            I => \N__39763\
        );

    \I__8692\ : InMux
    port map (
            O => \N__39766\,
            I => \N__39760\
        );

    \I__8691\ : LocalMux
    port map (
            O => \N__39763\,
            I => \N__39755\
        );

    \I__8690\ : LocalMux
    port map (
            O => \N__39760\,
            I => \N__39752\
        );

    \I__8689\ : InMux
    port map (
            O => \N__39759\,
            I => \N__39749\
        );

    \I__8688\ : InMux
    port map (
            O => \N__39758\,
            I => \N__39746\
        );

    \I__8687\ : Span12Mux_v
    port map (
            O => \N__39755\,
            I => \N__39743\
        );

    \I__8686\ : Span4Mux_h
    port map (
            O => \N__39752\,
            I => \N__39740\
        );

    \I__8685\ : LocalMux
    port map (
            O => \N__39749\,
            I => \N__39737\
        );

    \I__8684\ : LocalMux
    port map (
            O => \N__39746\,
            I => measured_delay_hc_4
        );

    \I__8683\ : Odrv12
    port map (
            O => \N__39743\,
            I => measured_delay_hc_4
        );

    \I__8682\ : Odrv4
    port map (
            O => \N__39740\,
            I => measured_delay_hc_4
        );

    \I__8681\ : Odrv4
    port map (
            O => \N__39737\,
            I => measured_delay_hc_4
        );

    \I__8680\ : CascadeMux
    port map (
            O => \N__39728\,
            I => \N__39725\
        );

    \I__8679\ : InMux
    port map (
            O => \N__39725\,
            I => \N__39719\
        );

    \I__8678\ : InMux
    port map (
            O => \N__39724\,
            I => \N__39716\
        );

    \I__8677\ : CascadeMux
    port map (
            O => \N__39723\,
            I => \N__39713\
        );

    \I__8676\ : InMux
    port map (
            O => \N__39722\,
            I => \N__39709\
        );

    \I__8675\ : LocalMux
    port map (
            O => \N__39719\,
            I => \N__39704\
        );

    \I__8674\ : LocalMux
    port map (
            O => \N__39716\,
            I => \N__39704\
        );

    \I__8673\ : InMux
    port map (
            O => \N__39713\,
            I => \N__39701\
        );

    \I__8672\ : CascadeMux
    port map (
            O => \N__39712\,
            I => \N__39698\
        );

    \I__8671\ : LocalMux
    port map (
            O => \N__39709\,
            I => \N__39695\
        );

    \I__8670\ : Span4Mux_v
    port map (
            O => \N__39704\,
            I => \N__39690\
        );

    \I__8669\ : LocalMux
    port map (
            O => \N__39701\,
            I => \N__39690\
        );

    \I__8668\ : InMux
    port map (
            O => \N__39698\,
            I => \N__39687\
        );

    \I__8667\ : Span4Mux_h
    port map (
            O => \N__39695\,
            I => \N__39682\
        );

    \I__8666\ : Span4Mux_h
    port map (
            O => \N__39690\,
            I => \N__39682\
        );

    \I__8665\ : LocalMux
    port map (
            O => \N__39687\,
            I => measured_delay_hc_14
        );

    \I__8664\ : Odrv4
    port map (
            O => \N__39682\,
            I => measured_delay_hc_14
        );

    \I__8663\ : InMux
    port map (
            O => \N__39677\,
            I => \N__39674\
        );

    \I__8662\ : LocalMux
    port map (
            O => \N__39674\,
            I => \N__39670\
        );

    \I__8661\ : InMux
    port map (
            O => \N__39673\,
            I => \N__39667\
        );

    \I__8660\ : Span4Mux_v
    port map (
            O => \N__39670\,
            I => \N__39664\
        );

    \I__8659\ : LocalMux
    port map (
            O => \N__39667\,
            I => measured_delay_hc_24
        );

    \I__8658\ : Odrv4
    port map (
            O => \N__39664\,
            I => measured_delay_hc_24
        );

    \I__8657\ : InMux
    port map (
            O => \N__39659\,
            I => \N__39656\
        );

    \I__8656\ : LocalMux
    port map (
            O => \N__39656\,
            I => \N__39652\
        );

    \I__8655\ : InMux
    port map (
            O => \N__39655\,
            I => \N__39649\
        );

    \I__8654\ : Span4Mux_h
    port map (
            O => \N__39652\,
            I => \N__39646\
        );

    \I__8653\ : LocalMux
    port map (
            O => \N__39649\,
            I => measured_delay_hc_25
        );

    \I__8652\ : Odrv4
    port map (
            O => \N__39646\,
            I => measured_delay_hc_25
        );

    \I__8651\ : CascadeMux
    port map (
            O => \N__39641\,
            I => \N__39638\
        );

    \I__8650\ : InMux
    port map (
            O => \N__39638\,
            I => \N__39635\
        );

    \I__8649\ : LocalMux
    port map (
            O => \N__39635\,
            I => \N__39631\
        );

    \I__8648\ : InMux
    port map (
            O => \N__39634\,
            I => \N__39628\
        );

    \I__8647\ : Span4Mux_h
    port map (
            O => \N__39631\,
            I => \N__39625\
        );

    \I__8646\ : LocalMux
    port map (
            O => \N__39628\,
            I => measured_delay_hc_26
        );

    \I__8645\ : Odrv4
    port map (
            O => \N__39625\,
            I => measured_delay_hc_26
        );

    \I__8644\ : InMux
    port map (
            O => \N__39620\,
            I => \N__39616\
        );

    \I__8643\ : InMux
    port map (
            O => \N__39619\,
            I => \N__39613\
        );

    \I__8642\ : LocalMux
    port map (
            O => \N__39616\,
            I => measured_delay_hc_28
        );

    \I__8641\ : LocalMux
    port map (
            O => \N__39613\,
            I => measured_delay_hc_28
        );

    \I__8640\ : InMux
    port map (
            O => \N__39608\,
            I => \N__39604\
        );

    \I__8639\ : InMux
    port map (
            O => \N__39607\,
            I => \N__39601\
        );

    \I__8638\ : LocalMux
    port map (
            O => \N__39604\,
            I => measured_delay_hc_30
        );

    \I__8637\ : LocalMux
    port map (
            O => \N__39601\,
            I => measured_delay_hc_30
        );

    \I__8636\ : InMux
    port map (
            O => \N__39596\,
            I => \N__39593\
        );

    \I__8635\ : LocalMux
    port map (
            O => \N__39593\,
            I => \N__39588\
        );

    \I__8634\ : InMux
    port map (
            O => \N__39592\,
            I => \N__39585\
        );

    \I__8633\ : InMux
    port map (
            O => \N__39591\,
            I => \N__39582\
        );

    \I__8632\ : Span12Mux_v
    port map (
            O => \N__39588\,
            I => \N__39578\
        );

    \I__8631\ : LocalMux
    port map (
            O => \N__39585\,
            I => \N__39575\
        );

    \I__8630\ : LocalMux
    port map (
            O => \N__39582\,
            I => \N__39572\
        );

    \I__8629\ : InMux
    port map (
            O => \N__39581\,
            I => \N__39569\
        );

    \I__8628\ : Span12Mux_h
    port map (
            O => \N__39578\,
            I => \N__39566\
        );

    \I__8627\ : Span4Mux_h
    port map (
            O => \N__39575\,
            I => \N__39563\
        );

    \I__8626\ : Span4Mux_h
    port map (
            O => \N__39572\,
            I => \N__39560\
        );

    \I__8625\ : LocalMux
    port map (
            O => \N__39569\,
            I => measured_delay_hc_0
        );

    \I__8624\ : Odrv12
    port map (
            O => \N__39566\,
            I => measured_delay_hc_0
        );

    \I__8623\ : Odrv4
    port map (
            O => \N__39563\,
            I => measured_delay_hc_0
        );

    \I__8622\ : Odrv4
    port map (
            O => \N__39560\,
            I => measured_delay_hc_0
        );

    \I__8621\ : InMux
    port map (
            O => \N__39551\,
            I => \N__39527\
        );

    \I__8620\ : InMux
    port map (
            O => \N__39550\,
            I => \N__39527\
        );

    \I__8619\ : InMux
    port map (
            O => \N__39549\,
            I => \N__39527\
        );

    \I__8618\ : InMux
    port map (
            O => \N__39548\,
            I => \N__39527\
        );

    \I__8617\ : InMux
    port map (
            O => \N__39547\,
            I => \N__39518\
        );

    \I__8616\ : InMux
    port map (
            O => \N__39546\,
            I => \N__39518\
        );

    \I__8615\ : InMux
    port map (
            O => \N__39545\,
            I => \N__39518\
        );

    \I__8614\ : InMux
    port map (
            O => \N__39544\,
            I => \N__39518\
        );

    \I__8613\ : InMux
    port map (
            O => \N__39543\,
            I => \N__39495\
        );

    \I__8612\ : InMux
    port map (
            O => \N__39542\,
            I => \N__39495\
        );

    \I__8611\ : InMux
    port map (
            O => \N__39541\,
            I => \N__39495\
        );

    \I__8610\ : InMux
    port map (
            O => \N__39540\,
            I => \N__39495\
        );

    \I__8609\ : InMux
    port map (
            O => \N__39539\,
            I => \N__39486\
        );

    \I__8608\ : InMux
    port map (
            O => \N__39538\,
            I => \N__39486\
        );

    \I__8607\ : InMux
    port map (
            O => \N__39537\,
            I => \N__39486\
        );

    \I__8606\ : InMux
    port map (
            O => \N__39536\,
            I => \N__39486\
        );

    \I__8605\ : LocalMux
    port map (
            O => \N__39527\,
            I => \N__39481\
        );

    \I__8604\ : LocalMux
    port map (
            O => \N__39518\,
            I => \N__39481\
        );

    \I__8603\ : InMux
    port map (
            O => \N__39517\,
            I => \N__39472\
        );

    \I__8602\ : InMux
    port map (
            O => \N__39516\,
            I => \N__39472\
        );

    \I__8601\ : InMux
    port map (
            O => \N__39515\,
            I => \N__39472\
        );

    \I__8600\ : InMux
    port map (
            O => \N__39514\,
            I => \N__39472\
        );

    \I__8599\ : InMux
    port map (
            O => \N__39513\,
            I => \N__39467\
        );

    \I__8598\ : InMux
    port map (
            O => \N__39512\,
            I => \N__39467\
        );

    \I__8597\ : InMux
    port map (
            O => \N__39511\,
            I => \N__39458\
        );

    \I__8596\ : InMux
    port map (
            O => \N__39510\,
            I => \N__39458\
        );

    \I__8595\ : InMux
    port map (
            O => \N__39509\,
            I => \N__39458\
        );

    \I__8594\ : InMux
    port map (
            O => \N__39508\,
            I => \N__39458\
        );

    \I__8593\ : InMux
    port map (
            O => \N__39507\,
            I => \N__39449\
        );

    \I__8592\ : InMux
    port map (
            O => \N__39506\,
            I => \N__39449\
        );

    \I__8591\ : InMux
    port map (
            O => \N__39505\,
            I => \N__39449\
        );

    \I__8590\ : InMux
    port map (
            O => \N__39504\,
            I => \N__39449\
        );

    \I__8589\ : LocalMux
    port map (
            O => \N__39495\,
            I => \N__39444\
        );

    \I__8588\ : LocalMux
    port map (
            O => \N__39486\,
            I => \N__39444\
        );

    \I__8587\ : Sp12to4
    port map (
            O => \N__39481\,
            I => \N__39435\
        );

    \I__8586\ : LocalMux
    port map (
            O => \N__39472\,
            I => \N__39435\
        );

    \I__8585\ : LocalMux
    port map (
            O => \N__39467\,
            I => \N__39435\
        );

    \I__8584\ : LocalMux
    port map (
            O => \N__39458\,
            I => \N__39435\
        );

    \I__8583\ : LocalMux
    port map (
            O => \N__39449\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__8582\ : Odrv4
    port map (
            O => \N__39444\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__8581\ : Odrv12
    port map (
            O => \N__39435\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__8580\ : InMux
    port map (
            O => \N__39428\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_28\
        );

    \I__8579\ : CEMux
    port map (
            O => \N__39425\,
            I => \N__39420\
        );

    \I__8578\ : CEMux
    port map (
            O => \N__39424\,
            I => \N__39417\
        );

    \I__8577\ : CEMux
    port map (
            O => \N__39423\,
            I => \N__39414\
        );

    \I__8576\ : LocalMux
    port map (
            O => \N__39420\,
            I => \N__39411\
        );

    \I__8575\ : LocalMux
    port map (
            O => \N__39417\,
            I => \N__39406\
        );

    \I__8574\ : LocalMux
    port map (
            O => \N__39414\,
            I => \N__39406\
        );

    \I__8573\ : Span4Mux_v
    port map (
            O => \N__39411\,
            I => \N__39402\
        );

    \I__8572\ : Span4Mux_v
    port map (
            O => \N__39406\,
            I => \N__39399\
        );

    \I__8571\ : CEMux
    port map (
            O => \N__39405\,
            I => \N__39396\
        );

    \I__8570\ : Odrv4
    port map (
            O => \N__39402\,
            I => \delay_measurement_inst.delay_hc_timer.N_336_i\
        );

    \I__8569\ : Odrv4
    port map (
            O => \N__39399\,
            I => \delay_measurement_inst.delay_hc_timer.N_336_i\
        );

    \I__8568\ : LocalMux
    port map (
            O => \N__39396\,
            I => \delay_measurement_inst.delay_hc_timer.N_336_i\
        );

    \I__8567\ : CascadeMux
    port map (
            O => \N__39389\,
            I => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_3_cascade_\
        );

    \I__8566\ : CascadeMux
    port map (
            O => \N__39386\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_a1_2_0_cascade_\
        );

    \I__8565\ : CascadeMux
    port map (
            O => \N__39383\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_a1_2_cascade_\
        );

    \I__8564\ : CascadeMux
    port map (
            O => \N__39380\,
            I => \N__39377\
        );

    \I__8563\ : InMux
    port map (
            O => \N__39377\,
            I => \N__39374\
        );

    \I__8562\ : LocalMux
    port map (
            O => \N__39374\,
            I => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1\
        );

    \I__8561\ : InMux
    port map (
            O => \N__39371\,
            I => \N__39368\
        );

    \I__8560\ : LocalMux
    port map (
            O => \N__39368\,
            I => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_4\
        );

    \I__8559\ : InMux
    port map (
            O => \N__39365\,
            I => \N__39361\
        );

    \I__8558\ : InMux
    port map (
            O => \N__39364\,
            I => \N__39358\
        );

    \I__8557\ : LocalMux
    port map (
            O => \N__39361\,
            I => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2\
        );

    \I__8556\ : LocalMux
    port map (
            O => \N__39358\,
            I => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2\
        );

    \I__8555\ : CascadeMux
    port map (
            O => \N__39353\,
            I => \N__39349\
        );

    \I__8554\ : InMux
    port map (
            O => \N__39352\,
            I => \N__39346\
        );

    \I__8553\ : InMux
    port map (
            O => \N__39349\,
            I => \N__39343\
        );

    \I__8552\ : LocalMux
    port map (
            O => \N__39346\,
            I => \N__39340\
        );

    \I__8551\ : LocalMux
    port map (
            O => \N__39343\,
            I => \N__39337\
        );

    \I__8550\ : Span4Mux_v
    port map (
            O => \N__39340\,
            I => \N__39332\
        );

    \I__8549\ : Span4Mux_h
    port map (
            O => \N__39337\,
            I => \N__39332\
        );

    \I__8548\ : Span4Mux_h
    port map (
            O => \N__39332\,
            I => \N__39329\
        );

    \I__8547\ : Span4Mux_h
    port map (
            O => \N__39329\,
            I => \N__39326\
        );

    \I__8546\ : Odrv4
    port map (
            O => \N__39326\,
            I => \delay_measurement_inst.delay_hc_reg3lto30_2\
        );

    \I__8545\ : InMux
    port map (
            O => \N__39323\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_19\
        );

    \I__8544\ : InMux
    port map (
            O => \N__39320\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_20\
        );

    \I__8543\ : InMux
    port map (
            O => \N__39317\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_21\
        );

    \I__8542\ : InMux
    port map (
            O => \N__39314\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_22\
        );

    \I__8541\ : InMux
    port map (
            O => \N__39311\,
            I => \bfn_16_10_0_\
        );

    \I__8540\ : InMux
    port map (
            O => \N__39308\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_24\
        );

    \I__8539\ : InMux
    port map (
            O => \N__39305\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_25\
        );

    \I__8538\ : InMux
    port map (
            O => \N__39302\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_26\
        );

    \I__8537\ : InMux
    port map (
            O => \N__39299\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_27\
        );

    \I__8536\ : InMux
    port map (
            O => \N__39296\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_10\
        );

    \I__8535\ : InMux
    port map (
            O => \N__39293\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_11\
        );

    \I__8534\ : InMux
    port map (
            O => \N__39290\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_12\
        );

    \I__8533\ : InMux
    port map (
            O => \N__39287\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_13\
        );

    \I__8532\ : InMux
    port map (
            O => \N__39284\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_14\
        );

    \I__8531\ : InMux
    port map (
            O => \N__39281\,
            I => \bfn_16_9_0_\
        );

    \I__8530\ : InMux
    port map (
            O => \N__39278\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_16\
        );

    \I__8529\ : InMux
    port map (
            O => \N__39275\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_17\
        );

    \I__8528\ : InMux
    port map (
            O => \N__39272\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_18\
        );

    \I__8527\ : InMux
    port map (
            O => \N__39269\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_1\
        );

    \I__8526\ : InMux
    port map (
            O => \N__39266\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_2\
        );

    \I__8525\ : InMux
    port map (
            O => \N__39263\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_3\
        );

    \I__8524\ : InMux
    port map (
            O => \N__39260\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_4\
        );

    \I__8523\ : InMux
    port map (
            O => \N__39257\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_5\
        );

    \I__8522\ : InMux
    port map (
            O => \N__39254\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_6\
        );

    \I__8521\ : InMux
    port map (
            O => \N__39251\,
            I => \bfn_16_8_0_\
        );

    \I__8520\ : InMux
    port map (
            O => \N__39248\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_8\
        );

    \I__8519\ : InMux
    port map (
            O => \N__39245\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_9\
        );

    \I__8518\ : InMux
    port map (
            O => \N__39242\,
            I => \N__39238\
        );

    \I__8517\ : InMux
    port map (
            O => \N__39241\,
            I => \N__39235\
        );

    \I__8516\ : LocalMux
    port map (
            O => \N__39238\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__8515\ : LocalMux
    port map (
            O => \N__39235\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__8514\ : InMux
    port map (
            O => \N__39230\,
            I => \N__39227\
        );

    \I__8513\ : LocalMux
    port map (
            O => \N__39227\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_19\
        );

    \I__8512\ : InMux
    port map (
            O => \N__39224\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__8511\ : InMux
    port map (
            O => \N__39221\,
            I => \N__39216\
        );

    \I__8510\ : InMux
    port map (
            O => \N__39220\,
            I => \N__39213\
        );

    \I__8509\ : InMux
    port map (
            O => \N__39219\,
            I => \N__39210\
        );

    \I__8508\ : LocalMux
    port map (
            O => \N__39216\,
            I => \N__39207\
        );

    \I__8507\ : LocalMux
    port map (
            O => \N__39213\,
            I => \N__39202\
        );

    \I__8506\ : LocalMux
    port map (
            O => \N__39210\,
            I => \N__39198\
        );

    \I__8505\ : Sp12to4
    port map (
            O => \N__39207\,
            I => \N__39195\
        );

    \I__8504\ : InMux
    port map (
            O => \N__39206\,
            I => \N__39190\
        );

    \I__8503\ : InMux
    port map (
            O => \N__39205\,
            I => \N__39190\
        );

    \I__8502\ : Span4Mux_h
    port map (
            O => \N__39202\,
            I => \N__39187\
        );

    \I__8501\ : InMux
    port map (
            O => \N__39201\,
            I => \N__39184\
        );

    \I__8500\ : Span12Mux_h
    port map (
            O => \N__39198\,
            I => \N__39179\
        );

    \I__8499\ : Span12Mux_v
    port map (
            O => \N__39195\,
            I => \N__39179\
        );

    \I__8498\ : LocalMux
    port map (
            O => \N__39190\,
            I => \N__39176\
        );

    \I__8497\ : Odrv4
    port map (
            O => \N__39187\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__8496\ : LocalMux
    port map (
            O => \N__39184\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__8495\ : Odrv12
    port map (
            O => \N__39179\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__8494\ : Odrv4
    port map (
            O => \N__39176\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__8493\ : CascadeMux
    port map (
            O => \N__39167\,
            I => \N__39164\
        );

    \I__8492\ : InMux
    port map (
            O => \N__39164\,
            I => \N__39161\
        );

    \I__8491\ : LocalMux
    port map (
            O => \N__39161\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\
        );

    \I__8490\ : CascadeMux
    port map (
            O => \N__39158\,
            I => \N__39155\
        );

    \I__8489\ : InMux
    port map (
            O => \N__39155\,
            I => \N__39152\
        );

    \I__8488\ : LocalMux
    port map (
            O => \N__39152\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\
        );

    \I__8487\ : CascadeMux
    port map (
            O => \N__39149\,
            I => \N__39146\
        );

    \I__8486\ : InMux
    port map (
            O => \N__39146\,
            I => \N__39143\
        );

    \I__8485\ : LocalMux
    port map (
            O => \N__39143\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\
        );

    \I__8484\ : InMux
    port map (
            O => \N__39140\,
            I => \N__39136\
        );

    \I__8483\ : InMux
    port map (
            O => \N__39139\,
            I => \N__39133\
        );

    \I__8482\ : LocalMux
    port map (
            O => \N__39136\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__8481\ : LocalMux
    port map (
            O => \N__39133\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__8480\ : InMux
    port map (
            O => \N__39128\,
            I => \N__39123\
        );

    \I__8479\ : InMux
    port map (
            O => \N__39127\,
            I => \N__39120\
        );

    \I__8478\ : InMux
    port map (
            O => \N__39126\,
            I => \N__39117\
        );

    \I__8477\ : LocalMux
    port map (
            O => \N__39123\,
            I => \N__39114\
        );

    \I__8476\ : LocalMux
    port map (
            O => \N__39120\,
            I => \N__39111\
        );

    \I__8475\ : LocalMux
    port map (
            O => \N__39117\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__8474\ : Odrv4
    port map (
            O => \N__39114\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__8473\ : Odrv4
    port map (
            O => \N__39111\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__8472\ : InMux
    port map (
            O => \N__39104\,
            I => \N__39098\
        );

    \I__8471\ : InMux
    port map (
            O => \N__39103\,
            I => \N__39095\
        );

    \I__8470\ : InMux
    port map (
            O => \N__39102\,
            I => \N__39090\
        );

    \I__8469\ : InMux
    port map (
            O => \N__39101\,
            I => \N__39090\
        );

    \I__8468\ : LocalMux
    port map (
            O => \N__39098\,
            I => \N__39087\
        );

    \I__8467\ : LocalMux
    port map (
            O => \N__39095\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__8466\ : LocalMux
    port map (
            O => \N__39090\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__8465\ : Odrv4
    port map (
            O => \N__39087\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__8464\ : InMux
    port map (
            O => \N__39080\,
            I => \bfn_16_7_0_\
        );

    \I__8463\ : InMux
    port map (
            O => \N__39077\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_0\
        );

    \I__8462\ : InMux
    port map (
            O => \N__39074\,
            I => \N__39070\
        );

    \I__8461\ : InMux
    port map (
            O => \N__39073\,
            I => \N__39067\
        );

    \I__8460\ : LocalMux
    port map (
            O => \N__39070\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__8459\ : LocalMux
    port map (
            O => \N__39067\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__8458\ : InMux
    port map (
            O => \N__39062\,
            I => \N__39059\
        );

    \I__8457\ : LocalMux
    port map (
            O => \N__39059\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\
        );

    \I__8456\ : InMux
    port map (
            O => \N__39056\,
            I => \N__39052\
        );

    \I__8455\ : InMux
    port map (
            O => \N__39055\,
            I => \N__39049\
        );

    \I__8454\ : LocalMux
    port map (
            O => \N__39052\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__8453\ : LocalMux
    port map (
            O => \N__39049\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__8452\ : InMux
    port map (
            O => \N__39044\,
            I => \N__39041\
        );

    \I__8451\ : LocalMux
    port map (
            O => \N__39041\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\
        );

    \I__8450\ : InMux
    port map (
            O => \N__39038\,
            I => \N__39034\
        );

    \I__8449\ : InMux
    port map (
            O => \N__39037\,
            I => \N__39031\
        );

    \I__8448\ : LocalMux
    port map (
            O => \N__39034\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__8447\ : LocalMux
    port map (
            O => \N__39031\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__8446\ : InMux
    port map (
            O => \N__39026\,
            I => \N__39023\
        );

    \I__8445\ : LocalMux
    port map (
            O => \N__39023\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\
        );

    \I__8444\ : InMux
    port map (
            O => \N__39020\,
            I => \N__39016\
        );

    \I__8443\ : InMux
    port map (
            O => \N__39019\,
            I => \N__39013\
        );

    \I__8442\ : LocalMux
    port map (
            O => \N__39016\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__8441\ : LocalMux
    port map (
            O => \N__39013\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__8440\ : InMux
    port map (
            O => \N__39008\,
            I => \N__39005\
        );

    \I__8439\ : LocalMux
    port map (
            O => \N__39005\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\
        );

    \I__8438\ : InMux
    port map (
            O => \N__39002\,
            I => \N__38998\
        );

    \I__8437\ : InMux
    port map (
            O => \N__39001\,
            I => \N__38995\
        );

    \I__8436\ : LocalMux
    port map (
            O => \N__38998\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__8435\ : LocalMux
    port map (
            O => \N__38995\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__8434\ : CascadeMux
    port map (
            O => \N__38990\,
            I => \N__38987\
        );

    \I__8433\ : InMux
    port map (
            O => \N__38987\,
            I => \N__38984\
        );

    \I__8432\ : LocalMux
    port map (
            O => \N__38984\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\
        );

    \I__8431\ : CascadeMux
    port map (
            O => \N__38981\,
            I => \N__38978\
        );

    \I__8430\ : InMux
    port map (
            O => \N__38978\,
            I => \N__38975\
        );

    \I__8429\ : LocalMux
    port map (
            O => \N__38975\,
            I => \N__38972\
        );

    \I__8428\ : Odrv4
    port map (
            O => \N__38972\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\
        );

    \I__8427\ : InMux
    port map (
            O => \N__38969\,
            I => \N__38965\
        );

    \I__8426\ : InMux
    port map (
            O => \N__38968\,
            I => \N__38962\
        );

    \I__8425\ : LocalMux
    port map (
            O => \N__38965\,
            I => \N__38959\
        );

    \I__8424\ : LocalMux
    port map (
            O => \N__38962\,
            I => \N__38954\
        );

    \I__8423\ : Span4Mux_h
    port map (
            O => \N__38959\,
            I => \N__38954\
        );

    \I__8422\ : Odrv4
    port map (
            O => \N__38954\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__8421\ : InMux
    port map (
            O => \N__38951\,
            I => \N__38948\
        );

    \I__8420\ : LocalMux
    port map (
            O => \N__38948\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_16\
        );

    \I__8419\ : InMux
    port map (
            O => \N__38945\,
            I => \N__38941\
        );

    \I__8418\ : InMux
    port map (
            O => \N__38944\,
            I => \N__38938\
        );

    \I__8417\ : LocalMux
    port map (
            O => \N__38941\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__8416\ : LocalMux
    port map (
            O => \N__38938\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__8415\ : InMux
    port map (
            O => \N__38933\,
            I => \N__38930\
        );

    \I__8414\ : LocalMux
    port map (
            O => \N__38930\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_17\
        );

    \I__8413\ : InMux
    port map (
            O => \N__38927\,
            I => \N__38923\
        );

    \I__8412\ : InMux
    port map (
            O => \N__38926\,
            I => \N__38920\
        );

    \I__8411\ : LocalMux
    port map (
            O => \N__38923\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__8410\ : LocalMux
    port map (
            O => \N__38920\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__8409\ : InMux
    port map (
            O => \N__38915\,
            I => \N__38912\
        );

    \I__8408\ : LocalMux
    port map (
            O => \N__38912\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_18\
        );

    \I__8407\ : InMux
    port map (
            O => \N__38909\,
            I => \N__38905\
        );

    \I__8406\ : InMux
    port map (
            O => \N__38908\,
            I => \N__38902\
        );

    \I__8405\ : LocalMux
    port map (
            O => \N__38905\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__8404\ : LocalMux
    port map (
            O => \N__38902\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__8403\ : InMux
    port map (
            O => \N__38897\,
            I => \N__38894\
        );

    \I__8402\ : LocalMux
    port map (
            O => \N__38894\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\
        );

    \I__8401\ : InMux
    port map (
            O => \N__38891\,
            I => \N__38887\
        );

    \I__8400\ : InMux
    port map (
            O => \N__38890\,
            I => \N__38884\
        );

    \I__8399\ : LocalMux
    port map (
            O => \N__38887\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__8398\ : LocalMux
    port map (
            O => \N__38884\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__8397\ : InMux
    port map (
            O => \N__38879\,
            I => \N__38876\
        );

    \I__8396\ : LocalMux
    port map (
            O => \N__38876\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\
        );

    \I__8395\ : InMux
    port map (
            O => \N__38873\,
            I => \N__38869\
        );

    \I__8394\ : InMux
    port map (
            O => \N__38872\,
            I => \N__38866\
        );

    \I__8393\ : LocalMux
    port map (
            O => \N__38869\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__8392\ : LocalMux
    port map (
            O => \N__38866\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__8391\ : CascadeMux
    port map (
            O => \N__38861\,
            I => \N__38858\
        );

    \I__8390\ : InMux
    port map (
            O => \N__38858\,
            I => \N__38855\
        );

    \I__8389\ : LocalMux
    port map (
            O => \N__38855\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\
        );

    \I__8388\ : InMux
    port map (
            O => \N__38852\,
            I => \N__38848\
        );

    \I__8387\ : InMux
    port map (
            O => \N__38851\,
            I => \N__38845\
        );

    \I__8386\ : LocalMux
    port map (
            O => \N__38848\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__8385\ : LocalMux
    port map (
            O => \N__38845\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__8384\ : InMux
    port map (
            O => \N__38840\,
            I => \N__38837\
        );

    \I__8383\ : LocalMux
    port map (
            O => \N__38837\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\
        );

    \I__8382\ : InMux
    port map (
            O => \N__38834\,
            I => \N__38830\
        );

    \I__8381\ : InMux
    port map (
            O => \N__38833\,
            I => \N__38827\
        );

    \I__8380\ : LocalMux
    port map (
            O => \N__38830\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__8379\ : LocalMux
    port map (
            O => \N__38827\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__8378\ : InMux
    port map (
            O => \N__38822\,
            I => \N__38819\
        );

    \I__8377\ : LocalMux
    port map (
            O => \N__38819\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\
        );

    \I__8376\ : CascadeMux
    port map (
            O => \N__38816\,
            I => \N__38813\
        );

    \I__8375\ : InMux
    port map (
            O => \N__38813\,
            I => \N__38809\
        );

    \I__8374\ : InMux
    port map (
            O => \N__38812\,
            I => \N__38806\
        );

    \I__8373\ : LocalMux
    port map (
            O => \N__38809\,
            I => \N__38803\
        );

    \I__8372\ : LocalMux
    port map (
            O => \N__38806\,
            I => \N__38800\
        );

    \I__8371\ : Odrv4
    port map (
            O => \N__38803\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__8370\ : Odrv4
    port map (
            O => \N__38800\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__8369\ : InMux
    port map (
            O => \N__38795\,
            I => \N__38792\
        );

    \I__8368\ : LocalMux
    port map (
            O => \N__38792\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\
        );

    \I__8367\ : InMux
    port map (
            O => \N__38789\,
            I => \N__38785\
        );

    \I__8366\ : InMux
    port map (
            O => \N__38788\,
            I => \N__38782\
        );

    \I__8365\ : LocalMux
    port map (
            O => \N__38785\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__8364\ : LocalMux
    port map (
            O => \N__38782\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__8363\ : InMux
    port map (
            O => \N__38777\,
            I => \N__38774\
        );

    \I__8362\ : LocalMux
    port map (
            O => \N__38774\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\
        );

    \I__8361\ : InMux
    port map (
            O => \N__38771\,
            I => \N__38768\
        );

    \I__8360\ : LocalMux
    port map (
            O => \N__38768\,
            I => \N__38764\
        );

    \I__8359\ : InMux
    port map (
            O => \N__38767\,
            I => \N__38761\
        );

    \I__8358\ : Span4Mux_h
    port map (
            O => \N__38764\,
            I => \N__38758\
        );

    \I__8357\ : LocalMux
    port map (
            O => \N__38761\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__8356\ : Odrv4
    port map (
            O => \N__38758\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__8355\ : InMux
    port map (
            O => \N__38753\,
            I => \N__38750\
        );

    \I__8354\ : LocalMux
    port map (
            O => \N__38750\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_17\
        );

    \I__8353\ : InMux
    port map (
            O => \N__38747\,
            I => \N__38744\
        );

    \I__8352\ : LocalMux
    port map (
            O => \N__38744\,
            I => \N__38740\
        );

    \I__8351\ : InMux
    port map (
            O => \N__38743\,
            I => \N__38737\
        );

    \I__8350\ : Span4Mux_h
    port map (
            O => \N__38740\,
            I => \N__38734\
        );

    \I__8349\ : LocalMux
    port map (
            O => \N__38737\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__8348\ : Odrv4
    port map (
            O => \N__38734\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__8347\ : InMux
    port map (
            O => \N__38729\,
            I => \N__38726\
        );

    \I__8346\ : LocalMux
    port map (
            O => \N__38726\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_18\
        );

    \I__8345\ : InMux
    port map (
            O => \N__38723\,
            I => \N__38719\
        );

    \I__8344\ : InMux
    port map (
            O => \N__38722\,
            I => \N__38716\
        );

    \I__8343\ : LocalMux
    port map (
            O => \N__38719\,
            I => \N__38713\
        );

    \I__8342\ : LocalMux
    port map (
            O => \N__38716\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__8341\ : Odrv4
    port map (
            O => \N__38713\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__8340\ : InMux
    port map (
            O => \N__38708\,
            I => \N__38705\
        );

    \I__8339\ : LocalMux
    port map (
            O => \N__38705\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_19\
        );

    \I__8338\ : InMux
    port map (
            O => \N__38702\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__8337\ : InMux
    port map (
            O => \N__38699\,
            I => \N__38692\
        );

    \I__8336\ : InMux
    port map (
            O => \N__38698\,
            I => \N__38692\
        );

    \I__8335\ : InMux
    port map (
            O => \N__38697\,
            I => \N__38689\
        );

    \I__8334\ : LocalMux
    port map (
            O => \N__38692\,
            I => \N__38686\
        );

    \I__8333\ : LocalMux
    port map (
            O => \N__38689\,
            I => \N__38683\
        );

    \I__8332\ : Span4Mux_v
    port map (
            O => \N__38686\,
            I => \N__38677\
        );

    \I__8331\ : Span4Mux_h
    port map (
            O => \N__38683\,
            I => \N__38674\
        );

    \I__8330\ : InMux
    port map (
            O => \N__38682\,
            I => \N__38671\
        );

    \I__8329\ : InMux
    port map (
            O => \N__38681\,
            I => \N__38668\
        );

    \I__8328\ : InMux
    port map (
            O => \N__38680\,
            I => \N__38665\
        );

    \I__8327\ : Span4Mux_v
    port map (
            O => \N__38677\,
            I => \N__38662\
        );

    \I__8326\ : Span4Mux_v
    port map (
            O => \N__38674\,
            I => \N__38659\
        );

    \I__8325\ : LocalMux
    port map (
            O => \N__38671\,
            I => \N__38656\
        );

    \I__8324\ : LocalMux
    port map (
            O => \N__38668\,
            I => \N__38651\
        );

    \I__8323\ : LocalMux
    port map (
            O => \N__38665\,
            I => \N__38651\
        );

    \I__8322\ : Odrv4
    port map (
            O => \N__38662\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__8321\ : Odrv4
    port map (
            O => \N__38659\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__8320\ : Odrv4
    port map (
            O => \N__38656\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__8319\ : Odrv12
    port map (
            O => \N__38651\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__8318\ : CascadeMux
    port map (
            O => \N__38642\,
            I => \N__38639\
        );

    \I__8317\ : InMux
    port map (
            O => \N__38639\,
            I => \N__38636\
        );

    \I__8316\ : LocalMux
    port map (
            O => \N__38636\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_17\
        );

    \I__8315\ : CascadeMux
    port map (
            O => \N__38633\,
            I => \N__38630\
        );

    \I__8314\ : InMux
    port map (
            O => \N__38630\,
            I => \N__38627\
        );

    \I__8313\ : LocalMux
    port map (
            O => \N__38627\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_18\
        );

    \I__8312\ : InMux
    port map (
            O => \N__38624\,
            I => \N__38621\
        );

    \I__8311\ : LocalMux
    port map (
            O => \N__38621\,
            I => \N__38617\
        );

    \I__8310\ : CascadeMux
    port map (
            O => \N__38620\,
            I => \N__38614\
        );

    \I__8309\ : Span12Mux_v
    port map (
            O => \N__38617\,
            I => \N__38610\
        );

    \I__8308\ : InMux
    port map (
            O => \N__38614\,
            I => \N__38607\
        );

    \I__8307\ : InMux
    port map (
            O => \N__38613\,
            I => \N__38604\
        );

    \I__8306\ : Odrv12
    port map (
            O => \N__38610\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__8305\ : LocalMux
    port map (
            O => \N__38607\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__8304\ : LocalMux
    port map (
            O => \N__38604\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__8303\ : InMux
    port map (
            O => \N__38597\,
            I => \N__38594\
        );

    \I__8302\ : LocalMux
    port map (
            O => \N__38594\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\
        );

    \I__8301\ : InMux
    port map (
            O => \N__38591\,
            I => \N__38587\
        );

    \I__8300\ : InMux
    port map (
            O => \N__38590\,
            I => \N__38584\
        );

    \I__8299\ : LocalMux
    port map (
            O => \N__38587\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__8298\ : LocalMux
    port map (
            O => \N__38584\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__8297\ : CascadeMux
    port map (
            O => \N__38579\,
            I => \N__38576\
        );

    \I__8296\ : InMux
    port map (
            O => \N__38576\,
            I => \N__38573\
        );

    \I__8295\ : LocalMux
    port map (
            O => \N__38573\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\
        );

    \I__8294\ : CascadeMux
    port map (
            O => \N__38570\,
            I => \N__38567\
        );

    \I__8293\ : InMux
    port map (
            O => \N__38567\,
            I => \N__38563\
        );

    \I__8292\ : InMux
    port map (
            O => \N__38566\,
            I => \N__38560\
        );

    \I__8291\ : LocalMux
    port map (
            O => \N__38563\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__8290\ : LocalMux
    port map (
            O => \N__38560\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__8289\ : InMux
    port map (
            O => \N__38555\,
            I => \N__38552\
        );

    \I__8288\ : LocalMux
    port map (
            O => \N__38552\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\
        );

    \I__8287\ : InMux
    port map (
            O => \N__38549\,
            I => \N__38545\
        );

    \I__8286\ : InMux
    port map (
            O => \N__38548\,
            I => \N__38542\
        );

    \I__8285\ : LocalMux
    port map (
            O => \N__38545\,
            I => \N__38539\
        );

    \I__8284\ : LocalMux
    port map (
            O => \N__38542\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__8283\ : Odrv4
    port map (
            O => \N__38539\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__8282\ : InMux
    port map (
            O => \N__38534\,
            I => \N__38531\
        );

    \I__8281\ : LocalMux
    port map (
            O => \N__38531\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_10\
        );

    \I__8280\ : InMux
    port map (
            O => \N__38528\,
            I => \N__38524\
        );

    \I__8279\ : InMux
    port map (
            O => \N__38527\,
            I => \N__38521\
        );

    \I__8278\ : LocalMux
    port map (
            O => \N__38524\,
            I => \N__38518\
        );

    \I__8277\ : LocalMux
    port map (
            O => \N__38521\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__8276\ : Odrv4
    port map (
            O => \N__38518\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__8275\ : InMux
    port map (
            O => \N__38513\,
            I => \N__38510\
        );

    \I__8274\ : LocalMux
    port map (
            O => \N__38510\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_11\
        );

    \I__8273\ : InMux
    port map (
            O => \N__38507\,
            I => \N__38503\
        );

    \I__8272\ : InMux
    port map (
            O => \N__38506\,
            I => \N__38500\
        );

    \I__8271\ : LocalMux
    port map (
            O => \N__38503\,
            I => \N__38497\
        );

    \I__8270\ : LocalMux
    port map (
            O => \N__38500\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__8269\ : Odrv4
    port map (
            O => \N__38497\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__8268\ : InMux
    port map (
            O => \N__38492\,
            I => \N__38489\
        );

    \I__8267\ : LocalMux
    port map (
            O => \N__38489\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_12\
        );

    \I__8266\ : InMux
    port map (
            O => \N__38486\,
            I => \N__38482\
        );

    \I__8265\ : InMux
    port map (
            O => \N__38485\,
            I => \N__38479\
        );

    \I__8264\ : LocalMux
    port map (
            O => \N__38482\,
            I => \N__38476\
        );

    \I__8263\ : LocalMux
    port map (
            O => \N__38479\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__8262\ : Odrv4
    port map (
            O => \N__38476\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__8261\ : InMux
    port map (
            O => \N__38471\,
            I => \N__38468\
        );

    \I__8260\ : LocalMux
    port map (
            O => \N__38468\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_13\
        );

    \I__8259\ : InMux
    port map (
            O => \N__38465\,
            I => \N__38461\
        );

    \I__8258\ : InMux
    port map (
            O => \N__38464\,
            I => \N__38458\
        );

    \I__8257\ : LocalMux
    port map (
            O => \N__38461\,
            I => \N__38455\
        );

    \I__8256\ : LocalMux
    port map (
            O => \N__38458\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__8255\ : Odrv4
    port map (
            O => \N__38455\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__8254\ : InMux
    port map (
            O => \N__38450\,
            I => \N__38447\
        );

    \I__8253\ : LocalMux
    port map (
            O => \N__38447\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_14\
        );

    \I__8252\ : InMux
    port map (
            O => \N__38444\,
            I => \N__38440\
        );

    \I__8251\ : InMux
    port map (
            O => \N__38443\,
            I => \N__38437\
        );

    \I__8250\ : LocalMux
    port map (
            O => \N__38440\,
            I => \N__38434\
        );

    \I__8249\ : LocalMux
    port map (
            O => \N__38437\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__8248\ : Odrv4
    port map (
            O => \N__38434\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__8247\ : CascadeMux
    port map (
            O => \N__38429\,
            I => \N__38426\
        );

    \I__8246\ : InMux
    port map (
            O => \N__38426\,
            I => \N__38423\
        );

    \I__8245\ : LocalMux
    port map (
            O => \N__38423\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_15\
        );

    \I__8244\ : CascadeMux
    port map (
            O => \N__38420\,
            I => \N__38417\
        );

    \I__8243\ : InMux
    port map (
            O => \N__38417\,
            I => \N__38414\
        );

    \I__8242\ : LocalMux
    port map (
            O => \N__38414\,
            I => \N__38411\
        );

    \I__8241\ : Odrv12
    port map (
            O => \N__38411\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_16\
        );

    \I__8240\ : InMux
    port map (
            O => \N__38408\,
            I => \N__38404\
        );

    \I__8239\ : CascadeMux
    port map (
            O => \N__38407\,
            I => \N__38401\
        );

    \I__8238\ : LocalMux
    port map (
            O => \N__38404\,
            I => \N__38398\
        );

    \I__8237\ : InMux
    port map (
            O => \N__38401\,
            I => \N__38395\
        );

    \I__8236\ : Span4Mux_v
    port map (
            O => \N__38398\,
            I => \N__38392\
        );

    \I__8235\ : LocalMux
    port map (
            O => \N__38395\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__8234\ : Odrv4
    port map (
            O => \N__38392\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__8233\ : InMux
    port map (
            O => \N__38387\,
            I => \N__38384\
        );

    \I__8232\ : LocalMux
    port map (
            O => \N__38384\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_16\
        );

    \I__8231\ : InMux
    port map (
            O => \N__38381\,
            I => \N__38378\
        );

    \I__8230\ : LocalMux
    port map (
            O => \N__38378\,
            I => \N__38374\
        );

    \I__8229\ : InMux
    port map (
            O => \N__38377\,
            I => \N__38371\
        );

    \I__8228\ : Odrv4
    port map (
            O => \N__38374\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__8227\ : LocalMux
    port map (
            O => \N__38371\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__8226\ : InMux
    port map (
            O => \N__38366\,
            I => \N__38363\
        );

    \I__8225\ : LocalMux
    port map (
            O => \N__38363\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_2\
        );

    \I__8224\ : CascadeMux
    port map (
            O => \N__38360\,
            I => \N__38357\
        );

    \I__8223\ : InMux
    port map (
            O => \N__38357\,
            I => \N__38354\
        );

    \I__8222\ : LocalMux
    port map (
            O => \N__38354\,
            I => \N__38350\
        );

    \I__8221\ : InMux
    port map (
            O => \N__38353\,
            I => \N__38347\
        );

    \I__8220\ : Odrv4
    port map (
            O => \N__38350\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__8219\ : LocalMux
    port map (
            O => \N__38347\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__8218\ : InMux
    port map (
            O => \N__38342\,
            I => \N__38339\
        );

    \I__8217\ : LocalMux
    port map (
            O => \N__38339\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_3\
        );

    \I__8216\ : InMux
    port map (
            O => \N__38336\,
            I => \N__38333\
        );

    \I__8215\ : LocalMux
    port map (
            O => \N__38333\,
            I => \N__38329\
        );

    \I__8214\ : InMux
    port map (
            O => \N__38332\,
            I => \N__38326\
        );

    \I__8213\ : Odrv4
    port map (
            O => \N__38329\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__8212\ : LocalMux
    port map (
            O => \N__38326\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__8211\ : InMux
    port map (
            O => \N__38321\,
            I => \N__38318\
        );

    \I__8210\ : LocalMux
    port map (
            O => \N__38318\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_4\
        );

    \I__8209\ : InMux
    port map (
            O => \N__38315\,
            I => \N__38312\
        );

    \I__8208\ : LocalMux
    port map (
            O => \N__38312\,
            I => \N__38308\
        );

    \I__8207\ : InMux
    port map (
            O => \N__38311\,
            I => \N__38305\
        );

    \I__8206\ : Odrv12
    port map (
            O => \N__38308\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__8205\ : LocalMux
    port map (
            O => \N__38305\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__8204\ : InMux
    port map (
            O => \N__38300\,
            I => \N__38297\
        );

    \I__8203\ : LocalMux
    port map (
            O => \N__38297\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_5\
        );

    \I__8202\ : CascadeMux
    port map (
            O => \N__38294\,
            I => \N__38291\
        );

    \I__8201\ : InMux
    port map (
            O => \N__38291\,
            I => \N__38288\
        );

    \I__8200\ : LocalMux
    port map (
            O => \N__38288\,
            I => \N__38284\
        );

    \I__8199\ : InMux
    port map (
            O => \N__38287\,
            I => \N__38281\
        );

    \I__8198\ : Odrv12
    port map (
            O => \N__38284\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__8197\ : LocalMux
    port map (
            O => \N__38281\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__8196\ : InMux
    port map (
            O => \N__38276\,
            I => \N__38273\
        );

    \I__8195\ : LocalMux
    port map (
            O => \N__38273\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_6\
        );

    \I__8194\ : InMux
    port map (
            O => \N__38270\,
            I => \N__38266\
        );

    \I__8193\ : InMux
    port map (
            O => \N__38269\,
            I => \N__38263\
        );

    \I__8192\ : LocalMux
    port map (
            O => \N__38266\,
            I => \N__38260\
        );

    \I__8191\ : LocalMux
    port map (
            O => \N__38263\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__8190\ : Odrv4
    port map (
            O => \N__38260\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__8189\ : InMux
    port map (
            O => \N__38255\,
            I => \N__38252\
        );

    \I__8188\ : LocalMux
    port map (
            O => \N__38252\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_7\
        );

    \I__8187\ : CascadeMux
    port map (
            O => \N__38249\,
            I => \N__38246\
        );

    \I__8186\ : InMux
    port map (
            O => \N__38246\,
            I => \N__38243\
        );

    \I__8185\ : LocalMux
    port map (
            O => \N__38243\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_8\
        );

    \I__8184\ : InMux
    port map (
            O => \N__38240\,
            I => \N__38236\
        );

    \I__8183\ : InMux
    port map (
            O => \N__38239\,
            I => \N__38233\
        );

    \I__8182\ : LocalMux
    port map (
            O => \N__38236\,
            I => \N__38230\
        );

    \I__8181\ : LocalMux
    port map (
            O => \N__38233\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__8180\ : Odrv4
    port map (
            O => \N__38230\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__8179\ : InMux
    port map (
            O => \N__38225\,
            I => \N__38222\
        );

    \I__8178\ : LocalMux
    port map (
            O => \N__38222\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_8\
        );

    \I__8177\ : InMux
    port map (
            O => \N__38219\,
            I => \N__38215\
        );

    \I__8176\ : InMux
    port map (
            O => \N__38218\,
            I => \N__38212\
        );

    \I__8175\ : LocalMux
    port map (
            O => \N__38215\,
            I => \N__38209\
        );

    \I__8174\ : LocalMux
    port map (
            O => \N__38212\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__8173\ : Odrv4
    port map (
            O => \N__38209\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__8172\ : InMux
    port map (
            O => \N__38204\,
            I => \N__38201\
        );

    \I__8171\ : LocalMux
    port map (
            O => \N__38201\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_9\
        );

    \I__8170\ : InMux
    port map (
            O => \N__38198\,
            I => \N__38195\
        );

    \I__8169\ : LocalMux
    port map (
            O => \N__38195\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10\
        );

    \I__8168\ : InMux
    port map (
            O => \N__38192\,
            I => \N__38186\
        );

    \I__8167\ : InMux
    port map (
            O => \N__38191\,
            I => \N__38183\
        );

    \I__8166\ : InMux
    port map (
            O => \N__38190\,
            I => \N__38180\
        );

    \I__8165\ : InMux
    port map (
            O => \N__38189\,
            I => \N__38177\
        );

    \I__8164\ : LocalMux
    port map (
            O => \N__38186\,
            I => \N__38170\
        );

    \I__8163\ : LocalMux
    port map (
            O => \N__38183\,
            I => \N__38170\
        );

    \I__8162\ : LocalMux
    port map (
            O => \N__38180\,
            I => \N__38170\
        );

    \I__8161\ : LocalMux
    port map (
            O => \N__38177\,
            I => \N__38167\
        );

    \I__8160\ : Span4Mux_v
    port map (
            O => \N__38170\,
            I => \N__38164\
        );

    \I__8159\ : Odrv4
    port map (
            O => \N__38167\,
            I => \phase_controller_slave.stoper_tr.time_passed11\
        );

    \I__8158\ : Odrv4
    port map (
            O => \N__38164\,
            I => \phase_controller_slave.stoper_tr.time_passed11\
        );

    \I__8157\ : CascadeMux
    port map (
            O => \N__38159\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\
        );

    \I__8156\ : InMux
    port map (
            O => \N__38156\,
            I => \N__38153\
        );

    \I__8155\ : LocalMux
    port map (
            O => \N__38153\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11\
        );

    \I__8154\ : InMux
    port map (
            O => \N__38150\,
            I => \N__38147\
        );

    \I__8153\ : LocalMux
    port map (
            O => \N__38147\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12\
        );

    \I__8152\ : InMux
    port map (
            O => \N__38144\,
            I => \N__38141\
        );

    \I__8151\ : LocalMux
    port map (
            O => \N__38141\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13\
        );

    \I__8150\ : InMux
    port map (
            O => \N__38138\,
            I => \N__38135\
        );

    \I__8149\ : LocalMux
    port map (
            O => \N__38135\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14\
        );

    \I__8148\ : CascadeMux
    port map (
            O => \N__38132\,
            I => \N__38126\
        );

    \I__8147\ : CascadeMux
    port map (
            O => \N__38131\,
            I => \N__38110\
        );

    \I__8146\ : CascadeMux
    port map (
            O => \N__38130\,
            I => \N__38107\
        );

    \I__8145\ : InMux
    port map (
            O => \N__38129\,
            I => \N__38089\
        );

    \I__8144\ : InMux
    port map (
            O => \N__38126\,
            I => \N__38089\
        );

    \I__8143\ : InMux
    port map (
            O => \N__38125\,
            I => \N__38089\
        );

    \I__8142\ : InMux
    port map (
            O => \N__38124\,
            I => \N__38089\
        );

    \I__8141\ : InMux
    port map (
            O => \N__38123\,
            I => \N__38089\
        );

    \I__8140\ : InMux
    port map (
            O => \N__38122\,
            I => \N__38089\
        );

    \I__8139\ : InMux
    port map (
            O => \N__38121\,
            I => \N__38089\
        );

    \I__8138\ : InMux
    port map (
            O => \N__38120\,
            I => \N__38072\
        );

    \I__8137\ : InMux
    port map (
            O => \N__38119\,
            I => \N__38072\
        );

    \I__8136\ : InMux
    port map (
            O => \N__38118\,
            I => \N__38072\
        );

    \I__8135\ : InMux
    port map (
            O => \N__38117\,
            I => \N__38072\
        );

    \I__8134\ : InMux
    port map (
            O => \N__38116\,
            I => \N__38072\
        );

    \I__8133\ : InMux
    port map (
            O => \N__38115\,
            I => \N__38072\
        );

    \I__8132\ : InMux
    port map (
            O => \N__38114\,
            I => \N__38072\
        );

    \I__8131\ : InMux
    port map (
            O => \N__38113\,
            I => \N__38072\
        );

    \I__8130\ : InMux
    port map (
            O => \N__38110\,
            I => \N__38063\
        );

    \I__8129\ : InMux
    port map (
            O => \N__38107\,
            I => \N__38063\
        );

    \I__8128\ : InMux
    port map (
            O => \N__38106\,
            I => \N__38063\
        );

    \I__8127\ : InMux
    port map (
            O => \N__38105\,
            I => \N__38063\
        );

    \I__8126\ : CascadeMux
    port map (
            O => \N__38104\,
            I => \N__38059\
        );

    \I__8125\ : LocalMux
    port map (
            O => \N__38089\,
            I => \N__38055\
        );

    \I__8124\ : LocalMux
    port map (
            O => \N__38072\,
            I => \N__38052\
        );

    \I__8123\ : LocalMux
    port map (
            O => \N__38063\,
            I => \N__38049\
        );

    \I__8122\ : InMux
    port map (
            O => \N__38062\,
            I => \N__38042\
        );

    \I__8121\ : InMux
    port map (
            O => \N__38059\,
            I => \N__38042\
        );

    \I__8120\ : InMux
    port map (
            O => \N__38058\,
            I => \N__38039\
        );

    \I__8119\ : Span4Mux_v
    port map (
            O => \N__38055\,
            I => \N__38034\
        );

    \I__8118\ : Span4Mux_v
    port map (
            O => \N__38052\,
            I => \N__38034\
        );

    \I__8117\ : Span4Mux_h
    port map (
            O => \N__38049\,
            I => \N__38031\
        );

    \I__8116\ : InMux
    port map (
            O => \N__38048\,
            I => \N__38026\
        );

    \I__8115\ : InMux
    port map (
            O => \N__38047\,
            I => \N__38026\
        );

    \I__8114\ : LocalMux
    port map (
            O => \N__38042\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__8113\ : LocalMux
    port map (
            O => \N__38039\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__8112\ : Odrv4
    port map (
            O => \N__38034\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__8111\ : Odrv4
    port map (
            O => \N__38031\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__8110\ : LocalMux
    port map (
            O => \N__38026\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__8109\ : CascadeMux
    port map (
            O => \N__38015\,
            I => \N__38004\
        );

    \I__8108\ : CascadeMux
    port map (
            O => \N__38014\,
            I => \N__38001\
        );

    \I__8107\ : CascadeMux
    port map (
            O => \N__38013\,
            I => \N__37998\
        );

    \I__8106\ : CascadeMux
    port map (
            O => \N__38012\,
            I => \N__37995\
        );

    \I__8105\ : CascadeMux
    port map (
            O => \N__38011\,
            I => \N__37988\
        );

    \I__8104\ : CascadeMux
    port map (
            O => \N__38010\,
            I => \N__37985\
        );

    \I__8103\ : CascadeMux
    port map (
            O => \N__38009\,
            I => \N__37982\
        );

    \I__8102\ : CascadeMux
    port map (
            O => \N__38008\,
            I => \N__37975\
        );

    \I__8101\ : InMux
    port map (
            O => \N__38007\,
            I => \N__37969\
        );

    \I__8100\ : InMux
    port map (
            O => \N__38004\,
            I => \N__37952\
        );

    \I__8099\ : InMux
    port map (
            O => \N__38001\,
            I => \N__37952\
        );

    \I__8098\ : InMux
    port map (
            O => \N__37998\,
            I => \N__37952\
        );

    \I__8097\ : InMux
    port map (
            O => \N__37995\,
            I => \N__37952\
        );

    \I__8096\ : InMux
    port map (
            O => \N__37994\,
            I => \N__37952\
        );

    \I__8095\ : InMux
    port map (
            O => \N__37993\,
            I => \N__37952\
        );

    \I__8094\ : InMux
    port map (
            O => \N__37992\,
            I => \N__37952\
        );

    \I__8093\ : InMux
    port map (
            O => \N__37991\,
            I => \N__37952\
        );

    \I__8092\ : InMux
    port map (
            O => \N__37988\,
            I => \N__37939\
        );

    \I__8091\ : InMux
    port map (
            O => \N__37985\,
            I => \N__37939\
        );

    \I__8090\ : InMux
    port map (
            O => \N__37982\,
            I => \N__37939\
        );

    \I__8089\ : InMux
    port map (
            O => \N__37981\,
            I => \N__37939\
        );

    \I__8088\ : InMux
    port map (
            O => \N__37980\,
            I => \N__37939\
        );

    \I__8087\ : InMux
    port map (
            O => \N__37979\,
            I => \N__37939\
        );

    \I__8086\ : CascadeMux
    port map (
            O => \N__37978\,
            I => \N__37935\
        );

    \I__8085\ : InMux
    port map (
            O => \N__37975\,
            I => \N__37928\
        );

    \I__8084\ : InMux
    port map (
            O => \N__37974\,
            I => \N__37928\
        );

    \I__8083\ : InMux
    port map (
            O => \N__37973\,
            I => \N__37925\
        );

    \I__8082\ : CascadeMux
    port map (
            O => \N__37972\,
            I => \N__37922\
        );

    \I__8081\ : LocalMux
    port map (
            O => \N__37969\,
            I => \N__37914\
        );

    \I__8080\ : LocalMux
    port map (
            O => \N__37952\,
            I => \N__37914\
        );

    \I__8079\ : LocalMux
    port map (
            O => \N__37939\,
            I => \N__37914\
        );

    \I__8078\ : InMux
    port map (
            O => \N__37938\,
            I => \N__37905\
        );

    \I__8077\ : InMux
    port map (
            O => \N__37935\,
            I => \N__37905\
        );

    \I__8076\ : InMux
    port map (
            O => \N__37934\,
            I => \N__37905\
        );

    \I__8075\ : InMux
    port map (
            O => \N__37933\,
            I => \N__37905\
        );

    \I__8074\ : LocalMux
    port map (
            O => \N__37928\,
            I => \N__37900\
        );

    \I__8073\ : LocalMux
    port map (
            O => \N__37925\,
            I => \N__37900\
        );

    \I__8072\ : InMux
    port map (
            O => \N__37922\,
            I => \N__37897\
        );

    \I__8071\ : InMux
    port map (
            O => \N__37921\,
            I => \N__37894\
        );

    \I__8070\ : Span4Mux_v
    port map (
            O => \N__37914\,
            I => \N__37891\
        );

    \I__8069\ : LocalMux
    port map (
            O => \N__37905\,
            I => \N__37888\
        );

    \I__8068\ : Span4Mux_v
    port map (
            O => \N__37900\,
            I => \N__37885\
        );

    \I__8067\ : LocalMux
    port map (
            O => \N__37897\,
            I => \phase_controller_slave.start_timer_trZ0\
        );

    \I__8066\ : LocalMux
    port map (
            O => \N__37894\,
            I => \phase_controller_slave.start_timer_trZ0\
        );

    \I__8065\ : Odrv4
    port map (
            O => \N__37891\,
            I => \phase_controller_slave.start_timer_trZ0\
        );

    \I__8064\ : Odrv4
    port map (
            O => \N__37888\,
            I => \phase_controller_slave.start_timer_trZ0\
        );

    \I__8063\ : Odrv4
    port map (
            O => \N__37885\,
            I => \phase_controller_slave.start_timer_trZ0\
        );

    \I__8062\ : CascadeMux
    port map (
            O => \N__37874\,
            I => \N__37866\
        );

    \I__8061\ : CascadeMux
    port map (
            O => \N__37873\,
            I => \N__37863\
        );

    \I__8060\ : CascadeMux
    port map (
            O => \N__37872\,
            I => \N__37855\
        );

    \I__8059\ : CascadeMux
    port map (
            O => \N__37871\,
            I => \N__37852\
        );

    \I__8058\ : CascadeMux
    port map (
            O => \N__37870\,
            I => \N__37849\
        );

    \I__8057\ : CascadeMux
    port map (
            O => \N__37869\,
            I => \N__37846\
        );

    \I__8056\ : InMux
    port map (
            O => \N__37866\,
            I => \N__37833\
        );

    \I__8055\ : InMux
    port map (
            O => \N__37863\,
            I => \N__37833\
        );

    \I__8054\ : InMux
    port map (
            O => \N__37862\,
            I => \N__37822\
        );

    \I__8053\ : InMux
    port map (
            O => \N__37861\,
            I => \N__37822\
        );

    \I__8052\ : InMux
    port map (
            O => \N__37860\,
            I => \N__37822\
        );

    \I__8051\ : InMux
    port map (
            O => \N__37859\,
            I => \N__37822\
        );

    \I__8050\ : InMux
    port map (
            O => \N__37858\,
            I => \N__37822\
        );

    \I__8049\ : InMux
    port map (
            O => \N__37855\,
            I => \N__37813\
        );

    \I__8048\ : InMux
    port map (
            O => \N__37852\,
            I => \N__37813\
        );

    \I__8047\ : InMux
    port map (
            O => \N__37849\,
            I => \N__37813\
        );

    \I__8046\ : InMux
    port map (
            O => \N__37846\,
            I => \N__37813\
        );

    \I__8045\ : InMux
    port map (
            O => \N__37845\,
            I => \N__37804\
        );

    \I__8044\ : InMux
    port map (
            O => \N__37844\,
            I => \N__37804\
        );

    \I__8043\ : InMux
    port map (
            O => \N__37843\,
            I => \N__37804\
        );

    \I__8042\ : InMux
    port map (
            O => \N__37842\,
            I => \N__37804\
        );

    \I__8041\ : InMux
    port map (
            O => \N__37841\,
            I => \N__37799\
        );

    \I__8040\ : InMux
    port map (
            O => \N__37840\,
            I => \N__37799\
        );

    \I__8039\ : InMux
    port map (
            O => \N__37839\,
            I => \N__37794\
        );

    \I__8038\ : InMux
    port map (
            O => \N__37838\,
            I => \N__37794\
        );

    \I__8037\ : LocalMux
    port map (
            O => \N__37833\,
            I => \N__37786\
        );

    \I__8036\ : LocalMux
    port map (
            O => \N__37822\,
            I => \N__37786\
        );

    \I__8035\ : LocalMux
    port map (
            O => \N__37813\,
            I => \N__37781\
        );

    \I__8034\ : LocalMux
    port map (
            O => \N__37804\,
            I => \N__37781\
        );

    \I__8033\ : LocalMux
    port map (
            O => \N__37799\,
            I => \N__37775\
        );

    \I__8032\ : LocalMux
    port map (
            O => \N__37794\,
            I => \N__37775\
        );

    \I__8031\ : InMux
    port map (
            O => \N__37793\,
            I => \N__37769\
        );

    \I__8030\ : InMux
    port map (
            O => \N__37792\,
            I => \N__37769\
        );

    \I__8029\ : InMux
    port map (
            O => \N__37791\,
            I => \N__37766\
        );

    \I__8028\ : Span4Mux_h
    port map (
            O => \N__37786\,
            I => \N__37761\
        );

    \I__8027\ : Span4Mux_v
    port map (
            O => \N__37781\,
            I => \N__37761\
        );

    \I__8026\ : InMux
    port map (
            O => \N__37780\,
            I => \N__37758\
        );

    \I__8025\ : Span4Mux_h
    port map (
            O => \N__37775\,
            I => \N__37755\
        );

    \I__8024\ : InMux
    port map (
            O => \N__37774\,
            I => \N__37752\
        );

    \I__8023\ : LocalMux
    port map (
            O => \N__37769\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__8022\ : LocalMux
    port map (
            O => \N__37766\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__8021\ : Odrv4
    port map (
            O => \N__37761\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__8020\ : LocalMux
    port map (
            O => \N__37758\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__8019\ : Odrv4
    port map (
            O => \N__37755\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__8018\ : LocalMux
    port map (
            O => \N__37752\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__8017\ : InMux
    port map (
            O => \N__37739\,
            I => \N__37736\
        );

    \I__8016\ : LocalMux
    port map (
            O => \N__37736\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15\
        );

    \I__8015\ : CascadeMux
    port map (
            O => \N__37733\,
            I => \N__37730\
        );

    \I__8014\ : InMux
    port map (
            O => \N__37730\,
            I => \N__37726\
        );

    \I__8013\ : InMux
    port map (
            O => \N__37729\,
            I => \N__37722\
        );

    \I__8012\ : LocalMux
    port map (
            O => \N__37726\,
            I => \N__37719\
        );

    \I__8011\ : InMux
    port map (
            O => \N__37725\,
            I => \N__37716\
        );

    \I__8010\ : LocalMux
    port map (
            O => \N__37722\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__8009\ : Odrv4
    port map (
            O => \N__37719\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__8008\ : LocalMux
    port map (
            O => \N__37716\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__8007\ : InMux
    port map (
            O => \N__37709\,
            I => \N__37706\
        );

    \I__8006\ : LocalMux
    port map (
            O => \N__37706\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_1\
        );

    \I__8005\ : InMux
    port map (
            O => \N__37703\,
            I => \N__37700\
        );

    \I__8004\ : LocalMux
    port map (
            O => \N__37700\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_19\
        );

    \I__8003\ : CascadeMux
    port map (
            O => \N__37697\,
            I => \N__37694\
        );

    \I__8002\ : InMux
    port map (
            O => \N__37694\,
            I => \N__37691\
        );

    \I__8001\ : LocalMux
    port map (
            O => \N__37691\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_19\
        );

    \I__8000\ : InMux
    port map (
            O => \N__37688\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__7999\ : InMux
    port map (
            O => \N__37685\,
            I => \N__37682\
        );

    \I__7998\ : LocalMux
    port map (
            O => \N__37682\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6\
        );

    \I__7997\ : InMux
    port map (
            O => \N__37679\,
            I => \N__37676\
        );

    \I__7996\ : LocalMux
    port map (
            O => \N__37676\,
            I => \N__37673\
        );

    \I__7995\ : Span4Mux_v
    port map (
            O => \N__37673\,
            I => \N__37670\
        );

    \I__7994\ : Odrv4
    port map (
            O => \N__37670\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0\
        );

    \I__7993\ : InMux
    port map (
            O => \N__37667\,
            I => \N__37664\
        );

    \I__7992\ : LocalMux
    port map (
            O => \N__37664\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7\
        );

    \I__7991\ : InMux
    port map (
            O => \N__37661\,
            I => \N__37658\
        );

    \I__7990\ : LocalMux
    port map (
            O => \N__37658\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8\
        );

    \I__7989\ : InMux
    port map (
            O => \N__37655\,
            I => \N__37652\
        );

    \I__7988\ : LocalMux
    port map (
            O => \N__37652\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9\
        );

    \I__7987\ : InMux
    port map (
            O => \N__37649\,
            I => \N__37646\
        );

    \I__7986\ : LocalMux
    port map (
            O => \N__37646\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2\
        );

    \I__7985\ : CascadeMux
    port map (
            O => \N__37643\,
            I => \N__37640\
        );

    \I__7984\ : InMux
    port map (
            O => \N__37640\,
            I => \N__37637\
        );

    \I__7983\ : LocalMux
    port map (
            O => \N__37637\,
            I => \N__37634\
        );

    \I__7982\ : Span4Mux_h
    port map (
            O => \N__37634\,
            I => \N__37631\
        );

    \I__7981\ : Odrv4
    port map (
            O => \N__37631\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_11\
        );

    \I__7980\ : InMux
    port map (
            O => \N__37628\,
            I => \N__37625\
        );

    \I__7979\ : LocalMux
    port map (
            O => \N__37625\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_11\
        );

    \I__7978\ : CascadeMux
    port map (
            O => \N__37622\,
            I => \N__37619\
        );

    \I__7977\ : InMux
    port map (
            O => \N__37619\,
            I => \N__37616\
        );

    \I__7976\ : LocalMux
    port map (
            O => \N__37616\,
            I => \N__37613\
        );

    \I__7975\ : Odrv4
    port map (
            O => \N__37613\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_12\
        );

    \I__7974\ : InMux
    port map (
            O => \N__37610\,
            I => \N__37607\
        );

    \I__7973\ : LocalMux
    port map (
            O => \N__37607\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_12\
        );

    \I__7972\ : CascadeMux
    port map (
            O => \N__37604\,
            I => \N__37601\
        );

    \I__7971\ : InMux
    port map (
            O => \N__37601\,
            I => \N__37598\
        );

    \I__7970\ : LocalMux
    port map (
            O => \N__37598\,
            I => \N__37595\
        );

    \I__7969\ : Odrv4
    port map (
            O => \N__37595\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_13\
        );

    \I__7968\ : InMux
    port map (
            O => \N__37592\,
            I => \N__37589\
        );

    \I__7967\ : LocalMux
    port map (
            O => \N__37589\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_13\
        );

    \I__7966\ : CascadeMux
    port map (
            O => \N__37586\,
            I => \N__37583\
        );

    \I__7965\ : InMux
    port map (
            O => \N__37583\,
            I => \N__37580\
        );

    \I__7964\ : LocalMux
    port map (
            O => \N__37580\,
            I => \N__37577\
        );

    \I__7963\ : Span4Mux_v
    port map (
            O => \N__37577\,
            I => \N__37574\
        );

    \I__7962\ : Odrv4
    port map (
            O => \N__37574\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_14\
        );

    \I__7961\ : InMux
    port map (
            O => \N__37571\,
            I => \N__37568\
        );

    \I__7960\ : LocalMux
    port map (
            O => \N__37568\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_14\
        );

    \I__7959\ : CascadeMux
    port map (
            O => \N__37565\,
            I => \N__37562\
        );

    \I__7958\ : InMux
    port map (
            O => \N__37562\,
            I => \N__37559\
        );

    \I__7957\ : LocalMux
    port map (
            O => \N__37559\,
            I => \N__37556\
        );

    \I__7956\ : Odrv4
    port map (
            O => \N__37556\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_15\
        );

    \I__7955\ : InMux
    port map (
            O => \N__37553\,
            I => \N__37550\
        );

    \I__7954\ : LocalMux
    port map (
            O => \N__37550\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_15\
        );

    \I__7953\ : CascadeMux
    port map (
            O => \N__37547\,
            I => \N__37544\
        );

    \I__7952\ : InMux
    port map (
            O => \N__37544\,
            I => \N__37541\
        );

    \I__7951\ : LocalMux
    port map (
            O => \N__37541\,
            I => \N__37538\
        );

    \I__7950\ : Span4Mux_h
    port map (
            O => \N__37538\,
            I => \N__37535\
        );

    \I__7949\ : Odrv4
    port map (
            O => \N__37535\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_16\
        );

    \I__7948\ : InMux
    port map (
            O => \N__37532\,
            I => \N__37529\
        );

    \I__7947\ : LocalMux
    port map (
            O => \N__37529\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_16\
        );

    \I__7946\ : CascadeMux
    port map (
            O => \N__37526\,
            I => \N__37523\
        );

    \I__7945\ : InMux
    port map (
            O => \N__37523\,
            I => \N__37520\
        );

    \I__7944\ : LocalMux
    port map (
            O => \N__37520\,
            I => \N__37517\
        );

    \I__7943\ : Span4Mux_h
    port map (
            O => \N__37517\,
            I => \N__37514\
        );

    \I__7942\ : Odrv4
    port map (
            O => \N__37514\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_17\
        );

    \I__7941\ : InMux
    port map (
            O => \N__37511\,
            I => \N__37508\
        );

    \I__7940\ : LocalMux
    port map (
            O => \N__37508\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_17\
        );

    \I__7939\ : CascadeMux
    port map (
            O => \N__37505\,
            I => \N__37502\
        );

    \I__7938\ : InMux
    port map (
            O => \N__37502\,
            I => \N__37499\
        );

    \I__7937\ : LocalMux
    port map (
            O => \N__37499\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_18\
        );

    \I__7936\ : InMux
    port map (
            O => \N__37496\,
            I => \N__37493\
        );

    \I__7935\ : LocalMux
    port map (
            O => \N__37493\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_18\
        );

    \I__7934\ : CascadeMux
    port map (
            O => \N__37490\,
            I => \N__37487\
        );

    \I__7933\ : InMux
    port map (
            O => \N__37487\,
            I => \N__37484\
        );

    \I__7932\ : LocalMux
    port map (
            O => \N__37484\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_4\
        );

    \I__7931\ : InMux
    port map (
            O => \N__37481\,
            I => \N__37478\
        );

    \I__7930\ : LocalMux
    port map (
            O => \N__37478\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_4\
        );

    \I__7929\ : CascadeMux
    port map (
            O => \N__37475\,
            I => \N__37472\
        );

    \I__7928\ : InMux
    port map (
            O => \N__37472\,
            I => \N__37469\
        );

    \I__7927\ : LocalMux
    port map (
            O => \N__37469\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_5\
        );

    \I__7926\ : InMux
    port map (
            O => \N__37466\,
            I => \N__37463\
        );

    \I__7925\ : LocalMux
    port map (
            O => \N__37463\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_5\
        );

    \I__7924\ : CascadeMux
    port map (
            O => \N__37460\,
            I => \N__37457\
        );

    \I__7923\ : InMux
    port map (
            O => \N__37457\,
            I => \N__37454\
        );

    \I__7922\ : LocalMux
    port map (
            O => \N__37454\,
            I => \phase_controller_slave.stoper_hc.target_timeZ1Z_6\
        );

    \I__7921\ : InMux
    port map (
            O => \N__37451\,
            I => \N__37448\
        );

    \I__7920\ : LocalMux
    port map (
            O => \N__37448\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_6\
        );

    \I__7919\ : CascadeMux
    port map (
            O => \N__37445\,
            I => \N__37442\
        );

    \I__7918\ : InMux
    port map (
            O => \N__37442\,
            I => \N__37439\
        );

    \I__7917\ : LocalMux
    port map (
            O => \N__37439\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_7\
        );

    \I__7916\ : InMux
    port map (
            O => \N__37436\,
            I => \N__37433\
        );

    \I__7915\ : LocalMux
    port map (
            O => \N__37433\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_7\
        );

    \I__7914\ : CascadeMux
    port map (
            O => \N__37430\,
            I => \N__37427\
        );

    \I__7913\ : InMux
    port map (
            O => \N__37427\,
            I => \N__37424\
        );

    \I__7912\ : LocalMux
    port map (
            O => \N__37424\,
            I => \N__37421\
        );

    \I__7911\ : Odrv12
    port map (
            O => \N__37421\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_8\
        );

    \I__7910\ : InMux
    port map (
            O => \N__37418\,
            I => \N__37415\
        );

    \I__7909\ : LocalMux
    port map (
            O => \N__37415\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_8\
        );

    \I__7908\ : CascadeMux
    port map (
            O => \N__37412\,
            I => \N__37409\
        );

    \I__7907\ : InMux
    port map (
            O => \N__37409\,
            I => \N__37406\
        );

    \I__7906\ : LocalMux
    port map (
            O => \N__37406\,
            I => \N__37403\
        );

    \I__7905\ : Odrv4
    port map (
            O => \N__37403\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_9\
        );

    \I__7904\ : InMux
    port map (
            O => \N__37400\,
            I => \N__37397\
        );

    \I__7903\ : LocalMux
    port map (
            O => \N__37397\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_9\
        );

    \I__7902\ : CascadeMux
    port map (
            O => \N__37394\,
            I => \N__37391\
        );

    \I__7901\ : InMux
    port map (
            O => \N__37391\,
            I => \N__37388\
        );

    \I__7900\ : LocalMux
    port map (
            O => \N__37388\,
            I => \N__37385\
        );

    \I__7899\ : Odrv4
    port map (
            O => \N__37385\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_10\
        );

    \I__7898\ : InMux
    port map (
            O => \N__37382\,
            I => \N__37379\
        );

    \I__7897\ : LocalMux
    port map (
            O => \N__37379\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_10\
        );

    \I__7896\ : InMux
    port map (
            O => \N__37376\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\
        );

    \I__7895\ : InMux
    port map (
            O => \N__37373\,
            I => \N__37369\
        );

    \I__7894\ : InMux
    port map (
            O => \N__37372\,
            I => \N__37366\
        );

    \I__7893\ : LocalMux
    port map (
            O => \N__37369\,
            I => \N__37363\
        );

    \I__7892\ : LocalMux
    port map (
            O => \N__37366\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__7891\ : Odrv4
    port map (
            O => \N__37363\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__7890\ : CascadeMux
    port map (
            O => \N__37358\,
            I => \N__37355\
        );

    \I__7889\ : InMux
    port map (
            O => \N__37355\,
            I => \N__37352\
        );

    \I__7888\ : LocalMux
    port map (
            O => \N__37352\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16\
        );

    \I__7887\ : InMux
    port map (
            O => \N__37349\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\
        );

    \I__7886\ : InMux
    port map (
            O => \N__37346\,
            I => \N__37342\
        );

    \I__7885\ : InMux
    port map (
            O => \N__37345\,
            I => \N__37339\
        );

    \I__7884\ : LocalMux
    port map (
            O => \N__37342\,
            I => \N__37336\
        );

    \I__7883\ : LocalMux
    port map (
            O => \N__37339\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__7882\ : Odrv4
    port map (
            O => \N__37336\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__7881\ : InMux
    port map (
            O => \N__37331\,
            I => \N__37328\
        );

    \I__7880\ : LocalMux
    port map (
            O => \N__37328\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17\
        );

    \I__7879\ : InMux
    port map (
            O => \N__37325\,
            I => \bfn_15_15_0_\
        );

    \I__7878\ : InMux
    port map (
            O => \N__37322\,
            I => \N__37318\
        );

    \I__7877\ : InMux
    port map (
            O => \N__37321\,
            I => \N__37315\
        );

    \I__7876\ : LocalMux
    port map (
            O => \N__37318\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__7875\ : LocalMux
    port map (
            O => \N__37315\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__7874\ : CascadeMux
    port map (
            O => \N__37310\,
            I => \N__37307\
        );

    \I__7873\ : InMux
    port map (
            O => \N__37307\,
            I => \N__37304\
        );

    \I__7872\ : LocalMux
    port map (
            O => \N__37304\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18\
        );

    \I__7871\ : InMux
    port map (
            O => \N__37301\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\
        );

    \I__7870\ : InMux
    port map (
            O => \N__37298\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17\
        );

    \I__7869\ : CascadeMux
    port map (
            O => \N__37295\,
            I => \N__37292\
        );

    \I__7868\ : InMux
    port map (
            O => \N__37292\,
            I => \N__37289\
        );

    \I__7867\ : LocalMux
    port map (
            O => \N__37289\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_0\
        );

    \I__7866\ : CascadeMux
    port map (
            O => \N__37286\,
            I => \N__37283\
        );

    \I__7865\ : InMux
    port map (
            O => \N__37283\,
            I => \N__37280\
        );

    \I__7864\ : LocalMux
    port map (
            O => \N__37280\,
            I => \N__37277\
        );

    \I__7863\ : Odrv4
    port map (
            O => \N__37277\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_1\
        );

    \I__7862\ : InMux
    port map (
            O => \N__37274\,
            I => \N__37271\
        );

    \I__7861\ : LocalMux
    port map (
            O => \N__37271\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_1\
        );

    \I__7860\ : CascadeMux
    port map (
            O => \N__37268\,
            I => \N__37265\
        );

    \I__7859\ : InMux
    port map (
            O => \N__37265\,
            I => \N__37262\
        );

    \I__7858\ : LocalMux
    port map (
            O => \N__37262\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_2\
        );

    \I__7857\ : InMux
    port map (
            O => \N__37259\,
            I => \N__37256\
        );

    \I__7856\ : LocalMux
    port map (
            O => \N__37256\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_2\
        );

    \I__7855\ : CascadeMux
    port map (
            O => \N__37253\,
            I => \N__37250\
        );

    \I__7854\ : InMux
    port map (
            O => \N__37250\,
            I => \N__37247\
        );

    \I__7853\ : LocalMux
    port map (
            O => \N__37247\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_3\
        );

    \I__7852\ : InMux
    port map (
            O => \N__37244\,
            I => \N__37241\
        );

    \I__7851\ : LocalMux
    port map (
            O => \N__37241\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_3\
        );

    \I__7850\ : InMux
    port map (
            O => \N__37238\,
            I => \N__37235\
        );

    \I__7849\ : LocalMux
    port map (
            O => \N__37235\,
            I => \N__37232\
        );

    \I__7848\ : Span4Mux_h
    port map (
            O => \N__37232\,
            I => \N__37228\
        );

    \I__7847\ : InMux
    port map (
            O => \N__37231\,
            I => \N__37225\
        );

    \I__7846\ : Odrv4
    port map (
            O => \N__37228\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__7845\ : LocalMux
    port map (
            O => \N__37225\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__7844\ : InMux
    port map (
            O => \N__37220\,
            I => \N__37217\
        );

    \I__7843\ : LocalMux
    port map (
            O => \N__37217\,
            I => \N__37214\
        );

    \I__7842\ : Span4Mux_h
    port map (
            O => \N__37214\,
            I => \N__37211\
        );

    \I__7841\ : Odrv4
    port map (
            O => \N__37211\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7\
        );

    \I__7840\ : InMux
    port map (
            O => \N__37208\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\
        );

    \I__7839\ : InMux
    port map (
            O => \N__37205\,
            I => \N__37201\
        );

    \I__7838\ : InMux
    port map (
            O => \N__37204\,
            I => \N__37198\
        );

    \I__7837\ : LocalMux
    port map (
            O => \N__37201\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__7836\ : LocalMux
    port map (
            O => \N__37198\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__7835\ : CascadeMux
    port map (
            O => \N__37193\,
            I => \N__37190\
        );

    \I__7834\ : InMux
    port map (
            O => \N__37190\,
            I => \N__37187\
        );

    \I__7833\ : LocalMux
    port map (
            O => \N__37187\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8\
        );

    \I__7832\ : InMux
    port map (
            O => \N__37184\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\
        );

    \I__7831\ : InMux
    port map (
            O => \N__37181\,
            I => \N__37178\
        );

    \I__7830\ : LocalMux
    port map (
            O => \N__37178\,
            I => \N__37174\
        );

    \I__7829\ : InMux
    port map (
            O => \N__37177\,
            I => \N__37171\
        );

    \I__7828\ : Odrv4
    port map (
            O => \N__37174\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__7827\ : LocalMux
    port map (
            O => \N__37171\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__7826\ : InMux
    port map (
            O => \N__37166\,
            I => \N__37163\
        );

    \I__7825\ : LocalMux
    port map (
            O => \N__37163\,
            I => \N__37160\
        );

    \I__7824\ : Odrv12
    port map (
            O => \N__37160\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9\
        );

    \I__7823\ : InMux
    port map (
            O => \N__37157\,
            I => \bfn_15_14_0_\
        );

    \I__7822\ : InMux
    port map (
            O => \N__37154\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\
        );

    \I__7821\ : InMux
    port map (
            O => \N__37151\,
            I => \N__37148\
        );

    \I__7820\ : LocalMux
    port map (
            O => \N__37148\,
            I => \N__37144\
        );

    \I__7819\ : InMux
    port map (
            O => \N__37147\,
            I => \N__37141\
        );

    \I__7818\ : Odrv4
    port map (
            O => \N__37144\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__7817\ : LocalMux
    port map (
            O => \N__37141\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__7816\ : CascadeMux
    port map (
            O => \N__37136\,
            I => \N__37133\
        );

    \I__7815\ : InMux
    port map (
            O => \N__37133\,
            I => \N__37130\
        );

    \I__7814\ : LocalMux
    port map (
            O => \N__37130\,
            I => \N__37127\
        );

    \I__7813\ : Odrv4
    port map (
            O => \N__37127\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11\
        );

    \I__7812\ : InMux
    port map (
            O => \N__37124\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\
        );

    \I__7811\ : InMux
    port map (
            O => \N__37121\,
            I => \N__37117\
        );

    \I__7810\ : InMux
    port map (
            O => \N__37120\,
            I => \N__37114\
        );

    \I__7809\ : LocalMux
    port map (
            O => \N__37117\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__7808\ : LocalMux
    port map (
            O => \N__37114\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__7807\ : InMux
    port map (
            O => \N__37109\,
            I => \N__37106\
        );

    \I__7806\ : LocalMux
    port map (
            O => \N__37106\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12\
        );

    \I__7805\ : InMux
    port map (
            O => \N__37103\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\
        );

    \I__7804\ : InMux
    port map (
            O => \N__37100\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\
        );

    \I__7803\ : InMux
    port map (
            O => \N__37097\,
            I => \N__37093\
        );

    \I__7802\ : InMux
    port map (
            O => \N__37096\,
            I => \N__37090\
        );

    \I__7801\ : LocalMux
    port map (
            O => \N__37093\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__7800\ : LocalMux
    port map (
            O => \N__37090\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__7799\ : InMux
    port map (
            O => \N__37085\,
            I => \N__37082\
        );

    \I__7798\ : LocalMux
    port map (
            O => \N__37082\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14\
        );

    \I__7797\ : InMux
    port map (
            O => \N__37079\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\
        );

    \I__7796\ : InMux
    port map (
            O => \N__37076\,
            I => \N__37072\
        );

    \I__7795\ : InMux
    port map (
            O => \N__37075\,
            I => \N__37069\
        );

    \I__7794\ : LocalMux
    port map (
            O => \N__37072\,
            I => measured_delay_hc_29
        );

    \I__7793\ : LocalMux
    port map (
            O => \N__37069\,
            I => measured_delay_hc_29
        );

    \I__7792\ : InMux
    port map (
            O => \N__37064\,
            I => \N__37061\
        );

    \I__7791\ : LocalMux
    port map (
            O => \N__37061\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_4\
        );

    \I__7790\ : CascadeMux
    port map (
            O => \N__37058\,
            I => \N__37054\
        );

    \I__7789\ : InMux
    port map (
            O => \N__37057\,
            I => \N__37051\
        );

    \I__7788\ : InMux
    port map (
            O => \N__37054\,
            I => \N__37048\
        );

    \I__7787\ : LocalMux
    port map (
            O => \N__37051\,
            I => measured_delay_hc_27
        );

    \I__7786\ : LocalMux
    port map (
            O => \N__37048\,
            I => measured_delay_hc_27
        );

    \I__7785\ : InMux
    port map (
            O => \N__37043\,
            I => \N__37040\
        );

    \I__7784\ : LocalMux
    port map (
            O => \N__37040\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0\
        );

    \I__7783\ : CascadeMux
    port map (
            O => \N__37037\,
            I => \N__37034\
        );

    \I__7782\ : InMux
    port map (
            O => \N__37034\,
            I => \N__37031\
        );

    \I__7781\ : LocalMux
    port map (
            O => \N__37031\,
            I => \N__37027\
        );

    \I__7780\ : InMux
    port map (
            O => \N__37030\,
            I => \N__37023\
        );

    \I__7779\ : Span4Mux_h
    port map (
            O => \N__37027\,
            I => \N__37020\
        );

    \I__7778\ : InMux
    port map (
            O => \N__37026\,
            I => \N__37017\
        );

    \I__7777\ : LocalMux
    port map (
            O => \N__37023\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__7776\ : Odrv4
    port map (
            O => \N__37020\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__7775\ : LocalMux
    port map (
            O => \N__37017\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__7774\ : InMux
    port map (
            O => \N__37010\,
            I => \N__37006\
        );

    \I__7773\ : InMux
    port map (
            O => \N__37009\,
            I => \N__37003\
        );

    \I__7772\ : LocalMux
    port map (
            O => \N__37006\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__7771\ : LocalMux
    port map (
            O => \N__37003\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__7770\ : CascadeMux
    port map (
            O => \N__36998\,
            I => \N__36995\
        );

    \I__7769\ : InMux
    port map (
            O => \N__36995\,
            I => \N__36992\
        );

    \I__7768\ : LocalMux
    port map (
            O => \N__36992\,
            I => \N__36989\
        );

    \I__7767\ : Span4Mux_h
    port map (
            O => \N__36989\,
            I => \N__36986\
        );

    \I__7766\ : Odrv4
    port map (
            O => \N__36986\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2\
        );

    \I__7765\ : InMux
    port map (
            O => \N__36983\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\
        );

    \I__7764\ : InMux
    port map (
            O => \N__36980\,
            I => \N__36977\
        );

    \I__7763\ : LocalMux
    port map (
            O => \N__36977\,
            I => \N__36974\
        );

    \I__7762\ : Span4Mux_v
    port map (
            O => \N__36974\,
            I => \N__36971\
        );

    \I__7761\ : Odrv4
    port map (
            O => \N__36971\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0\
        );

    \I__7760\ : CascadeMux
    port map (
            O => \N__36968\,
            I => \N__36965\
        );

    \I__7759\ : InMux
    port map (
            O => \N__36965\,
            I => \N__36961\
        );

    \I__7758\ : InMux
    port map (
            O => \N__36964\,
            I => \N__36958\
        );

    \I__7757\ : LocalMux
    port map (
            O => \N__36961\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__7756\ : LocalMux
    port map (
            O => \N__36958\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__7755\ : InMux
    port map (
            O => \N__36953\,
            I => \N__36950\
        );

    \I__7754\ : LocalMux
    port map (
            O => \N__36950\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3\
        );

    \I__7753\ : InMux
    port map (
            O => \N__36947\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\
        );

    \I__7752\ : InMux
    port map (
            O => \N__36944\,
            I => \N__36941\
        );

    \I__7751\ : LocalMux
    port map (
            O => \N__36941\,
            I => \N__36938\
        );

    \I__7750\ : Span4Mux_v
    port map (
            O => \N__36938\,
            I => \N__36934\
        );

    \I__7749\ : InMux
    port map (
            O => \N__36937\,
            I => \N__36931\
        );

    \I__7748\ : Odrv4
    port map (
            O => \N__36934\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__7747\ : LocalMux
    port map (
            O => \N__36931\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__7746\ : CascadeMux
    port map (
            O => \N__36926\,
            I => \N__36923\
        );

    \I__7745\ : InMux
    port map (
            O => \N__36923\,
            I => \N__36920\
        );

    \I__7744\ : LocalMux
    port map (
            O => \N__36920\,
            I => \N__36917\
        );

    \I__7743\ : Span4Mux_h
    port map (
            O => \N__36917\,
            I => \N__36914\
        );

    \I__7742\ : Odrv4
    port map (
            O => \N__36914\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4\
        );

    \I__7741\ : InMux
    port map (
            O => \N__36911\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\
        );

    \I__7740\ : InMux
    port map (
            O => \N__36908\,
            I => \N__36905\
        );

    \I__7739\ : LocalMux
    port map (
            O => \N__36905\,
            I => \N__36902\
        );

    \I__7738\ : Span4Mux_h
    port map (
            O => \N__36902\,
            I => \N__36898\
        );

    \I__7737\ : InMux
    port map (
            O => \N__36901\,
            I => \N__36895\
        );

    \I__7736\ : Odrv4
    port map (
            O => \N__36898\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__7735\ : LocalMux
    port map (
            O => \N__36895\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__7734\ : InMux
    port map (
            O => \N__36890\,
            I => \N__36887\
        );

    \I__7733\ : LocalMux
    port map (
            O => \N__36887\,
            I => \N__36884\
        );

    \I__7732\ : Span4Mux_v
    port map (
            O => \N__36884\,
            I => \N__36881\
        );

    \I__7731\ : Odrv4
    port map (
            O => \N__36881\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5\
        );

    \I__7730\ : InMux
    port map (
            O => \N__36878\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\
        );

    \I__7729\ : InMux
    port map (
            O => \N__36875\,
            I => \N__36871\
        );

    \I__7728\ : InMux
    port map (
            O => \N__36874\,
            I => \N__36868\
        );

    \I__7727\ : LocalMux
    port map (
            O => \N__36871\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__7726\ : LocalMux
    port map (
            O => \N__36868\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__7725\ : CascadeMux
    port map (
            O => \N__36863\,
            I => \N__36860\
        );

    \I__7724\ : InMux
    port map (
            O => \N__36860\,
            I => \N__36857\
        );

    \I__7723\ : LocalMux
    port map (
            O => \N__36857\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6\
        );

    \I__7722\ : InMux
    port map (
            O => \N__36854\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\
        );

    \I__7721\ : CascadeMux
    port map (
            O => \N__36851\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto6_c_cascade_\
        );

    \I__7720\ : CascadeMux
    port map (
            O => \N__36848\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto6_0_0_cascade_\
        );

    \I__7719\ : InMux
    port map (
            O => \N__36845\,
            I => \N__36842\
        );

    \I__7718\ : LocalMux
    port map (
            O => \N__36842\,
            I => \N__36839\
        );

    \I__7717\ : Span12Mux_v
    port map (
            O => \N__36839\,
            I => \N__36836\
        );

    \I__7716\ : Odrv12
    port map (
            O => \N__36836\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt13\
        );

    \I__7715\ : CascadeMux
    port map (
            O => \N__36833\,
            I => \N__36830\
        );

    \I__7714\ : InMux
    port map (
            O => \N__36830\,
            I => \N__36827\
        );

    \I__7713\ : LocalMux
    port map (
            O => \N__36827\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt9\
        );

    \I__7712\ : InMux
    port map (
            O => \N__36824\,
            I => \N__36820\
        );

    \I__7711\ : InMux
    port map (
            O => \N__36823\,
            I => \N__36816\
        );

    \I__7710\ : LocalMux
    port map (
            O => \N__36820\,
            I => \N__36813\
        );

    \I__7709\ : InMux
    port map (
            O => \N__36819\,
            I => \N__36810\
        );

    \I__7708\ : LocalMux
    port map (
            O => \N__36816\,
            I => \N__36805\
        );

    \I__7707\ : Span12Mux_s10_h
    port map (
            O => \N__36813\,
            I => \N__36805\
        );

    \I__7706\ : LocalMux
    port map (
            O => \N__36810\,
            I => measured_delay_hc_21
        );

    \I__7705\ : Odrv12
    port map (
            O => \N__36805\,
            I => measured_delay_hc_21
        );

    \I__7704\ : InMux
    port map (
            O => \N__36800\,
            I => \N__36796\
        );

    \I__7703\ : InMux
    port map (
            O => \N__36799\,
            I => \N__36793\
        );

    \I__7702\ : LocalMux
    port map (
            O => \N__36796\,
            I => \N__36789\
        );

    \I__7701\ : LocalMux
    port map (
            O => \N__36793\,
            I => \N__36786\
        );

    \I__7700\ : InMux
    port map (
            O => \N__36792\,
            I => \N__36783\
        );

    \I__7699\ : Span12Mux_v
    port map (
            O => \N__36789\,
            I => \N__36780\
        );

    \I__7698\ : Span4Mux_v
    port map (
            O => \N__36786\,
            I => \N__36777\
        );

    \I__7697\ : LocalMux
    port map (
            O => \N__36783\,
            I => \N__36774\
        );

    \I__7696\ : Odrv12
    port map (
            O => \N__36780\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1\
        );

    \I__7695\ : Odrv4
    port map (
            O => \N__36777\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1\
        );

    \I__7694\ : Odrv4
    port map (
            O => \N__36774\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1\
        );

    \I__7693\ : CascadeMux
    port map (
            O => \N__36767\,
            I => \N__36764\
        );

    \I__7692\ : InMux
    port map (
            O => \N__36764\,
            I => \N__36759\
        );

    \I__7691\ : InMux
    port map (
            O => \N__36763\,
            I => \N__36754\
        );

    \I__7690\ : InMux
    port map (
            O => \N__36762\,
            I => \N__36754\
        );

    \I__7689\ : LocalMux
    port map (
            O => \N__36759\,
            I => \N__36751\
        );

    \I__7688\ : LocalMux
    port map (
            O => \N__36754\,
            I => measured_delay_hc_20
        );

    \I__7687\ : Odrv4
    port map (
            O => \N__36751\,
            I => measured_delay_hc_20
        );

    \I__7686\ : CascadeMux
    port map (
            O => \N__36746\,
            I => \N__36743\
        );

    \I__7685\ : InMux
    port map (
            O => \N__36743\,
            I => \N__36738\
        );

    \I__7684\ : InMux
    port map (
            O => \N__36742\,
            I => \N__36733\
        );

    \I__7683\ : InMux
    port map (
            O => \N__36741\,
            I => \N__36733\
        );

    \I__7682\ : LocalMux
    port map (
            O => \N__36738\,
            I => measured_delay_hc_19
        );

    \I__7681\ : LocalMux
    port map (
            O => \N__36733\,
            I => measured_delay_hc_19
        );

    \I__7680\ : CascadeMux
    port map (
            O => \N__36728\,
            I => \N__36725\
        );

    \I__7679\ : InMux
    port map (
            O => \N__36725\,
            I => \N__36720\
        );

    \I__7678\ : InMux
    port map (
            O => \N__36724\,
            I => \N__36717\
        );

    \I__7677\ : InMux
    port map (
            O => \N__36723\,
            I => \N__36714\
        );

    \I__7676\ : LocalMux
    port map (
            O => \N__36720\,
            I => \N__36709\
        );

    \I__7675\ : LocalMux
    port map (
            O => \N__36717\,
            I => \N__36709\
        );

    \I__7674\ : LocalMux
    port map (
            O => \N__36714\,
            I => measured_delay_hc_22
        );

    \I__7673\ : Odrv4
    port map (
            O => \N__36709\,
            I => measured_delay_hc_22
        );

    \I__7672\ : InMux
    port map (
            O => \N__36704\,
            I => \N__36701\
        );

    \I__7671\ : LocalMux
    port map (
            O => \N__36701\,
            I => \N__36693\
        );

    \I__7670\ : InMux
    port map (
            O => \N__36700\,
            I => \N__36686\
        );

    \I__7669\ : InMux
    port map (
            O => \N__36699\,
            I => \N__36686\
        );

    \I__7668\ : InMux
    port map (
            O => \N__36698\,
            I => \N__36686\
        );

    \I__7667\ : InMux
    port map (
            O => \N__36697\,
            I => \N__36681\
        );

    \I__7666\ : InMux
    port map (
            O => \N__36696\,
            I => \N__36681\
        );

    \I__7665\ : Span4Mux_v
    port map (
            O => \N__36693\,
            I => \N__36676\
        );

    \I__7664\ : LocalMux
    port map (
            O => \N__36686\,
            I => \N__36676\
        );

    \I__7663\ : LocalMux
    port map (
            O => \N__36681\,
            I => \N__36673\
        );

    \I__7662\ : Span4Mux_h
    port map (
            O => \N__36676\,
            I => \N__36670\
        );

    \I__7661\ : Span4Mux_v
    port map (
            O => \N__36673\,
            I => \N__36667\
        );

    \I__7660\ : Span4Mux_v
    port map (
            O => \N__36670\,
            I => \N__36664\
        );

    \I__7659\ : Span4Mux_h
    port map (
            O => \N__36667\,
            I => \N__36661\
        );

    \I__7658\ : Span4Mux_h
    port map (
            O => \N__36664\,
            I => \N__36658\
        );

    \I__7657\ : Span4Mux_h
    port map (
            O => \N__36661\,
            I => \N__36655\
        );

    \I__7656\ : Odrv4
    port map (
            O => \N__36658\,
            I => \delay_measurement_inst.delay_hc_reg3lto31_0_0\
        );

    \I__7655\ : Odrv4
    port map (
            O => \N__36655\,
            I => \delay_measurement_inst.delay_hc_reg3lto31_0_0\
        );

    \I__7654\ : CascadeMux
    port map (
            O => \N__36650\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6_cascade_\
        );

    \I__7653\ : InMux
    port map (
            O => \N__36647\,
            I => \N__36642\
        );

    \I__7652\ : InMux
    port map (
            O => \N__36646\,
            I => \N__36637\
        );

    \I__7651\ : InMux
    port map (
            O => \N__36645\,
            I => \N__36637\
        );

    \I__7650\ : LocalMux
    port map (
            O => \N__36642\,
            I => \N__36634\
        );

    \I__7649\ : LocalMux
    port map (
            O => \N__36637\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__7648\ : Odrv4
    port map (
            O => \N__36634\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__7647\ : InMux
    port map (
            O => \N__36629\,
            I => \N__36626\
        );

    \I__7646\ : LocalMux
    port map (
            O => \N__36626\,
            I => \N__36623\
        );

    \I__7645\ : Odrv4
    port map (
            O => \N__36623\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9\
        );

    \I__7644\ : InMux
    port map (
            O => \N__36620\,
            I => \N__36617\
        );

    \I__7643\ : LocalMux
    port map (
            O => \N__36617\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_12\
        );

    \I__7642\ : InMux
    port map (
            O => \N__36614\,
            I => \N__36611\
        );

    \I__7641\ : LocalMux
    port map (
            O => \N__36611\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_11\
        );

    \I__7640\ : InMux
    port map (
            O => \N__36608\,
            I => \N__36605\
        );

    \I__7639\ : LocalMux
    port map (
            O => \N__36605\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt15_0\
        );

    \I__7638\ : CascadeMux
    port map (
            O => \N__36602\,
            I => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_3_cascade_\
        );

    \I__7637\ : InMux
    port map (
            O => \N__36599\,
            I => \N__36593\
        );

    \I__7636\ : InMux
    port map (
            O => \N__36598\,
            I => \N__36590\
        );

    \I__7635\ : InMux
    port map (
            O => \N__36597\,
            I => \N__36585\
        );

    \I__7634\ : InMux
    port map (
            O => \N__36596\,
            I => \N__36585\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__36593\,
            I => \N__36582\
        );

    \I__7632\ : LocalMux
    port map (
            O => \N__36590\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__7631\ : LocalMux
    port map (
            O => \N__36585\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__7630\ : Odrv4
    port map (
            O => \N__36582\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__7629\ : InMux
    port map (
            O => \N__36575\,
            I => \N__36570\
        );

    \I__7628\ : InMux
    port map (
            O => \N__36574\,
            I => \N__36567\
        );

    \I__7627\ : InMux
    port map (
            O => \N__36573\,
            I => \N__36564\
        );

    \I__7626\ : LocalMux
    port map (
            O => \N__36570\,
            I => \delay_measurement_inst.prev_hc_sigZ0\
        );

    \I__7625\ : LocalMux
    port map (
            O => \N__36567\,
            I => \delay_measurement_inst.prev_hc_sigZ0\
        );

    \I__7624\ : LocalMux
    port map (
            O => \N__36564\,
            I => \delay_measurement_inst.prev_hc_sigZ0\
        );

    \I__7623\ : InMux
    port map (
            O => \N__36557\,
            I => \N__36554\
        );

    \I__7622\ : LocalMux
    port map (
            O => \N__36554\,
            I => \N__36549\
        );

    \I__7621\ : InMux
    port map (
            O => \N__36553\,
            I => \N__36546\
        );

    \I__7620\ : InMux
    port map (
            O => \N__36552\,
            I => \N__36543\
        );

    \I__7619\ : Odrv4
    port map (
            O => \N__36549\,
            I => \delay_measurement_inst.hc_stateZ0Z_0\
        );

    \I__7618\ : LocalMux
    port map (
            O => \N__36546\,
            I => \delay_measurement_inst.hc_stateZ0Z_0\
        );

    \I__7617\ : LocalMux
    port map (
            O => \N__36543\,
            I => \delay_measurement_inst.hc_stateZ0Z_0\
        );

    \I__7616\ : InMux
    port map (
            O => \N__36536\,
            I => \N__36531\
        );

    \I__7615\ : InMux
    port map (
            O => \N__36535\,
            I => \N__36526\
        );

    \I__7614\ : InMux
    port map (
            O => \N__36534\,
            I => \N__36526\
        );

    \I__7613\ : LocalMux
    port map (
            O => \N__36531\,
            I => \N__36520\
        );

    \I__7612\ : LocalMux
    port map (
            O => \N__36526\,
            I => \N__36520\
        );

    \I__7611\ : InMux
    port map (
            O => \N__36525\,
            I => \N__36517\
        );

    \I__7610\ : Odrv4
    port map (
            O => \N__36520\,
            I => delay_tr_d2
        );

    \I__7609\ : LocalMux
    port map (
            O => \N__36517\,
            I => delay_tr_d2
        );

    \I__7608\ : InMux
    port map (
            O => \N__36512\,
            I => \N__36509\
        );

    \I__7607\ : LocalMux
    port map (
            O => \N__36509\,
            I => \N__36504\
        );

    \I__7606\ : InMux
    port map (
            O => \N__36508\,
            I => \N__36501\
        );

    \I__7605\ : InMux
    port map (
            O => \N__36507\,
            I => \N__36498\
        );

    \I__7604\ : Odrv4
    port map (
            O => \N__36504\,
            I => \delay_measurement_inst.tr_stateZ0Z_0\
        );

    \I__7603\ : LocalMux
    port map (
            O => \N__36501\,
            I => \delay_measurement_inst.tr_stateZ0Z_0\
        );

    \I__7602\ : LocalMux
    port map (
            O => \N__36498\,
            I => \delay_measurement_inst.tr_stateZ0Z_0\
        );

    \I__7601\ : InMux
    port map (
            O => \N__36491\,
            I => \N__36486\
        );

    \I__7600\ : InMux
    port map (
            O => \N__36490\,
            I => \N__36483\
        );

    \I__7599\ : InMux
    port map (
            O => \N__36489\,
            I => \N__36480\
        );

    \I__7598\ : LocalMux
    port map (
            O => \N__36486\,
            I => \delay_measurement_inst.prev_tr_sigZ0\
        );

    \I__7597\ : LocalMux
    port map (
            O => \N__36483\,
            I => \delay_measurement_inst.prev_tr_sigZ0\
        );

    \I__7596\ : LocalMux
    port map (
            O => \N__36480\,
            I => \delay_measurement_inst.prev_tr_sigZ0\
        );

    \I__7595\ : InMux
    port map (
            O => \N__36473\,
            I => \N__36470\
        );

    \I__7594\ : LocalMux
    port map (
            O => \N__36470\,
            I => \N__36467\
        );

    \I__7593\ : Span4Mux_h
    port map (
            O => \N__36467\,
            I => \N__36464\
        );

    \I__7592\ : Sp12to4
    port map (
            O => \N__36464\,
            I => \N__36461\
        );

    \I__7591\ : Odrv12
    port map (
            O => \N__36461\,
            I => delay_hc_input_c
        );

    \I__7590\ : InMux
    port map (
            O => \N__36458\,
            I => \N__36455\
        );

    \I__7589\ : LocalMux
    port map (
            O => \N__36455\,
            I => delay_hc_d1
        );

    \I__7588\ : InMux
    port map (
            O => \N__36452\,
            I => \N__36448\
        );

    \I__7587\ : InMux
    port map (
            O => \N__36451\,
            I => \N__36445\
        );

    \I__7586\ : LocalMux
    port map (
            O => \N__36448\,
            I => \N__36442\
        );

    \I__7585\ : LocalMux
    port map (
            O => \N__36445\,
            I => \N__36437\
        );

    \I__7584\ : Span4Mux_h
    port map (
            O => \N__36442\,
            I => \N__36434\
        );

    \I__7583\ : InMux
    port map (
            O => \N__36441\,
            I => \N__36431\
        );

    \I__7582\ : InMux
    port map (
            O => \N__36440\,
            I => \N__36428\
        );

    \I__7581\ : Odrv4
    port map (
            O => \N__36437\,
            I => delay_hc_d2
        );

    \I__7580\ : Odrv4
    port map (
            O => \N__36434\,
            I => delay_hc_d2
        );

    \I__7579\ : LocalMux
    port map (
            O => \N__36431\,
            I => delay_hc_d2
        );

    \I__7578\ : LocalMux
    port map (
            O => \N__36428\,
            I => delay_hc_d2
        );

    \I__7577\ : CascadeMux
    port map (
            O => \N__36419\,
            I => \N__36414\
        );

    \I__7576\ : InMux
    port map (
            O => \N__36418\,
            I => \N__36410\
        );

    \I__7575\ : InMux
    port map (
            O => \N__36417\,
            I => \N__36407\
        );

    \I__7574\ : InMux
    port map (
            O => \N__36414\,
            I => \N__36404\
        );

    \I__7573\ : CascadeMux
    port map (
            O => \N__36413\,
            I => \N__36400\
        );

    \I__7572\ : LocalMux
    port map (
            O => \N__36410\,
            I => \N__36397\
        );

    \I__7571\ : LocalMux
    port map (
            O => \N__36407\,
            I => \N__36394\
        );

    \I__7570\ : LocalMux
    port map (
            O => \N__36404\,
            I => \N__36391\
        );

    \I__7569\ : InMux
    port map (
            O => \N__36403\,
            I => \N__36388\
        );

    \I__7568\ : InMux
    port map (
            O => \N__36400\,
            I => \N__36385\
        );

    \I__7567\ : Span12Mux_s11_h
    port map (
            O => \N__36397\,
            I => \N__36382\
        );

    \I__7566\ : Sp12to4
    port map (
            O => \N__36394\,
            I => \N__36379\
        );

    \I__7565\ : Span4Mux_v
    port map (
            O => \N__36391\,
            I => \N__36374\
        );

    \I__7564\ : LocalMux
    port map (
            O => \N__36388\,
            I => \N__36374\
        );

    \I__7563\ : LocalMux
    port map (
            O => \N__36385\,
            I => measured_delay_hc_9
        );

    \I__7562\ : Odrv12
    port map (
            O => \N__36382\,
            I => measured_delay_hc_9
        );

    \I__7561\ : Odrv12
    port map (
            O => \N__36379\,
            I => measured_delay_hc_9
        );

    \I__7560\ : Odrv4
    port map (
            O => \N__36374\,
            I => measured_delay_hc_9
        );

    \I__7559\ : InMux
    port map (
            O => \N__36365\,
            I => \N__36361\
        );

    \I__7558\ : InMux
    port map (
            O => \N__36364\,
            I => \N__36358\
        );

    \I__7557\ : LocalMux
    port map (
            O => \N__36361\,
            I => \N__36353\
        );

    \I__7556\ : LocalMux
    port map (
            O => \N__36358\,
            I => \N__36353\
        );

    \I__7555\ : Odrv4
    port map (
            O => \N__36353\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__7554\ : InMux
    port map (
            O => \N__36350\,
            I => \N__36347\
        );

    \I__7553\ : LocalMux
    port map (
            O => \N__36347\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18\
        );

    \I__7552\ : InMux
    port map (
            O => \N__36344\,
            I => \N__36341\
        );

    \I__7551\ : LocalMux
    port map (
            O => \N__36341\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14\
        );

    \I__7550\ : InMux
    port map (
            O => \N__36338\,
            I => \N__36335\
        );

    \I__7549\ : LocalMux
    port map (
            O => \N__36335\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11\
        );

    \I__7548\ : InMux
    port map (
            O => \N__36332\,
            I => \N__36329\
        );

    \I__7547\ : LocalMux
    port map (
            O => \N__36329\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13\
        );

    \I__7546\ : InMux
    port map (
            O => \N__36326\,
            I => \N__36312\
        );

    \I__7545\ : InMux
    port map (
            O => \N__36325\,
            I => \N__36295\
        );

    \I__7544\ : InMux
    port map (
            O => \N__36324\,
            I => \N__36295\
        );

    \I__7543\ : InMux
    port map (
            O => \N__36323\,
            I => \N__36295\
        );

    \I__7542\ : InMux
    port map (
            O => \N__36322\,
            I => \N__36295\
        );

    \I__7541\ : InMux
    port map (
            O => \N__36321\,
            I => \N__36295\
        );

    \I__7540\ : InMux
    port map (
            O => \N__36320\,
            I => \N__36295\
        );

    \I__7539\ : InMux
    port map (
            O => \N__36319\,
            I => \N__36295\
        );

    \I__7538\ : InMux
    port map (
            O => \N__36318\,
            I => \N__36295\
        );

    \I__7537\ : InMux
    port map (
            O => \N__36317\,
            I => \N__36280\
        );

    \I__7536\ : InMux
    port map (
            O => \N__36316\,
            I => \N__36280\
        );

    \I__7535\ : InMux
    port map (
            O => \N__36315\,
            I => \N__36280\
        );

    \I__7534\ : LocalMux
    port map (
            O => \N__36312\,
            I => \N__36273\
        );

    \I__7533\ : LocalMux
    port map (
            O => \N__36295\,
            I => \N__36273\
        );

    \I__7532\ : InMux
    port map (
            O => \N__36294\,
            I => \N__36256\
        );

    \I__7531\ : InMux
    port map (
            O => \N__36293\,
            I => \N__36256\
        );

    \I__7530\ : InMux
    port map (
            O => \N__36292\,
            I => \N__36256\
        );

    \I__7529\ : InMux
    port map (
            O => \N__36291\,
            I => \N__36256\
        );

    \I__7528\ : InMux
    port map (
            O => \N__36290\,
            I => \N__36256\
        );

    \I__7527\ : InMux
    port map (
            O => \N__36289\,
            I => \N__36256\
        );

    \I__7526\ : InMux
    port map (
            O => \N__36288\,
            I => \N__36256\
        );

    \I__7525\ : InMux
    port map (
            O => \N__36287\,
            I => \N__36256\
        );

    \I__7524\ : LocalMux
    port map (
            O => \N__36280\,
            I => \N__36252\
        );

    \I__7523\ : InMux
    port map (
            O => \N__36279\,
            I => \N__36249\
        );

    \I__7522\ : InMux
    port map (
            O => \N__36278\,
            I => \N__36246\
        );

    \I__7521\ : Span4Mux_v
    port map (
            O => \N__36273\,
            I => \N__36240\
        );

    \I__7520\ : LocalMux
    port map (
            O => \N__36256\,
            I => \N__36240\
        );

    \I__7519\ : InMux
    port map (
            O => \N__36255\,
            I => \N__36237\
        );

    \I__7518\ : Span4Mux_h
    port map (
            O => \N__36252\,
            I => \N__36232\
        );

    \I__7517\ : LocalMux
    port map (
            O => \N__36249\,
            I => \N__36232\
        );

    \I__7516\ : LocalMux
    port map (
            O => \N__36246\,
            I => \N__36229\
        );

    \I__7515\ : InMux
    port map (
            O => \N__36245\,
            I => \N__36226\
        );

    \I__7514\ : Span4Mux_v
    port map (
            O => \N__36240\,
            I => \N__36223\
        );

    \I__7513\ : LocalMux
    port map (
            O => \N__36237\,
            I => \N__36216\
        );

    \I__7512\ : Sp12to4
    port map (
            O => \N__36232\,
            I => \N__36216\
        );

    \I__7511\ : Sp12to4
    port map (
            O => \N__36229\,
            I => \N__36216\
        );

    \I__7510\ : LocalMux
    port map (
            O => \N__36226\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__7509\ : Odrv4
    port map (
            O => \N__36223\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__7508\ : Odrv12
    port map (
            O => \N__36216\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__7507\ : CascadeMux
    port map (
            O => \N__36209\,
            I => \N__36201\
        );

    \I__7506\ : CascadeMux
    port map (
            O => \N__36208\,
            I => \N__36198\
        );

    \I__7505\ : CascadeMux
    port map (
            O => \N__36207\,
            I => \N__36194\
        );

    \I__7504\ : CascadeMux
    port map (
            O => \N__36206\,
            I => \N__36188\
        );

    \I__7503\ : CascadeMux
    port map (
            O => \N__36205\,
            I => \N__36185\
        );

    \I__7502\ : CascadeMux
    port map (
            O => \N__36204\,
            I => \N__36177\
        );

    \I__7501\ : InMux
    port map (
            O => \N__36201\,
            I => \N__36173\
        );

    \I__7500\ : InMux
    port map (
            O => \N__36198\,
            I => \N__36156\
        );

    \I__7499\ : InMux
    port map (
            O => \N__36197\,
            I => \N__36156\
        );

    \I__7498\ : InMux
    port map (
            O => \N__36194\,
            I => \N__36156\
        );

    \I__7497\ : InMux
    port map (
            O => \N__36193\,
            I => \N__36156\
        );

    \I__7496\ : InMux
    port map (
            O => \N__36192\,
            I => \N__36156\
        );

    \I__7495\ : InMux
    port map (
            O => \N__36191\,
            I => \N__36156\
        );

    \I__7494\ : InMux
    port map (
            O => \N__36188\,
            I => \N__36156\
        );

    \I__7493\ : InMux
    port map (
            O => \N__36185\,
            I => \N__36156\
        );

    \I__7492\ : CascadeMux
    port map (
            O => \N__36184\,
            I => \N__36152\
        );

    \I__7491\ : CascadeMux
    port map (
            O => \N__36183\,
            I => \N__36149\
        );

    \I__7490\ : CascadeMux
    port map (
            O => \N__36182\,
            I => \N__36145\
        );

    \I__7489\ : CascadeMux
    port map (
            O => \N__36181\,
            I => \N__36140\
        );

    \I__7488\ : CascadeMux
    port map (
            O => \N__36180\,
            I => \N__36137\
        );

    \I__7487\ : InMux
    port map (
            O => \N__36177\,
            I => \N__36134\
        );

    \I__7486\ : CascadeMux
    port map (
            O => \N__36176\,
            I => \N__36131\
        );

    \I__7485\ : LocalMux
    port map (
            O => \N__36173\,
            I => \N__36126\
        );

    \I__7484\ : LocalMux
    port map (
            O => \N__36156\,
            I => \N__36126\
        );

    \I__7483\ : InMux
    port map (
            O => \N__36155\,
            I => \N__36109\
        );

    \I__7482\ : InMux
    port map (
            O => \N__36152\,
            I => \N__36109\
        );

    \I__7481\ : InMux
    port map (
            O => \N__36149\,
            I => \N__36109\
        );

    \I__7480\ : InMux
    port map (
            O => \N__36148\,
            I => \N__36109\
        );

    \I__7479\ : InMux
    port map (
            O => \N__36145\,
            I => \N__36109\
        );

    \I__7478\ : InMux
    port map (
            O => \N__36144\,
            I => \N__36109\
        );

    \I__7477\ : InMux
    port map (
            O => \N__36143\,
            I => \N__36109\
        );

    \I__7476\ : InMux
    port map (
            O => \N__36140\,
            I => \N__36109\
        );

    \I__7475\ : InMux
    port map (
            O => \N__36137\,
            I => \N__36106\
        );

    \I__7474\ : LocalMux
    port map (
            O => \N__36134\,
            I => \N__36099\
        );

    \I__7473\ : InMux
    port map (
            O => \N__36131\,
            I => \N__36096\
        );

    \I__7472\ : Span4Mux_v
    port map (
            O => \N__36126\,
            I => \N__36091\
        );

    \I__7471\ : LocalMux
    port map (
            O => \N__36109\,
            I => \N__36091\
        );

    \I__7470\ : LocalMux
    port map (
            O => \N__36106\,
            I => \N__36088\
        );

    \I__7469\ : InMux
    port map (
            O => \N__36105\,
            I => \N__36081\
        );

    \I__7468\ : InMux
    port map (
            O => \N__36104\,
            I => \N__36081\
        );

    \I__7467\ : InMux
    port map (
            O => \N__36103\,
            I => \N__36081\
        );

    \I__7466\ : InMux
    port map (
            O => \N__36102\,
            I => \N__36078\
        );

    \I__7465\ : Odrv12
    port map (
            O => \N__36099\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__7464\ : LocalMux
    port map (
            O => \N__36096\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__7463\ : Odrv4
    port map (
            O => \N__36091\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__7462\ : Odrv4
    port map (
            O => \N__36088\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__7461\ : LocalMux
    port map (
            O => \N__36081\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__7460\ : LocalMux
    port map (
            O => \N__36078\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__7459\ : InMux
    port map (
            O => \N__36065\,
            I => \N__36057\
        );

    \I__7458\ : CascadeMux
    port map (
            O => \N__36064\,
            I => \N__36047\
        );

    \I__7457\ : CascadeMux
    port map (
            O => \N__36063\,
            I => \N__36044\
        );

    \I__7456\ : CascadeMux
    port map (
            O => \N__36062\,
            I => \N__36041\
        );

    \I__7455\ : CascadeMux
    port map (
            O => \N__36061\,
            I => \N__36038\
        );

    \I__7454\ : InMux
    port map (
            O => \N__36060\,
            I => \N__36031\
        );

    \I__7453\ : LocalMux
    port map (
            O => \N__36057\,
            I => \N__36028\
        );

    \I__7452\ : CascadeMux
    port map (
            O => \N__36056\,
            I => \N__36025\
        );

    \I__7451\ : CascadeMux
    port map (
            O => \N__36055\,
            I => \N__36022\
        );

    \I__7450\ : InMux
    port map (
            O => \N__36054\,
            I => \N__36018\
        );

    \I__7449\ : CascadeMux
    port map (
            O => \N__36053\,
            I => \N__36013\
        );

    \I__7448\ : CascadeMux
    port map (
            O => \N__36052\,
            I => \N__36010\
        );

    \I__7447\ : CascadeMux
    port map (
            O => \N__36051\,
            I => \N__36007\
        );

    \I__7446\ : CascadeMux
    port map (
            O => \N__36050\,
            I => \N__36004\
        );

    \I__7445\ : InMux
    port map (
            O => \N__36047\,
            I => \N__35991\
        );

    \I__7444\ : InMux
    port map (
            O => \N__36044\,
            I => \N__35991\
        );

    \I__7443\ : InMux
    port map (
            O => \N__36041\,
            I => \N__35991\
        );

    \I__7442\ : InMux
    port map (
            O => \N__36038\,
            I => \N__35991\
        );

    \I__7441\ : InMux
    port map (
            O => \N__36037\,
            I => \N__35982\
        );

    \I__7440\ : InMux
    port map (
            O => \N__36036\,
            I => \N__35982\
        );

    \I__7439\ : InMux
    port map (
            O => \N__36035\,
            I => \N__35982\
        );

    \I__7438\ : InMux
    port map (
            O => \N__36034\,
            I => \N__35982\
        );

    \I__7437\ : LocalMux
    port map (
            O => \N__36031\,
            I => \N__35979\
        );

    \I__7436\ : Span4Mux_v
    port map (
            O => \N__36028\,
            I => \N__35976\
        );

    \I__7435\ : InMux
    port map (
            O => \N__36025\,
            I => \N__35969\
        );

    \I__7434\ : InMux
    port map (
            O => \N__36022\,
            I => \N__35969\
        );

    \I__7433\ : InMux
    port map (
            O => \N__36021\,
            I => \N__35969\
        );

    \I__7432\ : LocalMux
    port map (
            O => \N__36018\,
            I => \N__35966\
        );

    \I__7431\ : InMux
    port map (
            O => \N__36017\,
            I => \N__35963\
        );

    \I__7430\ : InMux
    port map (
            O => \N__36016\,
            I => \N__35960\
        );

    \I__7429\ : InMux
    port map (
            O => \N__36013\,
            I => \N__35951\
        );

    \I__7428\ : InMux
    port map (
            O => \N__36010\,
            I => \N__35951\
        );

    \I__7427\ : InMux
    port map (
            O => \N__36007\,
            I => \N__35951\
        );

    \I__7426\ : InMux
    port map (
            O => \N__36004\,
            I => \N__35951\
        );

    \I__7425\ : InMux
    port map (
            O => \N__36003\,
            I => \N__35942\
        );

    \I__7424\ : InMux
    port map (
            O => \N__36002\,
            I => \N__35942\
        );

    \I__7423\ : InMux
    port map (
            O => \N__36001\,
            I => \N__35942\
        );

    \I__7422\ : InMux
    port map (
            O => \N__36000\,
            I => \N__35942\
        );

    \I__7421\ : LocalMux
    port map (
            O => \N__35991\,
            I => \N__35933\
        );

    \I__7420\ : LocalMux
    port map (
            O => \N__35982\,
            I => \N__35933\
        );

    \I__7419\ : Span4Mux_h
    port map (
            O => \N__35979\,
            I => \N__35933\
        );

    \I__7418\ : Span4Mux_v
    port map (
            O => \N__35976\,
            I => \N__35933\
        );

    \I__7417\ : LocalMux
    port map (
            O => \N__35969\,
            I => \N__35930\
        );

    \I__7416\ : Span4Mux_v
    port map (
            O => \N__35966\,
            I => \N__35925\
        );

    \I__7415\ : LocalMux
    port map (
            O => \N__35963\,
            I => \N__35925\
        );

    \I__7414\ : LocalMux
    port map (
            O => \N__35960\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__7413\ : LocalMux
    port map (
            O => \N__35951\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__7412\ : LocalMux
    port map (
            O => \N__35942\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__7411\ : Odrv4
    port map (
            O => \N__35933\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__7410\ : Odrv12
    port map (
            O => \N__35930\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__7409\ : Odrv4
    port map (
            O => \N__35925\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__7408\ : InMux
    port map (
            O => \N__35912\,
            I => \N__35909\
        );

    \I__7407\ : LocalMux
    port map (
            O => \N__35909\,
            I => \N__35906\
        );

    \I__7406\ : Odrv12
    port map (
            O => \N__35906\,
            I => delay_tr_input_c
        );

    \I__7405\ : InMux
    port map (
            O => \N__35903\,
            I => \N__35900\
        );

    \I__7404\ : LocalMux
    port map (
            O => \N__35900\,
            I => delay_tr_d1
        );

    \I__7403\ : CEMux
    port map (
            O => \N__35897\,
            I => \N__35894\
        );

    \I__7402\ : LocalMux
    port map (
            O => \N__35894\,
            I => \N__35891\
        );

    \I__7401\ : Span4Mux_h
    port map (
            O => \N__35891\,
            I => \N__35888\
        );

    \I__7400\ : Span4Mux_v
    port map (
            O => \N__35888\,
            I => \N__35884\
        );

    \I__7399\ : CEMux
    port map (
            O => \N__35887\,
            I => \N__35881\
        );

    \I__7398\ : Span4Mux_v
    port map (
            O => \N__35884\,
            I => \N__35874\
        );

    \I__7397\ : LocalMux
    port map (
            O => \N__35881\,
            I => \N__35874\
        );

    \I__7396\ : IoInMux
    port map (
            O => \N__35880\,
            I => \N__35871\
        );

    \I__7395\ : CEMux
    port map (
            O => \N__35879\,
            I => \N__35868\
        );

    \I__7394\ : Span4Mux_v
    port map (
            O => \N__35874\,
            I => \N__35865\
        );

    \I__7393\ : LocalMux
    port map (
            O => \N__35871\,
            I => \N__35862\
        );

    \I__7392\ : LocalMux
    port map (
            O => \N__35868\,
            I => \N__35858\
        );

    \I__7391\ : Span4Mux_v
    port map (
            O => \N__35865\,
            I => \N__35855\
        );

    \I__7390\ : IoSpan4Mux
    port map (
            O => \N__35862\,
            I => \N__35852\
        );

    \I__7389\ : CEMux
    port map (
            O => \N__35861\,
            I => \N__35849\
        );

    \I__7388\ : Span12Mux_h
    port map (
            O => \N__35858\,
            I => \N__35846\
        );

    \I__7387\ : Span4Mux_v
    port map (
            O => \N__35855\,
            I => \N__35841\
        );

    \I__7386\ : Span4Mux_s0_v
    port map (
            O => \N__35852\,
            I => \N__35841\
        );

    \I__7385\ : LocalMux
    port map (
            O => \N__35849\,
            I => \N__35838\
        );

    \I__7384\ : Span12Mux_v
    port map (
            O => \N__35846\,
            I => \N__35833\
        );

    \I__7383\ : Span4Mux_v
    port map (
            O => \N__35841\,
            I => \N__35828\
        );

    \I__7382\ : Span4Mux_h
    port map (
            O => \N__35838\,
            I => \N__35828\
        );

    \I__7381\ : CEMux
    port map (
            O => \N__35837\,
            I => \N__35825\
        );

    \I__7380\ : CEMux
    port map (
            O => \N__35836\,
            I => \N__35822\
        );

    \I__7379\ : Odrv12
    port map (
            O => \N__35833\,
            I => red_c_i
        );

    \I__7378\ : Odrv4
    port map (
            O => \N__35828\,
            I => red_c_i
        );

    \I__7377\ : LocalMux
    port map (
            O => \N__35825\,
            I => red_c_i
        );

    \I__7376\ : LocalMux
    port map (
            O => \N__35822\,
            I => red_c_i
        );

    \I__7375\ : InMux
    port map (
            O => \N__35813\,
            I => \N__35810\
        );

    \I__7374\ : LocalMux
    port map (
            O => \N__35810\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2\
        );

    \I__7373\ : InMux
    port map (
            O => \N__35807\,
            I => \N__35804\
        );

    \I__7372\ : LocalMux
    port map (
            O => \N__35804\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3\
        );

    \I__7371\ : InMux
    port map (
            O => \N__35801\,
            I => \N__35798\
        );

    \I__7370\ : LocalMux
    port map (
            O => \N__35798\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4\
        );

    \I__7369\ : InMux
    port map (
            O => \N__35795\,
            I => \N__35792\
        );

    \I__7368\ : LocalMux
    port map (
            O => \N__35792\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15\
        );

    \I__7367\ : InMux
    port map (
            O => \N__35789\,
            I => \N__35786\
        );

    \I__7366\ : LocalMux
    port map (
            O => \N__35786\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6\
        );

    \I__7365\ : InMux
    port map (
            O => \N__35783\,
            I => \N__35780\
        );

    \I__7364\ : LocalMux
    port map (
            O => \N__35780\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10\
        );

    \I__7363\ : InMux
    port map (
            O => \N__35777\,
            I => \N__35774\
        );

    \I__7362\ : LocalMux
    port map (
            O => \N__35774\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17\
        );

    \I__7361\ : InMux
    port map (
            O => \N__35771\,
            I => \N__35768\
        );

    \I__7360\ : LocalMux
    port map (
            O => \N__35768\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5\
        );

    \I__7359\ : InMux
    port map (
            O => \N__35765\,
            I => \N__35762\
        );

    \I__7358\ : LocalMux
    port map (
            O => \N__35762\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19\
        );

    \I__7357\ : InMux
    port map (
            O => \N__35759\,
            I => \N__35756\
        );

    \I__7356\ : LocalMux
    port map (
            O => \N__35756\,
            I => \N__35753\
        );

    \I__7355\ : Odrv4
    port map (
            O => \N__35753\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6\
        );

    \I__7354\ : InMux
    port map (
            O => \N__35750\,
            I => \N__35747\
        );

    \I__7353\ : LocalMux
    port map (
            O => \N__35747\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7\
        );

    \I__7352\ : InMux
    port map (
            O => \N__35744\,
            I => \N__35741\
        );

    \I__7351\ : LocalMux
    port map (
            O => \N__35741\,
            I => \N__35738\
        );

    \I__7350\ : Odrv4
    port map (
            O => \N__35738\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9\
        );

    \I__7349\ : InMux
    port map (
            O => \N__35735\,
            I => \N__35732\
        );

    \I__7348\ : LocalMux
    port map (
            O => \N__35732\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8\
        );

    \I__7347\ : InMux
    port map (
            O => \N__35729\,
            I => \N__35726\
        );

    \I__7346\ : LocalMux
    port map (
            O => \N__35726\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12\
        );

    \I__7345\ : InMux
    port map (
            O => \N__35723\,
            I => \N__35720\
        );

    \I__7344\ : LocalMux
    port map (
            O => \N__35720\,
            I => \N__35717\
        );

    \I__7343\ : Span12Mux_s9_v
    port map (
            O => \N__35717\,
            I => \N__35714\
        );

    \I__7342\ : Odrv12
    port map (
            O => \N__35714\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0\
        );

    \I__7341\ : InMux
    port map (
            O => \N__35711\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16\
        );

    \I__7340\ : InMux
    port map (
            O => \N__35708\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17\
        );

    \I__7339\ : InMux
    port map (
            O => \N__35705\,
            I => \N__35702\
        );

    \I__7338\ : LocalMux
    port map (
            O => \N__35702\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17\
        );

    \I__7337\ : InMux
    port map (
            O => \N__35699\,
            I => \N__35696\
        );

    \I__7336\ : LocalMux
    port map (
            O => \N__35696\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18\
        );

    \I__7335\ : InMux
    port map (
            O => \N__35693\,
            I => \N__35690\
        );

    \I__7334\ : LocalMux
    port map (
            O => \N__35690\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19\
        );

    \I__7333\ : InMux
    port map (
            O => \N__35687\,
            I => \N__35684\
        );

    \I__7332\ : LocalMux
    port map (
            O => \N__35684\,
            I => \N__35681\
        );

    \I__7331\ : Odrv12
    port map (
            O => \N__35681\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2\
        );

    \I__7330\ : InMux
    port map (
            O => \N__35678\,
            I => \N__35675\
        );

    \I__7329\ : LocalMux
    port map (
            O => \N__35675\,
            I => \N__35672\
        );

    \I__7328\ : Odrv4
    port map (
            O => \N__35672\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3\
        );

    \I__7327\ : InMux
    port map (
            O => \N__35669\,
            I => \N__35666\
        );

    \I__7326\ : LocalMux
    port map (
            O => \N__35666\,
            I => \N__35663\
        );

    \I__7325\ : Odrv4
    port map (
            O => \N__35663\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4\
        );

    \I__7324\ : InMux
    port map (
            O => \N__35660\,
            I => \N__35657\
        );

    \I__7323\ : LocalMux
    port map (
            O => \N__35657\,
            I => \N__35654\
        );

    \I__7322\ : Odrv4
    port map (
            O => \N__35654\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5\
        );

    \I__7321\ : InMux
    port map (
            O => \N__35651\,
            I => \bfn_14_19_0_\
        );

    \I__7320\ : InMux
    port map (
            O => \N__35648\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8\
        );

    \I__7319\ : InMux
    port map (
            O => \N__35645\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9\
        );

    \I__7318\ : InMux
    port map (
            O => \N__35642\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10\
        );

    \I__7317\ : InMux
    port map (
            O => \N__35639\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11\
        );

    \I__7316\ : InMux
    port map (
            O => \N__35636\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12\
        );

    \I__7315\ : InMux
    port map (
            O => \N__35633\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13\
        );

    \I__7314\ : InMux
    port map (
            O => \N__35630\,
            I => \N__35627\
        );

    \I__7313\ : LocalMux
    port map (
            O => \N__35627\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16\
        );

    \I__7312\ : InMux
    port map (
            O => \N__35624\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14\
        );

    \I__7311\ : InMux
    port map (
            O => \N__35621\,
            I => \bfn_14_20_0_\
        );

    \I__7310\ : CascadeMux
    port map (
            O => \N__35618\,
            I => \N__35612\
        );

    \I__7309\ : InMux
    port map (
            O => \N__35617\,
            I => \N__35605\
        );

    \I__7308\ : InMux
    port map (
            O => \N__35616\,
            I => \N__35605\
        );

    \I__7307\ : CascadeMux
    port map (
            O => \N__35615\,
            I => \N__35601\
        );

    \I__7306\ : InMux
    port map (
            O => \N__35612\,
            I => \N__35587\
        );

    \I__7305\ : InMux
    port map (
            O => \N__35611\,
            I => \N__35587\
        );

    \I__7304\ : InMux
    port map (
            O => \N__35610\,
            I => \N__35587\
        );

    \I__7303\ : LocalMux
    port map (
            O => \N__35605\,
            I => \N__35580\
        );

    \I__7302\ : InMux
    port map (
            O => \N__35604\,
            I => \N__35577\
        );

    \I__7301\ : InMux
    port map (
            O => \N__35601\,
            I => \N__35568\
        );

    \I__7300\ : InMux
    port map (
            O => \N__35600\,
            I => \N__35568\
        );

    \I__7299\ : InMux
    port map (
            O => \N__35599\,
            I => \N__35568\
        );

    \I__7298\ : InMux
    port map (
            O => \N__35598\,
            I => \N__35568\
        );

    \I__7297\ : InMux
    port map (
            O => \N__35597\,
            I => \N__35559\
        );

    \I__7296\ : InMux
    port map (
            O => \N__35596\,
            I => \N__35559\
        );

    \I__7295\ : InMux
    port map (
            O => \N__35595\,
            I => \N__35559\
        );

    \I__7294\ : InMux
    port map (
            O => \N__35594\,
            I => \N__35559\
        );

    \I__7293\ : LocalMux
    port map (
            O => \N__35587\,
            I => \N__35556\
        );

    \I__7292\ : InMux
    port map (
            O => \N__35586\,
            I => \N__35547\
        );

    \I__7291\ : InMux
    port map (
            O => \N__35585\,
            I => \N__35547\
        );

    \I__7290\ : InMux
    port map (
            O => \N__35584\,
            I => \N__35547\
        );

    \I__7289\ : InMux
    port map (
            O => \N__35583\,
            I => \N__35547\
        );

    \I__7288\ : Span4Mux_h
    port map (
            O => \N__35580\,
            I => \N__35544\
        );

    \I__7287\ : LocalMux
    port map (
            O => \N__35577\,
            I => \N__35537\
        );

    \I__7286\ : LocalMux
    port map (
            O => \N__35568\,
            I => \N__35528\
        );

    \I__7285\ : LocalMux
    port map (
            O => \N__35559\,
            I => \N__35528\
        );

    \I__7284\ : Span4Mux_v
    port map (
            O => \N__35556\,
            I => \N__35528\
        );

    \I__7283\ : LocalMux
    port map (
            O => \N__35547\,
            I => \N__35528\
        );

    \I__7282\ : Span4Mux_h
    port map (
            O => \N__35544\,
            I => \N__35525\
        );

    \I__7281\ : InMux
    port map (
            O => \N__35543\,
            I => \N__35516\
        );

    \I__7280\ : InMux
    port map (
            O => \N__35542\,
            I => \N__35516\
        );

    \I__7279\ : InMux
    port map (
            O => \N__35541\,
            I => \N__35516\
        );

    \I__7278\ : InMux
    port map (
            O => \N__35540\,
            I => \N__35516\
        );

    \I__7277\ : Span4Mux_h
    port map (
            O => \N__35537\,
            I => \N__35513\
        );

    \I__7276\ : Span4Mux_v
    port map (
            O => \N__35528\,
            I => \N__35508\
        );

    \I__7275\ : Span4Mux_h
    port map (
            O => \N__35525\,
            I => \N__35508\
        );

    \I__7274\ : LocalMux
    port map (
            O => \N__35516\,
            I => \phase_controller_inst1.stoper_hc.un2_startlt31\
        );

    \I__7273\ : Odrv4
    port map (
            O => \N__35513\,
            I => \phase_controller_inst1.stoper_hc.un2_startlt31\
        );

    \I__7272\ : Odrv4
    port map (
            O => \N__35508\,
            I => \phase_controller_inst1.stoper_hc.un2_startlt31\
        );

    \I__7271\ : InMux
    port map (
            O => \N__35501\,
            I => \N__35496\
        );

    \I__7270\ : CascadeMux
    port map (
            O => \N__35500\,
            I => \N__35493\
        );

    \I__7269\ : InMux
    port map (
            O => \N__35499\,
            I => \N__35490\
        );

    \I__7268\ : LocalMux
    port map (
            O => \N__35496\,
            I => \N__35485\
        );

    \I__7267\ : InMux
    port map (
            O => \N__35493\,
            I => \N__35482\
        );

    \I__7266\ : LocalMux
    port map (
            O => \N__35490\,
            I => \N__35479\
        );

    \I__7265\ : InMux
    port map (
            O => \N__35489\,
            I => \N__35476\
        );

    \I__7264\ : InMux
    port map (
            O => \N__35488\,
            I => \N__35473\
        );

    \I__7263\ : Span4Mux_v
    port map (
            O => \N__35485\,
            I => \N__35470\
        );

    \I__7262\ : LocalMux
    port map (
            O => \N__35482\,
            I => \N__35467\
        );

    \I__7261\ : Span4Mux_v
    port map (
            O => \N__35479\,
            I => \N__35462\
        );

    \I__7260\ : LocalMux
    port map (
            O => \N__35476\,
            I => \N__35462\
        );

    \I__7259\ : LocalMux
    port map (
            O => \N__35473\,
            I => measured_delay_hc_8
        );

    \I__7258\ : Odrv4
    port map (
            O => \N__35470\,
            I => measured_delay_hc_8
        );

    \I__7257\ : Odrv12
    port map (
            O => \N__35467\,
            I => measured_delay_hc_8
        );

    \I__7256\ : Odrv4
    port map (
            O => \N__35462\,
            I => measured_delay_hc_8
        );

    \I__7255\ : InMux
    port map (
            O => \N__35453\,
            I => \N__35440\
        );

    \I__7254\ : InMux
    port map (
            O => \N__35452\,
            I => \N__35440\
        );

    \I__7253\ : InMux
    port map (
            O => \N__35451\,
            I => \N__35440\
        );

    \I__7252\ : InMux
    port map (
            O => \N__35450\,
            I => \N__35427\
        );

    \I__7251\ : InMux
    port map (
            O => \N__35449\,
            I => \N__35427\
        );

    \I__7250\ : InMux
    port map (
            O => \N__35448\,
            I => \N__35427\
        );

    \I__7249\ : InMux
    port map (
            O => \N__35447\,
            I => \N__35427\
        );

    \I__7248\ : LocalMux
    port map (
            O => \N__35440\,
            I => \N__35424\
        );

    \I__7247\ : InMux
    port map (
            O => \N__35439\,
            I => \N__35415\
        );

    \I__7246\ : InMux
    port map (
            O => \N__35438\,
            I => \N__35415\
        );

    \I__7245\ : InMux
    port map (
            O => \N__35437\,
            I => \N__35415\
        );

    \I__7244\ : InMux
    port map (
            O => \N__35436\,
            I => \N__35415\
        );

    \I__7243\ : LocalMux
    port map (
            O => \N__35427\,
            I => \N__35409\
        );

    \I__7242\ : Span4Mux_v
    port map (
            O => \N__35424\,
            I => \N__35404\
        );

    \I__7241\ : LocalMux
    port map (
            O => \N__35415\,
            I => \N__35404\
        );

    \I__7240\ : InMux
    port map (
            O => \N__35414\,
            I => \N__35397\
        );

    \I__7239\ : InMux
    port map (
            O => \N__35413\,
            I => \N__35397\
        );

    \I__7238\ : InMux
    port map (
            O => \N__35412\,
            I => \N__35397\
        );

    \I__7237\ : Odrv12
    port map (
            O => \N__35409\,
            I => \phase_controller_inst1.stoper_hc.un1_start\
        );

    \I__7236\ : Odrv4
    port map (
            O => \N__35404\,
            I => \phase_controller_inst1.stoper_hc.un1_start\
        );

    \I__7235\ : LocalMux
    port map (
            O => \N__35397\,
            I => \phase_controller_inst1.stoper_hc.un1_start\
        );

    \I__7234\ : InMux
    port map (
            O => \N__35390\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0\
        );

    \I__7233\ : InMux
    port map (
            O => \N__35387\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1\
        );

    \I__7232\ : InMux
    port map (
            O => \N__35384\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2\
        );

    \I__7231\ : InMux
    port map (
            O => \N__35381\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3\
        );

    \I__7230\ : InMux
    port map (
            O => \N__35378\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4\
        );

    \I__7229\ : InMux
    port map (
            O => \N__35375\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5\
        );

    \I__7228\ : InMux
    port map (
            O => \N__35372\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6\
        );

    \I__7227\ : InMux
    port map (
            O => \N__35369\,
            I => \N__35365\
        );

    \I__7226\ : CascadeMux
    port map (
            O => \N__35368\,
            I => \N__35361\
        );

    \I__7225\ : LocalMux
    port map (
            O => \N__35365\,
            I => \N__35357\
        );

    \I__7224\ : InMux
    port map (
            O => \N__35364\,
            I => \N__35354\
        );

    \I__7223\ : InMux
    port map (
            O => \N__35361\,
            I => \N__35351\
        );

    \I__7222\ : CascadeMux
    port map (
            O => \N__35360\,
            I => \N__35347\
        );

    \I__7221\ : Sp12to4
    port map (
            O => \N__35357\,
            I => \N__35342\
        );

    \I__7220\ : LocalMux
    port map (
            O => \N__35354\,
            I => \N__35342\
        );

    \I__7219\ : LocalMux
    port map (
            O => \N__35351\,
            I => \N__35339\
        );

    \I__7218\ : CascadeMux
    port map (
            O => \N__35350\,
            I => \N__35336\
        );

    \I__7217\ : InMux
    port map (
            O => \N__35347\,
            I => \N__35333\
        );

    \I__7216\ : Span12Mux_v
    port map (
            O => \N__35342\,
            I => \N__35330\
        );

    \I__7215\ : Span4Mux_h
    port map (
            O => \N__35339\,
            I => \N__35327\
        );

    \I__7214\ : InMux
    port map (
            O => \N__35336\,
            I => \N__35324\
        );

    \I__7213\ : LocalMux
    port map (
            O => \N__35333\,
            I => measured_delay_hc_12
        );

    \I__7212\ : Odrv12
    port map (
            O => \N__35330\,
            I => measured_delay_hc_12
        );

    \I__7211\ : Odrv4
    port map (
            O => \N__35327\,
            I => measured_delay_hc_12
        );

    \I__7210\ : LocalMux
    port map (
            O => \N__35324\,
            I => measured_delay_hc_12
        );

    \I__7209\ : InMux
    port map (
            O => \N__35315\,
            I => \N__35312\
        );

    \I__7208\ : LocalMux
    port map (
            O => \N__35312\,
            I => \N__35308\
        );

    \I__7207\ : InMux
    port map (
            O => \N__35311\,
            I => \N__35305\
        );

    \I__7206\ : Span4Mux_v
    port map (
            O => \N__35308\,
            I => \N__35298\
        );

    \I__7205\ : LocalMux
    port map (
            O => \N__35305\,
            I => \N__35298\
        );

    \I__7204\ : InMux
    port map (
            O => \N__35304\,
            I => \N__35295\
        );

    \I__7203\ : InMux
    port map (
            O => \N__35303\,
            I => \N__35292\
        );

    \I__7202\ : Span4Mux_h
    port map (
            O => \N__35298\,
            I => \N__35289\
        );

    \I__7201\ : LocalMux
    port map (
            O => \N__35295\,
            I => \N__35286\
        );

    \I__7200\ : LocalMux
    port map (
            O => \N__35292\,
            I => measured_delay_hc_1
        );

    \I__7199\ : Odrv4
    port map (
            O => \N__35289\,
            I => measured_delay_hc_1
        );

    \I__7198\ : Odrv12
    port map (
            O => \N__35286\,
            I => measured_delay_hc_1
        );

    \I__7197\ : CascadeMux
    port map (
            O => \N__35279\,
            I => \N__35275\
        );

    \I__7196\ : CascadeMux
    port map (
            O => \N__35278\,
            I => \N__35271\
        );

    \I__7195\ : InMux
    port map (
            O => \N__35275\,
            I => \N__35268\
        );

    \I__7194\ : CascadeMux
    port map (
            O => \N__35274\,
            I => \N__35264\
        );

    \I__7193\ : InMux
    port map (
            O => \N__35271\,
            I => \N__35261\
        );

    \I__7192\ : LocalMux
    port map (
            O => \N__35268\,
            I => \N__35258\
        );

    \I__7191\ : InMux
    port map (
            O => \N__35267\,
            I => \N__35253\
        );

    \I__7190\ : InMux
    port map (
            O => \N__35264\,
            I => \N__35253\
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__35261\,
            I => \N__35249\
        );

    \I__7188\ : Span4Mux_v
    port map (
            O => \N__35258\,
            I => \N__35244\
        );

    \I__7187\ : LocalMux
    port map (
            O => \N__35253\,
            I => \N__35244\
        );

    \I__7186\ : InMux
    port map (
            O => \N__35252\,
            I => \N__35241\
        );

    \I__7185\ : Span12Mux_h
    port map (
            O => \N__35249\,
            I => \N__35238\
        );

    \I__7184\ : Span4Mux_v
    port map (
            O => \N__35244\,
            I => \N__35235\
        );

    \I__7183\ : LocalMux
    port map (
            O => \N__35241\,
            I => measured_delay_hc_3
        );

    \I__7182\ : Odrv12
    port map (
            O => \N__35238\,
            I => measured_delay_hc_3
        );

    \I__7181\ : Odrv4
    port map (
            O => \N__35235\,
            I => measured_delay_hc_3
        );

    \I__7180\ : InMux
    port map (
            O => \N__35228\,
            I => \N__35225\
        );

    \I__7179\ : LocalMux
    port map (
            O => \N__35225\,
            I => \N__35222\
        );

    \I__7178\ : Span4Mux_h
    port map (
            O => \N__35222\,
            I => \N__35218\
        );

    \I__7177\ : InMux
    port map (
            O => \N__35221\,
            I => \N__35215\
        );

    \I__7176\ : Span4Mux_v
    port map (
            O => \N__35218\,
            I => \N__35210\
        );

    \I__7175\ : LocalMux
    port map (
            O => \N__35215\,
            I => \N__35207\
        );

    \I__7174\ : InMux
    port map (
            O => \N__35214\,
            I => \N__35202\
        );

    \I__7173\ : InMux
    port map (
            O => \N__35213\,
            I => \N__35202\
        );

    \I__7172\ : Odrv4
    port map (
            O => \N__35210\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_2\
        );

    \I__7171\ : Odrv12
    port map (
            O => \N__35207\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_2\
        );

    \I__7170\ : LocalMux
    port map (
            O => \N__35202\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_2\
        );

    \I__7169\ : InMux
    port map (
            O => \N__35195\,
            I => \N__35191\
        );

    \I__7168\ : CascadeMux
    port map (
            O => \N__35194\,
            I => \N__35188\
        );

    \I__7167\ : LocalMux
    port map (
            O => \N__35191\,
            I => \N__35184\
        );

    \I__7166\ : InMux
    port map (
            O => \N__35188\,
            I => \N__35181\
        );

    \I__7165\ : InMux
    port map (
            O => \N__35187\,
            I => \N__35177\
        );

    \I__7164\ : Span4Mux_v
    port map (
            O => \N__35184\,
            I => \N__35173\
        );

    \I__7163\ : LocalMux
    port map (
            O => \N__35181\,
            I => \N__35170\
        );

    \I__7162\ : InMux
    port map (
            O => \N__35180\,
            I => \N__35167\
        );

    \I__7161\ : LocalMux
    port map (
            O => \N__35177\,
            I => \N__35164\
        );

    \I__7160\ : InMux
    port map (
            O => \N__35176\,
            I => \N__35161\
        );

    \I__7159\ : Span4Mux_v
    port map (
            O => \N__35173\,
            I => \N__35158\
        );

    \I__7158\ : Span4Mux_v
    port map (
            O => \N__35170\,
            I => \N__35151\
        );

    \I__7157\ : LocalMux
    port map (
            O => \N__35167\,
            I => \N__35151\
        );

    \I__7156\ : Span4Mux_h
    port map (
            O => \N__35164\,
            I => \N__35151\
        );

    \I__7155\ : LocalMux
    port map (
            O => \N__35161\,
            I => measured_delay_hc_15
        );

    \I__7154\ : Odrv4
    port map (
            O => \N__35158\,
            I => measured_delay_hc_15
        );

    \I__7153\ : Odrv4
    port map (
            O => \N__35151\,
            I => measured_delay_hc_15
        );

    \I__7152\ : InMux
    port map (
            O => \N__35144\,
            I => \N__35140\
        );

    \I__7151\ : InMux
    port map (
            O => \N__35143\,
            I => \N__35137\
        );

    \I__7150\ : LocalMux
    port map (
            O => \N__35140\,
            I => \N__35133\
        );

    \I__7149\ : LocalMux
    port map (
            O => \N__35137\,
            I => \N__35128\
        );

    \I__7148\ : InMux
    port map (
            O => \N__35136\,
            I => \N__35125\
        );

    \I__7147\ : Span4Mux_v
    port map (
            O => \N__35133\,
            I => \N__35122\
        );

    \I__7146\ : InMux
    port map (
            O => \N__35132\,
            I => \N__35119\
        );

    \I__7145\ : InMux
    port map (
            O => \N__35131\,
            I => \N__35116\
        );

    \I__7144\ : Span12Mux_v
    port map (
            O => \N__35128\,
            I => \N__35113\
        );

    \I__7143\ : LocalMux
    port map (
            O => \N__35125\,
            I => \N__35110\
        );

    \I__7142\ : Span4Mux_v
    port map (
            O => \N__35122\,
            I => \N__35105\
        );

    \I__7141\ : LocalMux
    port map (
            O => \N__35119\,
            I => \N__35105\
        );

    \I__7140\ : LocalMux
    port map (
            O => \N__35116\,
            I => measured_delay_hc_13
        );

    \I__7139\ : Odrv12
    port map (
            O => \N__35113\,
            I => measured_delay_hc_13
        );

    \I__7138\ : Odrv12
    port map (
            O => \N__35110\,
            I => measured_delay_hc_13
        );

    \I__7137\ : Odrv4
    port map (
            O => \N__35105\,
            I => measured_delay_hc_13
        );

    \I__7136\ : InMux
    port map (
            O => \N__35096\,
            I => \N__35092\
        );

    \I__7135\ : CascadeMux
    port map (
            O => \N__35095\,
            I => \N__35086\
        );

    \I__7134\ : LocalMux
    port map (
            O => \N__35092\,
            I => \N__35083\
        );

    \I__7133\ : InMux
    port map (
            O => \N__35091\,
            I => \N__35080\
        );

    \I__7132\ : InMux
    port map (
            O => \N__35090\,
            I => \N__35075\
        );

    \I__7131\ : InMux
    port map (
            O => \N__35089\,
            I => \N__35075\
        );

    \I__7130\ : InMux
    port map (
            O => \N__35086\,
            I => \N__35072\
        );

    \I__7129\ : Sp12to4
    port map (
            O => \N__35083\,
            I => \N__35067\
        );

    \I__7128\ : LocalMux
    port map (
            O => \N__35080\,
            I => \N__35067\
        );

    \I__7127\ : LocalMux
    port map (
            O => \N__35075\,
            I => \N__35064\
        );

    \I__7126\ : LocalMux
    port map (
            O => \N__35072\,
            I => measured_delay_hc_18
        );

    \I__7125\ : Odrv12
    port map (
            O => \N__35067\,
            I => measured_delay_hc_18
        );

    \I__7124\ : Odrv4
    port map (
            O => \N__35064\,
            I => measured_delay_hc_18
        );

    \I__7123\ : InMux
    port map (
            O => \N__35057\,
            I => \N__35053\
        );

    \I__7122\ : InMux
    port map (
            O => \N__35056\,
            I => \N__35050\
        );

    \I__7121\ : LocalMux
    port map (
            O => \N__35053\,
            I => \N__35047\
        );

    \I__7120\ : LocalMux
    port map (
            O => \N__35050\,
            I => \N__35040\
        );

    \I__7119\ : Span4Mux_h
    port map (
            O => \N__35047\,
            I => \N__35040\
        );

    \I__7118\ : InMux
    port map (
            O => \N__35046\,
            I => \N__35036\
        );

    \I__7117\ : InMux
    port map (
            O => \N__35045\,
            I => \N__35033\
        );

    \I__7116\ : Span4Mux_v
    port map (
            O => \N__35040\,
            I => \N__35030\
        );

    \I__7115\ : InMux
    port map (
            O => \N__35039\,
            I => \N__35027\
        );

    \I__7114\ : LocalMux
    port map (
            O => \N__35036\,
            I => \N__35024\
        );

    \I__7113\ : LocalMux
    port map (
            O => \N__35033\,
            I => measured_delay_hc_6
        );

    \I__7112\ : Odrv4
    port map (
            O => \N__35030\,
            I => measured_delay_hc_6
        );

    \I__7111\ : LocalMux
    port map (
            O => \N__35027\,
            I => measured_delay_hc_6
        );

    \I__7110\ : Odrv4
    port map (
            O => \N__35024\,
            I => measured_delay_hc_6
        );

    \I__7109\ : InMux
    port map (
            O => \N__35015\,
            I => \N__35002\
        );

    \I__7108\ : InMux
    port map (
            O => \N__35014\,
            I => \N__35002\
        );

    \I__7107\ : InMux
    port map (
            O => \N__35013\,
            I => \N__35002\
        );

    \I__7106\ : InMux
    port map (
            O => \N__35012\,
            I => \N__34993\
        );

    \I__7105\ : InMux
    port map (
            O => \N__35011\,
            I => \N__34993\
        );

    \I__7104\ : InMux
    port map (
            O => \N__35010\,
            I => \N__34993\
        );

    \I__7103\ : InMux
    port map (
            O => \N__35009\,
            I => \N__34993\
        );

    \I__7102\ : LocalMux
    port map (
            O => \N__35002\,
            I => \N__34982\
        );

    \I__7101\ : LocalMux
    port map (
            O => \N__34993\,
            I => \N__34979\
        );

    \I__7100\ : InMux
    port map (
            O => \N__34992\,
            I => \N__34976\
        );

    \I__7099\ : InMux
    port map (
            O => \N__34991\,
            I => \N__34969\
        );

    \I__7098\ : InMux
    port map (
            O => \N__34990\,
            I => \N__34969\
        );

    \I__7097\ : InMux
    port map (
            O => \N__34989\,
            I => \N__34969\
        );

    \I__7096\ : InMux
    port map (
            O => \N__34988\,
            I => \N__34964\
        );

    \I__7095\ : InMux
    port map (
            O => \N__34987\,
            I => \N__34964\
        );

    \I__7094\ : InMux
    port map (
            O => \N__34986\,
            I => \N__34958\
        );

    \I__7093\ : InMux
    port map (
            O => \N__34985\,
            I => \N__34958\
        );

    \I__7092\ : Span4Mux_h
    port map (
            O => \N__34982\,
            I => \N__34955\
        );

    \I__7091\ : Span4Mux_h
    port map (
            O => \N__34979\,
            I => \N__34950\
        );

    \I__7090\ : LocalMux
    port map (
            O => \N__34976\,
            I => \N__34950\
        );

    \I__7089\ : LocalMux
    port map (
            O => \N__34969\,
            I => \N__34945\
        );

    \I__7088\ : LocalMux
    port map (
            O => \N__34964\,
            I => \N__34942\
        );

    \I__7087\ : InMux
    port map (
            O => \N__34963\,
            I => \N__34939\
        );

    \I__7086\ : LocalMux
    port map (
            O => \N__34958\,
            I => \N__34936\
        );

    \I__7085\ : Span4Mux_v
    port map (
            O => \N__34955\,
            I => \N__34933\
        );

    \I__7084\ : Span4Mux_v
    port map (
            O => \N__34950\,
            I => \N__34930\
        );

    \I__7083\ : InMux
    port map (
            O => \N__34949\,
            I => \N__34925\
        );

    \I__7082\ : InMux
    port map (
            O => \N__34948\,
            I => \N__34925\
        );

    \I__7081\ : Span12Mux_s11_v
    port map (
            O => \N__34945\,
            I => \N__34922\
        );

    \I__7080\ : Span4Mux_v
    port map (
            O => \N__34942\,
            I => \N__34915\
        );

    \I__7079\ : LocalMux
    port map (
            O => \N__34939\,
            I => \N__34915\
        );

    \I__7078\ : Span4Mux_h
    port map (
            O => \N__34936\,
            I => \N__34915\
        );

    \I__7077\ : Odrv4
    port map (
            O => \N__34933\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt31_0\
        );

    \I__7076\ : Odrv4
    port map (
            O => \N__34930\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt31_0\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__34925\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt31_0\
        );

    \I__7074\ : Odrv12
    port map (
            O => \N__34922\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt31_0\
        );

    \I__7073\ : Odrv4
    port map (
            O => \N__34915\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt31_0\
        );

    \I__7072\ : InMux
    port map (
            O => \N__34904\,
            I => \N__34900\
        );

    \I__7071\ : InMux
    port map (
            O => \N__34903\,
            I => \N__34897\
        );

    \I__7070\ : LocalMux
    port map (
            O => \N__34900\,
            I => \N__34894\
        );

    \I__7069\ : LocalMux
    port map (
            O => \N__34897\,
            I => \N__34888\
        );

    \I__7068\ : Span4Mux_h
    port map (
            O => \N__34894\,
            I => \N__34888\
        );

    \I__7067\ : InMux
    port map (
            O => \N__34893\,
            I => \N__34885\
        );

    \I__7066\ : Span4Mux_v
    port map (
            O => \N__34888\,
            I => \N__34880\
        );

    \I__7065\ : LocalMux
    port map (
            O => \N__34885\,
            I => \N__34880\
        );

    \I__7064\ : Odrv4
    port map (
            O => \N__34880\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2\
        );

    \I__7063\ : InMux
    port map (
            O => \N__34877\,
            I => \N__34874\
        );

    \I__7062\ : LocalMux
    port map (
            O => \N__34874\,
            I => \N__34870\
        );

    \I__7061\ : InMux
    port map (
            O => \N__34873\,
            I => \N__34867\
        );

    \I__7060\ : Span4Mux_h
    port map (
            O => \N__34870\,
            I => \N__34864\
        );

    \I__7059\ : LocalMux
    port map (
            O => \N__34867\,
            I => \N__34861\
        );

    \I__7058\ : Odrv4
    port map (
            O => \N__34864\,
            I => \phase_controller_inst1.stoper_hc.un1_N_4\
        );

    \I__7057\ : Odrv12
    port map (
            O => \N__34861\,
            I => \phase_controller_inst1.stoper_hc.un1_N_4\
        );

    \I__7056\ : InMux
    port map (
            O => \N__34856\,
            I => \N__34853\
        );

    \I__7055\ : LocalMux
    port map (
            O => \N__34853\,
            I => \N__34850\
        );

    \I__7054\ : Span4Mux_h
    port map (
            O => \N__34850\,
            I => \N__34847\
        );

    \I__7053\ : Odrv4
    port map (
            O => \N__34847\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto31_dZ0Z_0\
        );

    \I__7052\ : InMux
    port map (
            O => \N__34844\,
            I => \N__34840\
        );

    \I__7051\ : InMux
    port map (
            O => \N__34843\,
            I => \N__34837\
        );

    \I__7050\ : LocalMux
    port map (
            O => \N__34840\,
            I => \N__34834\
        );

    \I__7049\ : LocalMux
    port map (
            O => \N__34837\,
            I => \N__34831\
        );

    \I__7048\ : Span4Mux_h
    port map (
            O => \N__34834\,
            I => \N__34828\
        );

    \I__7047\ : Odrv4
    port map (
            O => \N__34831\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__7046\ : Odrv4
    port map (
            O => \N__34828\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__7045\ : CascadeMux
    port map (
            O => \N__34823\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto31_dZ0Z_0_cascade_\
        );

    \I__7044\ : CascadeMux
    port map (
            O => \N__34820\,
            I => \N__34817\
        );

    \I__7043\ : InMux
    port map (
            O => \N__34817\,
            I => \N__34813\
        );

    \I__7042\ : InMux
    port map (
            O => \N__34816\,
            I => \N__34810\
        );

    \I__7041\ : LocalMux
    port map (
            O => \N__34813\,
            I => \N__34804\
        );

    \I__7040\ : LocalMux
    port map (
            O => \N__34810\,
            I => \N__34801\
        );

    \I__7039\ : InMux
    port map (
            O => \N__34809\,
            I => \N__34796\
        );

    \I__7038\ : InMux
    port map (
            O => \N__34808\,
            I => \N__34796\
        );

    \I__7037\ : CascadeMux
    port map (
            O => \N__34807\,
            I => \N__34793\
        );

    \I__7036\ : Span4Mux_h
    port map (
            O => \N__34804\,
            I => \N__34786\
        );

    \I__7035\ : Span4Mux_h
    port map (
            O => \N__34801\,
            I => \N__34786\
        );

    \I__7034\ : LocalMux
    port map (
            O => \N__34796\,
            I => \N__34786\
        );

    \I__7033\ : InMux
    port map (
            O => \N__34793\,
            I => \N__34783\
        );

    \I__7032\ : Span4Mux_v
    port map (
            O => \N__34786\,
            I => \N__34780\
        );

    \I__7031\ : LocalMux
    port map (
            O => \N__34783\,
            I => measured_delay_hc_16
        );

    \I__7030\ : Odrv4
    port map (
            O => \N__34780\,
            I => measured_delay_hc_16
        );

    \I__7029\ : InMux
    port map (
            O => \N__34775\,
            I => \N__34772\
        );

    \I__7028\ : LocalMux
    port map (
            O => \N__34772\,
            I => \N__34765\
        );

    \I__7027\ : InMux
    port map (
            O => \N__34771\,
            I => \N__34758\
        );

    \I__7026\ : InMux
    port map (
            O => \N__34770\,
            I => \N__34758\
        );

    \I__7025\ : InMux
    port map (
            O => \N__34769\,
            I => \N__34758\
        );

    \I__7024\ : InMux
    port map (
            O => \N__34768\,
            I => \N__34755\
        );

    \I__7023\ : Span4Mux_h
    port map (
            O => \N__34765\,
            I => \N__34752\
        );

    \I__7022\ : LocalMux
    port map (
            O => \N__34758\,
            I => \N__34749\
        );

    \I__7021\ : LocalMux
    port map (
            O => \N__34755\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto31_cZ0Z_0\
        );

    \I__7020\ : Odrv4
    port map (
            O => \N__34752\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto31_cZ0Z_0\
        );

    \I__7019\ : Odrv4
    port map (
            O => \N__34749\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto31_cZ0Z_0\
        );

    \I__7018\ : CascadeMux
    port map (
            O => \N__34742\,
            I => \N__34738\
        );

    \I__7017\ : CascadeMux
    port map (
            O => \N__34741\,
            I => \N__34733\
        );

    \I__7016\ : InMux
    port map (
            O => \N__34738\,
            I => \N__34729\
        );

    \I__7015\ : InMux
    port map (
            O => \N__34737\,
            I => \N__34726\
        );

    \I__7014\ : InMux
    port map (
            O => \N__34736\,
            I => \N__34721\
        );

    \I__7013\ : InMux
    port map (
            O => \N__34733\,
            I => \N__34721\
        );

    \I__7012\ : CascadeMux
    port map (
            O => \N__34732\,
            I => \N__34718\
        );

    \I__7011\ : LocalMux
    port map (
            O => \N__34729\,
            I => \N__34715\
        );

    \I__7010\ : LocalMux
    port map (
            O => \N__34726\,
            I => \N__34712\
        );

    \I__7009\ : LocalMux
    port map (
            O => \N__34721\,
            I => \N__34709\
        );

    \I__7008\ : InMux
    port map (
            O => \N__34718\,
            I => \N__34706\
        );

    \I__7007\ : Span12Mux_v
    port map (
            O => \N__34715\,
            I => \N__34703\
        );

    \I__7006\ : Span4Mux_v
    port map (
            O => \N__34712\,
            I => \N__34698\
        );

    \I__7005\ : Span4Mux_h
    port map (
            O => \N__34709\,
            I => \N__34698\
        );

    \I__7004\ : LocalMux
    port map (
            O => \N__34706\,
            I => measured_delay_hc_17
        );

    \I__7003\ : Odrv12
    port map (
            O => \N__34703\,
            I => measured_delay_hc_17
        );

    \I__7002\ : Odrv4
    port map (
            O => \N__34698\,
            I => measured_delay_hc_17
        );

    \I__7001\ : CascadeMux
    port map (
            O => \N__34691\,
            I => \N__34688\
        );

    \I__7000\ : InMux
    port map (
            O => \N__34688\,
            I => \N__34685\
        );

    \I__6999\ : LocalMux
    port map (
            O => \N__34685\,
            I => \N__34682\
        );

    \I__6998\ : Span12Mux_s8_v
    port map (
            O => \N__34682\,
            I => \N__34677\
        );

    \I__6997\ : InMux
    port map (
            O => \N__34681\,
            I => \N__34674\
        );

    \I__6996\ : InMux
    port map (
            O => \N__34680\,
            I => \N__34669\
        );

    \I__6995\ : Span12Mux_h
    port map (
            O => \N__34677\,
            I => \N__34664\
        );

    \I__6994\ : LocalMux
    port map (
            O => \N__34674\,
            I => \N__34664\
        );

    \I__6993\ : InMux
    port map (
            O => \N__34673\,
            I => \N__34661\
        );

    \I__6992\ : InMux
    port map (
            O => \N__34672\,
            I => \N__34658\
        );

    \I__6991\ : LocalMux
    port map (
            O => \N__34669\,
            I => measured_delay_hc_10
        );

    \I__6990\ : Odrv12
    port map (
            O => \N__34664\,
            I => measured_delay_hc_10
        );

    \I__6989\ : LocalMux
    port map (
            O => \N__34661\,
            I => measured_delay_hc_10
        );

    \I__6988\ : LocalMux
    port map (
            O => \N__34658\,
            I => measured_delay_hc_10
        );

    \I__6987\ : InMux
    port map (
            O => \N__34649\,
            I => \N__34645\
        );

    \I__6986\ : InMux
    port map (
            O => \N__34648\,
            I => \N__34642\
        );

    \I__6985\ : LocalMux
    port map (
            O => \N__34645\,
            I => \N__34637\
        );

    \I__6984\ : LocalMux
    port map (
            O => \N__34642\,
            I => \N__34633\
        );

    \I__6983\ : InMux
    port map (
            O => \N__34641\,
            I => \N__34630\
        );

    \I__6982\ : InMux
    port map (
            O => \N__34640\,
            I => \N__34627\
        );

    \I__6981\ : Span4Mux_v
    port map (
            O => \N__34637\,
            I => \N__34624\
        );

    \I__6980\ : InMux
    port map (
            O => \N__34636\,
            I => \N__34621\
        );

    \I__6979\ : Span4Mux_v
    port map (
            O => \N__34633\,
            I => \N__34616\
        );

    \I__6978\ : LocalMux
    port map (
            O => \N__34630\,
            I => \N__34616\
        );

    \I__6977\ : LocalMux
    port map (
            O => \N__34627\,
            I => measured_delay_hc_11
        );

    \I__6976\ : Odrv4
    port map (
            O => \N__34624\,
            I => measured_delay_hc_11
        );

    \I__6975\ : LocalMux
    port map (
            O => \N__34621\,
            I => measured_delay_hc_11
        );

    \I__6974\ : Odrv4
    port map (
            O => \N__34616\,
            I => measured_delay_hc_11
        );

    \I__6973\ : CascadeMux
    port map (
            O => \N__34607\,
            I => \N__34603\
        );

    \I__6972\ : CascadeMux
    port map (
            O => \N__34606\,
            I => \N__34600\
        );

    \I__6971\ : InMux
    port map (
            O => \N__34603\,
            I => \N__34597\
        );

    \I__6970\ : InMux
    port map (
            O => \N__34600\,
            I => \N__34592\
        );

    \I__6969\ : LocalMux
    port map (
            O => \N__34597\,
            I => \N__34589\
        );

    \I__6968\ : InMux
    port map (
            O => \N__34596\,
            I => \N__34586\
        );

    \I__6967\ : InMux
    port map (
            O => \N__34595\,
            I => \N__34583\
        );

    \I__6966\ : LocalMux
    port map (
            O => \N__34592\,
            I => \N__34578\
        );

    \I__6965\ : Span4Mux_v
    port map (
            O => \N__34589\,
            I => \N__34578\
        );

    \I__6964\ : LocalMux
    port map (
            O => \N__34586\,
            I => \N__34575\
        );

    \I__6963\ : LocalMux
    port map (
            O => \N__34583\,
            I => \N__34572\
        );

    \I__6962\ : Odrv4
    port map (
            O => \N__34578\,
            I => measured_delay_hc_2
        );

    \I__6961\ : Odrv12
    port map (
            O => \N__34575\,
            I => measured_delay_hc_2
        );

    \I__6960\ : Odrv4
    port map (
            O => \N__34572\,
            I => measured_delay_hc_2
        );

    \I__6959\ : CascadeMux
    port map (
            O => \N__34565\,
            I => \N__34562\
        );

    \I__6958\ : InMux
    port map (
            O => \N__34562\,
            I => \N__34558\
        );

    \I__6957\ : InMux
    port map (
            O => \N__34561\,
            I => \N__34553\
        );

    \I__6956\ : LocalMux
    port map (
            O => \N__34558\,
            I => \N__34550\
        );

    \I__6955\ : InMux
    port map (
            O => \N__34557\,
            I => \N__34547\
        );

    \I__6954\ : InMux
    port map (
            O => \N__34556\,
            I => \N__34544\
        );

    \I__6953\ : LocalMux
    port map (
            O => \N__34553\,
            I => \N__34540\
        );

    \I__6952\ : Span4Mux_v
    port map (
            O => \N__34550\,
            I => \N__34533\
        );

    \I__6951\ : LocalMux
    port map (
            O => \N__34547\,
            I => \N__34533\
        );

    \I__6950\ : LocalMux
    port map (
            O => \N__34544\,
            I => \N__34533\
        );

    \I__6949\ : InMux
    port map (
            O => \N__34543\,
            I => \N__34530\
        );

    \I__6948\ : Span4Mux_h
    port map (
            O => \N__34540\,
            I => \N__34527\
        );

    \I__6947\ : Span4Mux_v
    port map (
            O => \N__34533\,
            I => \N__34524\
        );

    \I__6946\ : LocalMux
    port map (
            O => \N__34530\,
            I => measured_delay_hc_7
        );

    \I__6945\ : Odrv4
    port map (
            O => \N__34527\,
            I => measured_delay_hc_7
        );

    \I__6944\ : Odrv4
    port map (
            O => \N__34524\,
            I => measured_delay_hc_7
        );

    \I__6943\ : InMux
    port map (
            O => \N__34517\,
            I => \N__34514\
        );

    \I__6942\ : LocalMux
    port map (
            O => \N__34514\,
            I => \N__34508\
        );

    \I__6941\ : InMux
    port map (
            O => \N__34513\,
            I => \N__34505\
        );

    \I__6940\ : InMux
    port map (
            O => \N__34512\,
            I => \N__34502\
        );

    \I__6939\ : InMux
    port map (
            O => \N__34511\,
            I => \N__34499\
        );

    \I__6938\ : Span12Mux_h
    port map (
            O => \N__34508\,
            I => \N__34492\
        );

    \I__6937\ : LocalMux
    port map (
            O => \N__34505\,
            I => \N__34492\
        );

    \I__6936\ : LocalMux
    port map (
            O => \N__34502\,
            I => \N__34492\
        );

    \I__6935\ : LocalMux
    port map (
            O => \N__34499\,
            I => measured_delay_hc_5
        );

    \I__6934\ : Odrv12
    port map (
            O => \N__34492\,
            I => measured_delay_hc_5
        );

    \I__6933\ : InMux
    port map (
            O => \N__34487\,
            I => \N__34483\
        );

    \I__6932\ : InMux
    port map (
            O => \N__34486\,
            I => \N__34480\
        );

    \I__6931\ : LocalMux
    port map (
            O => \N__34483\,
            I => \N__34477\
        );

    \I__6930\ : LocalMux
    port map (
            O => \N__34480\,
            I => measured_delay_hc_23
        );

    \I__6929\ : Odrv4
    port map (
            O => \N__34477\,
            I => measured_delay_hc_23
        );

    \I__6928\ : InMux
    port map (
            O => \N__34472\,
            I => \N__34469\
        );

    \I__6927\ : LocalMux
    port map (
            O => \N__34469\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_3\
        );

    \I__6926\ : CascadeMux
    port map (
            O => \N__34466\,
            I => \phase_controller_inst1.start_timer_hc_0_sqmuxa_cascade_\
        );

    \I__6925\ : InMux
    port map (
            O => \N__34463\,
            I => \N__34460\
        );

    \I__6924\ : LocalMux
    port map (
            O => \N__34460\,
            I => \phase_controller_inst1.start_timer_hc_RNOZ0Z_0\
        );

    \I__6923\ : InMux
    port map (
            O => \N__34457\,
            I => \N__34454\
        );

    \I__6922\ : LocalMux
    port map (
            O => \N__34454\,
            I => \N__34447\
        );

    \I__6921\ : InMux
    port map (
            O => \N__34453\,
            I => \N__34444\
        );

    \I__6920\ : InMux
    port map (
            O => \N__34452\,
            I => \N__34439\
        );

    \I__6919\ : InMux
    port map (
            O => \N__34451\,
            I => \N__34439\
        );

    \I__6918\ : CascadeMux
    port map (
            O => \N__34450\,
            I => \N__34436\
        );

    \I__6917\ : Span4Mux_v
    port map (
            O => \N__34447\,
            I => \N__34431\
        );

    \I__6916\ : LocalMux
    port map (
            O => \N__34444\,
            I => \N__34431\
        );

    \I__6915\ : LocalMux
    port map (
            O => \N__34439\,
            I => \N__34428\
        );

    \I__6914\ : InMux
    port map (
            O => \N__34436\,
            I => \N__34425\
        );

    \I__6913\ : Span4Mux_v
    port map (
            O => \N__34431\,
            I => \N__34422\
        );

    \I__6912\ : Span4Mux_h
    port map (
            O => \N__34428\,
            I => \N__34419\
        );

    \I__6911\ : LocalMux
    port map (
            O => \N__34425\,
            I => \phase_controller_inst1.stateZ0Z_3\
        );

    \I__6910\ : Odrv4
    port map (
            O => \N__34422\,
            I => \phase_controller_inst1.stateZ0Z_3\
        );

    \I__6909\ : Odrv4
    port map (
            O => \N__34419\,
            I => \phase_controller_inst1.stateZ0Z_3\
        );

    \I__6908\ : InMux
    port map (
            O => \N__34412\,
            I => \N__34407\
        );

    \I__6907\ : InMux
    port map (
            O => \N__34411\,
            I => \N__34404\
        );

    \I__6906\ : InMux
    port map (
            O => \N__34410\,
            I => \N__34401\
        );

    \I__6905\ : LocalMux
    port map (
            O => \N__34407\,
            I => \N__34396\
        );

    \I__6904\ : LocalMux
    port map (
            O => \N__34404\,
            I => \N__34396\
        );

    \I__6903\ : LocalMux
    port map (
            O => \N__34401\,
            I => \N__34393\
        );

    \I__6902\ : Span4Mux_v
    port map (
            O => \N__34396\,
            I => \N__34390\
        );

    \I__6901\ : Span12Mux_v
    port map (
            O => \N__34393\,
            I => \N__34387\
        );

    \I__6900\ : Span4Mux_h
    port map (
            O => \N__34390\,
            I => \N__34384\
        );

    \I__6899\ : Odrv12
    port map (
            O => \N__34387\,
            I => \il_max_comp1_D2\
        );

    \I__6898\ : Odrv4
    port map (
            O => \N__34384\,
            I => \il_max_comp1_D2\
        );

    \I__6897\ : InMux
    port map (
            O => \N__34379\,
            I => \N__34375\
        );

    \I__6896\ : CascadeMux
    port map (
            O => \N__34378\,
            I => \N__34372\
        );

    \I__6895\ : LocalMux
    port map (
            O => \N__34375\,
            I => \N__34368\
        );

    \I__6894\ : InMux
    port map (
            O => \N__34372\,
            I => \N__34363\
        );

    \I__6893\ : InMux
    port map (
            O => \N__34371\,
            I => \N__34363\
        );

    \I__6892\ : Odrv4
    port map (
            O => \N__34368\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__6891\ : LocalMux
    port map (
            O => \N__34363\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__6890\ : CascadeMux
    port map (
            O => \N__34358\,
            I => \N__34355\
        );

    \I__6889\ : InMux
    port map (
            O => \N__34355\,
            I => \N__34352\
        );

    \I__6888\ : LocalMux
    port map (
            O => \N__34352\,
            I => \N__34349\
        );

    \I__6887\ : Odrv4
    port map (
            O => \N__34349\,
            I => \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa\
        );

    \I__6886\ : InMux
    port map (
            O => \N__34346\,
            I => \N__34342\
        );

    \I__6885\ : InMux
    port map (
            O => \N__34345\,
            I => \N__34337\
        );

    \I__6884\ : LocalMux
    port map (
            O => \N__34342\,
            I => \N__34334\
        );

    \I__6883\ : InMux
    port map (
            O => \N__34341\,
            I => \N__34329\
        );

    \I__6882\ : InMux
    port map (
            O => \N__34340\,
            I => \N__34329\
        );

    \I__6881\ : LocalMux
    port map (
            O => \N__34337\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__6880\ : Odrv4
    port map (
            O => \N__34334\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__6879\ : LocalMux
    port map (
            O => \N__34329\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__6878\ : InMux
    port map (
            O => \N__34322\,
            I => \N__34318\
        );

    \I__6877\ : InMux
    port map (
            O => \N__34321\,
            I => \N__34315\
        );

    \I__6876\ : LocalMux
    port map (
            O => \N__34318\,
            I => \N__34309\
        );

    \I__6875\ : LocalMux
    port map (
            O => \N__34315\,
            I => \N__34309\
        );

    \I__6874\ : InMux
    port map (
            O => \N__34314\,
            I => \N__34306\
        );

    \I__6873\ : Span4Mux_h
    port map (
            O => \N__34309\,
            I => \N__34303\
        );

    \I__6872\ : LocalMux
    port map (
            O => \N__34306\,
            I => \phase_controller_inst1.stoper_hc.time_passed11\
        );

    \I__6871\ : Odrv4
    port map (
            O => \N__34303\,
            I => \phase_controller_inst1.stoper_hc.time_passed11\
        );

    \I__6870\ : CascadeMux
    port map (
            O => \N__34298\,
            I => \phase_controller_inst1.stoper_hc.time_passed11_cascade_\
        );

    \I__6869\ : InMux
    port map (
            O => \N__34295\,
            I => \N__34287\
        );

    \I__6868\ : InMux
    port map (
            O => \N__34294\,
            I => \N__34287\
        );

    \I__6867\ : InMux
    port map (
            O => \N__34293\,
            I => \N__34280\
        );

    \I__6866\ : InMux
    port map (
            O => \N__34292\,
            I => \N__34280\
        );

    \I__6865\ : LocalMux
    port map (
            O => \N__34287\,
            I => \N__34277\
        );

    \I__6864\ : InMux
    port map (
            O => \N__34286\,
            I => \N__34274\
        );

    \I__6863\ : InMux
    port map (
            O => \N__34285\,
            I => \N__34271\
        );

    \I__6862\ : LocalMux
    port map (
            O => \N__34280\,
            I => \N__34268\
        );

    \I__6861\ : Odrv4
    port map (
            O => \N__34277\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__6860\ : LocalMux
    port map (
            O => \N__34274\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__34271\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__6858\ : Odrv4
    port map (
            O => \N__34268\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__6857\ : InMux
    port map (
            O => \N__34259\,
            I => \N__34256\
        );

    \I__6856\ : LocalMux
    port map (
            O => \N__34256\,
            I => \N__34253\
        );

    \I__6855\ : Span4Mux_h
    port map (
            O => \N__34253\,
            I => \N__34249\
        );

    \I__6854\ : InMux
    port map (
            O => \N__34252\,
            I => \N__34245\
        );

    \I__6853\ : Span4Mux_v
    port map (
            O => \N__34249\,
            I => \N__34242\
        );

    \I__6852\ : CascadeMux
    port map (
            O => \N__34248\,
            I => \N__34239\
        );

    \I__6851\ : LocalMux
    port map (
            O => \N__34245\,
            I => \N__34235\
        );

    \I__6850\ : Sp12to4
    port map (
            O => \N__34242\,
            I => \N__34232\
        );

    \I__6849\ : InMux
    port map (
            O => \N__34239\,
            I => \N__34227\
        );

    \I__6848\ : InMux
    port map (
            O => \N__34238\,
            I => \N__34227\
        );

    \I__6847\ : Odrv4
    port map (
            O => \N__34235\,
            I => \phase_controller_inst1.stoper_tr.time_passed11\
        );

    \I__6846\ : Odrv12
    port map (
            O => \N__34232\,
            I => \phase_controller_inst1.stoper_tr.time_passed11\
        );

    \I__6845\ : LocalMux
    port map (
            O => \N__34227\,
            I => \phase_controller_inst1.stoper_tr.time_passed11\
        );

    \I__6844\ : InMux
    port map (
            O => \N__34220\,
            I => \N__34216\
        );

    \I__6843\ : InMux
    port map (
            O => \N__34219\,
            I => \N__34213\
        );

    \I__6842\ : LocalMux
    port map (
            O => \N__34216\,
            I => \phase_controller_inst1.stoper_hc.un1_m2_eZ0Z_1\
        );

    \I__6841\ : LocalMux
    port map (
            O => \N__34213\,
            I => \phase_controller_inst1.stoper_hc.un1_m2_eZ0Z_1\
        );

    \I__6840\ : InMux
    port map (
            O => \N__34208\,
            I => \N__34205\
        );

    \I__6839\ : LocalMux
    port map (
            O => \N__34205\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7\
        );

    \I__6838\ : InMux
    port map (
            O => \N__34202\,
            I => \N__34196\
        );

    \I__6837\ : InMux
    port map (
            O => \N__34201\,
            I => \N__34196\
        );

    \I__6836\ : LocalMux
    port map (
            O => \N__34196\,
            I => \phase_controller_inst1.stoper_hc.un1_m2_eZ0Z_2\
        );

    \I__6835\ : InMux
    port map (
            O => \N__34193\,
            I => \N__34190\
        );

    \I__6834\ : LocalMux
    port map (
            O => \N__34190\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8\
        );

    \I__6833\ : InMux
    port map (
            O => \N__34187\,
            I => \N__34184\
        );

    \I__6832\ : LocalMux
    port map (
            O => \N__34184\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8\
        );

    \I__6831\ : CascadeMux
    port map (
            O => \N__34181\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_2_cascade_\
        );

    \I__6830\ : InMux
    port map (
            O => \N__34178\,
            I => \N__34173\
        );

    \I__6829\ : InMux
    port map (
            O => \N__34177\,
            I => \N__34170\
        );

    \I__6828\ : InMux
    port map (
            O => \N__34176\,
            I => \N__34167\
        );

    \I__6827\ : LocalMux
    port map (
            O => \N__34173\,
            I => \N__34162\
        );

    \I__6826\ : LocalMux
    port map (
            O => \N__34170\,
            I => \N__34162\
        );

    \I__6825\ : LocalMux
    port map (
            O => \N__34167\,
            I => \N__34159\
        );

    \I__6824\ : Span4Mux_h
    port map (
            O => \N__34162\,
            I => \N__34156\
        );

    \I__6823\ : Span4Mux_h
    port map (
            O => \N__34159\,
            I => \N__34153\
        );

    \I__6822\ : Sp12to4
    port map (
            O => \N__34156\,
            I => \N__34150\
        );

    \I__6821\ : Sp12to4
    port map (
            O => \N__34153\,
            I => \N__34145\
        );

    \I__6820\ : Span12Mux_v
    port map (
            O => \N__34150\,
            I => \N__34145\
        );

    \I__6819\ : Odrv12
    port map (
            O => \N__34145\,
            I => \il_min_comp1_D2\
        );

    \I__6818\ : InMux
    port map (
            O => \N__34142\,
            I => \N__34137\
        );

    \I__6817\ : InMux
    port map (
            O => \N__34141\,
            I => \N__34133\
        );

    \I__6816\ : InMux
    port map (
            O => \N__34140\,
            I => \N__34130\
        );

    \I__6815\ : LocalMux
    port map (
            O => \N__34137\,
            I => \N__34127\
        );

    \I__6814\ : InMux
    port map (
            O => \N__34136\,
            I => \N__34124\
        );

    \I__6813\ : LocalMux
    port map (
            O => \N__34133\,
            I => \N__34120\
        );

    \I__6812\ : LocalMux
    port map (
            O => \N__34130\,
            I => \N__34113\
        );

    \I__6811\ : Span4Mux_v
    port map (
            O => \N__34127\,
            I => \N__34113\
        );

    \I__6810\ : LocalMux
    port map (
            O => \N__34124\,
            I => \N__34113\
        );

    \I__6809\ : CascadeMux
    port map (
            O => \N__34123\,
            I => \N__34110\
        );

    \I__6808\ : Sp12to4
    port map (
            O => \N__34120\,
            I => \N__34105\
        );

    \I__6807\ : Sp12to4
    port map (
            O => \N__34113\,
            I => \N__34105\
        );

    \I__6806\ : InMux
    port map (
            O => \N__34110\,
            I => \N__34102\
        );

    \I__6805\ : Span12Mux_s11_v
    port map (
            O => \N__34105\,
            I => \N__34099\
        );

    \I__6804\ : LocalMux
    port map (
            O => \N__34102\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__6803\ : Odrv12
    port map (
            O => \N__34099\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__6802\ : InMux
    port map (
            O => \N__34094\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17\
        );

    \I__6801\ : InMux
    port map (
            O => \N__34091\,
            I => \N__34088\
        );

    \I__6800\ : LocalMux
    port map (
            O => \N__34088\,
            I => \N__34085\
        );

    \I__6799\ : Odrv4
    port map (
            O => \N__34085\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0\
        );

    \I__6798\ : InMux
    port map (
            O => \N__34082\,
            I => \N__34079\
        );

    \I__6797\ : LocalMux
    port map (
            O => \N__34079\,
            I => \N__34076\
        );

    \I__6796\ : Odrv4
    port map (
            O => \N__34076\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0\
        );

    \I__6795\ : IoInMux
    port map (
            O => \N__34073\,
            I => \N__34070\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__34070\,
            I => s2_phy_c
        );

    \I__6793\ : IoInMux
    port map (
            O => \N__34067\,
            I => \N__34064\
        );

    \I__6792\ : LocalMux
    port map (
            O => \N__34064\,
            I => \N__34061\
        );

    \I__6791\ : Span4Mux_s3_v
    port map (
            O => \N__34061\,
            I => \N__34058\
        );

    \I__6790\ : Odrv4
    port map (
            O => \N__34058\,
            I => \delay_measurement_inst.delay_hc_timer.N_335_i\
        );

    \I__6789\ : InMux
    port map (
            O => \N__34055\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\
        );

    \I__6788\ : InMux
    port map (
            O => \N__34052\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\
        );

    \I__6787\ : InMux
    port map (
            O => \N__34049\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\
        );

    \I__6786\ : InMux
    port map (
            O => \N__34046\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\
        );

    \I__6785\ : InMux
    port map (
            O => \N__34043\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\
        );

    \I__6784\ : InMux
    port map (
            O => \N__34040\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\
        );

    \I__6783\ : InMux
    port map (
            O => \N__34037\,
            I => \N__34034\
        );

    \I__6782\ : LocalMux
    port map (
            O => \N__34034\,
            I => \N__34031\
        );

    \I__6781\ : Odrv4
    port map (
            O => \N__34031\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16\
        );

    \I__6780\ : InMux
    port map (
            O => \N__34028\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\
        );

    \I__6779\ : InMux
    port map (
            O => \N__34025\,
            I => \bfn_13_26_0_\
        );

    \I__6778\ : InMux
    port map (
            O => \N__34022\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\
        );

    \I__6777\ : InMux
    port map (
            O => \N__34019\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\
        );

    \I__6776\ : InMux
    port map (
            O => \N__34016\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\
        );

    \I__6775\ : InMux
    port map (
            O => \N__34013\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\
        );

    \I__6774\ : InMux
    port map (
            O => \N__34010\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\
        );

    \I__6773\ : InMux
    port map (
            O => \N__34007\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\
        );

    \I__6772\ : InMux
    port map (
            O => \N__34004\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\
        );

    \I__6771\ : InMux
    port map (
            O => \N__34001\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\
        );

    \I__6770\ : InMux
    port map (
            O => \N__33998\,
            I => \bfn_13_25_0_\
        );

    \I__6769\ : InMux
    port map (
            O => \N__33995\,
            I => \N__33991\
        );

    \I__6768\ : InMux
    port map (
            O => \N__33994\,
            I => \N__33988\
        );

    \I__6767\ : LocalMux
    port map (
            O => \N__33991\,
            I => \N__33984\
        );

    \I__6766\ : LocalMux
    port map (
            O => \N__33988\,
            I => \N__33981\
        );

    \I__6765\ : InMux
    port map (
            O => \N__33987\,
            I => \N__33978\
        );

    \I__6764\ : Span4Mux_v
    port map (
            O => \N__33984\,
            I => \N__33975\
        );

    \I__6763\ : Span4Mux_h
    port map (
            O => \N__33981\,
            I => \N__33972\
        );

    \I__6762\ : LocalMux
    port map (
            O => \N__33978\,
            I => \N__33969\
        );

    \I__6761\ : Span4Mux_v
    port map (
            O => \N__33975\,
            I => \N__33966\
        );

    \I__6760\ : Span4Mux_v
    port map (
            O => \N__33972\,
            I => \N__33961\
        );

    \I__6759\ : Span4Mux_v
    port map (
            O => \N__33969\,
            I => \N__33961\
        );

    \I__6758\ : Span4Mux_v
    port map (
            O => \N__33966\,
            I => \N__33958\
        );

    \I__6757\ : Span4Mux_v
    port map (
            O => \N__33961\,
            I => \N__33955\
        );

    \I__6756\ : Odrv4
    port map (
            O => \N__33958\,
            I => \il_min_comp2_D2\
        );

    \I__6755\ : Odrv4
    port map (
            O => \N__33955\,
            I => \il_min_comp2_D2\
        );

    \I__6754\ : InMux
    port map (
            O => \N__33950\,
            I => \N__33946\
        );

    \I__6753\ : CascadeMux
    port map (
            O => \N__33949\,
            I => \N__33942\
        );

    \I__6752\ : LocalMux
    port map (
            O => \N__33946\,
            I => \N__33938\
        );

    \I__6751\ : InMux
    port map (
            O => \N__33945\,
            I => \N__33935\
        );

    \I__6750\ : InMux
    port map (
            O => \N__33942\,
            I => \N__33930\
        );

    \I__6749\ : InMux
    port map (
            O => \N__33941\,
            I => \N__33930\
        );

    \I__6748\ : Span4Mux_h
    port map (
            O => \N__33938\,
            I => \N__33927\
        );

    \I__6747\ : LocalMux
    port map (
            O => \N__33935\,
            I => \phase_controller_slave.stateZ0Z_1\
        );

    \I__6746\ : LocalMux
    port map (
            O => \N__33930\,
            I => \phase_controller_slave.stateZ0Z_1\
        );

    \I__6745\ : Odrv4
    port map (
            O => \N__33927\,
            I => \phase_controller_slave.stateZ0Z_1\
        );

    \I__6744\ : CascadeMux
    port map (
            O => \N__33920\,
            I => \N__33917\
        );

    \I__6743\ : InMux
    port map (
            O => \N__33917\,
            I => \N__33914\
        );

    \I__6742\ : LocalMux
    port map (
            O => \N__33914\,
            I => \N__33911\
        );

    \I__6741\ : Odrv4
    port map (
            O => \N__33911\,
            I => \phase_controller_slave.start_timer_tr_0_sqmuxa\
        );

    \I__6740\ : InMux
    port map (
            O => \N__33908\,
            I => \N__33905\
        );

    \I__6739\ : LocalMux
    port map (
            O => \N__33905\,
            I => \phase_controller_slave.state_RNIVDE2Z0Z_0\
        );

    \I__6738\ : IoInMux
    port map (
            O => \N__33902\,
            I => \N__33899\
        );

    \I__6737\ : LocalMux
    port map (
            O => \N__33899\,
            I => \N__33896\
        );

    \I__6736\ : IoSpan4Mux
    port map (
            O => \N__33896\,
            I => \N__33892\
        );

    \I__6735\ : InMux
    port map (
            O => \N__33895\,
            I => \N__33889\
        );

    \I__6734\ : Span4Mux_s3_v
    port map (
            O => \N__33892\,
            I => \N__33884\
        );

    \I__6733\ : LocalMux
    port map (
            O => \N__33889\,
            I => \N__33884\
        );

    \I__6732\ : Span4Mux_v
    port map (
            O => \N__33884\,
            I => \N__33880\
        );

    \I__6731\ : InMux
    port map (
            O => \N__33883\,
            I => \N__33877\
        );

    \I__6730\ : Odrv4
    port map (
            O => \N__33880\,
            I => s3_phy_c
        );

    \I__6729\ : LocalMux
    port map (
            O => \N__33877\,
            I => s3_phy_c
        );

    \I__6728\ : CascadeMux
    port map (
            O => \N__33872\,
            I => \N__33868\
        );

    \I__6727\ : CascadeMux
    port map (
            O => \N__33871\,
            I => \N__33865\
        );

    \I__6726\ : InMux
    port map (
            O => \N__33868\,
            I => \N__33861\
        );

    \I__6725\ : InMux
    port map (
            O => \N__33865\,
            I => \N__33856\
        );

    \I__6724\ : InMux
    port map (
            O => \N__33864\,
            I => \N__33856\
        );

    \I__6723\ : LocalMux
    port map (
            O => \N__33861\,
            I => shift_flag_start
        );

    \I__6722\ : LocalMux
    port map (
            O => \N__33856\,
            I => shift_flag_start
        );

    \I__6721\ : InMux
    port map (
            O => \N__33851\,
            I => \N__33848\
        );

    \I__6720\ : LocalMux
    port map (
            O => \N__33848\,
            I => \N__33845\
        );

    \I__6719\ : Sp12to4
    port map (
            O => \N__33845\,
            I => \N__33841\
        );

    \I__6718\ : InMux
    port map (
            O => \N__33844\,
            I => \N__33838\
        );

    \I__6717\ : Odrv12
    port map (
            O => \N__33841\,
            I => \phase_controller_inst1.state_RNI7NN7Z0Z_0\
        );

    \I__6716\ : LocalMux
    port map (
            O => \N__33838\,
            I => \phase_controller_inst1.state_RNI7NN7Z0Z_0\
        );

    \I__6715\ : CascadeMux
    port map (
            O => \N__33833\,
            I => \N__33830\
        );

    \I__6714\ : InMux
    port map (
            O => \N__33830\,
            I => \N__33827\
        );

    \I__6713\ : LocalMux
    port map (
            O => \N__33827\,
            I => \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa\
        );

    \I__6712\ : InMux
    port map (
            O => \N__33824\,
            I => \N__33821\
        );

    \I__6711\ : LocalMux
    port map (
            O => \N__33821\,
            I => \phase_controller_inst1.start_timer_tr_0_sqmuxa\
        );

    \I__6710\ : CascadeMux
    port map (
            O => \N__33818\,
            I => \N__33814\
        );

    \I__6709\ : InMux
    port map (
            O => \N__33817\,
            I => \N__33806\
        );

    \I__6708\ : InMux
    port map (
            O => \N__33814\,
            I => \N__33806\
        );

    \I__6707\ : InMux
    port map (
            O => \N__33813\,
            I => \N__33806\
        );

    \I__6706\ : LocalMux
    port map (
            O => \N__33806\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__6705\ : InMux
    port map (
            O => \N__33803\,
            I => \N__33797\
        );

    \I__6704\ : InMux
    port map (
            O => \N__33802\,
            I => \N__33797\
        );

    \I__6703\ : LocalMux
    port map (
            O => \N__33797\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__6702\ : CascadeMux
    port map (
            O => \N__33794\,
            I => \N__33791\
        );

    \I__6701\ : InMux
    port map (
            O => \N__33791\,
            I => \N__33788\
        );

    \I__6700\ : LocalMux
    port map (
            O => \N__33788\,
            I => \N__33785\
        );

    \I__6699\ : Span4Mux_h
    port map (
            O => \N__33785\,
            I => \N__33782\
        );

    \I__6698\ : Odrv4
    port map (
            O => \N__33782\,
            I => \phase_controller_slave.stoper_tr.time_passed_1_sqmuxa\
        );

    \I__6697\ : CascadeMux
    port map (
            O => \N__33779\,
            I => \N__33775\
        );

    \I__6696\ : InMux
    port map (
            O => \N__33778\,
            I => \N__33771\
        );

    \I__6695\ : InMux
    port map (
            O => \N__33775\,
            I => \N__33766\
        );

    \I__6694\ : InMux
    port map (
            O => \N__33774\,
            I => \N__33766\
        );

    \I__6693\ : LocalMux
    port map (
            O => \N__33771\,
            I => \phase_controller_slave.tr_time_passed\
        );

    \I__6692\ : LocalMux
    port map (
            O => \N__33766\,
            I => \phase_controller_slave.tr_time_passed\
        );

    \I__6691\ : InMux
    port map (
            O => \N__33761\,
            I => \N__33755\
        );

    \I__6690\ : InMux
    port map (
            O => \N__33760\,
            I => \N__33755\
        );

    \I__6689\ : LocalMux
    port map (
            O => \N__33755\,
            I => \phase_controller_slave.stateZ0Z_0\
        );

    \I__6688\ : CascadeMux
    port map (
            O => \N__33752\,
            I => \phase_controller_slave.state_RNIVDE2Z0Z_0_cascade_\
        );

    \I__6687\ : InMux
    port map (
            O => \N__33749\,
            I => \N__33746\
        );

    \I__6686\ : LocalMux
    port map (
            O => \N__33746\,
            I => \N__33743\
        );

    \I__6685\ : Span4Mux_h
    port map (
            O => \N__33743\,
            I => \N__33739\
        );

    \I__6684\ : InMux
    port map (
            O => \N__33742\,
            I => \N__33736\
        );

    \I__6683\ : Odrv4
    port map (
            O => \N__33739\,
            I => state_ns_i_a2_1
        );

    \I__6682\ : LocalMux
    port map (
            O => \N__33736\,
            I => state_ns_i_a2_1
        );

    \I__6681\ : InMux
    port map (
            O => \N__33731\,
            I => \N__33726\
        );

    \I__6680\ : InMux
    port map (
            O => \N__33730\,
            I => \N__33723\
        );

    \I__6679\ : InMux
    port map (
            O => \N__33729\,
            I => \N__33719\
        );

    \I__6678\ : LocalMux
    port map (
            O => \N__33726\,
            I => \N__33715\
        );

    \I__6677\ : LocalMux
    port map (
            O => \N__33723\,
            I => \N__33712\
        );

    \I__6676\ : CascadeMux
    port map (
            O => \N__33722\,
            I => \N__33709\
        );

    \I__6675\ : LocalMux
    port map (
            O => \N__33719\,
            I => \N__33706\
        );

    \I__6674\ : InMux
    port map (
            O => \N__33718\,
            I => \N__33703\
        );

    \I__6673\ : Span4Mux_v
    port map (
            O => \N__33715\,
            I => \N__33700\
        );

    \I__6672\ : Span4Mux_h
    port map (
            O => \N__33712\,
            I => \N__33697\
        );

    \I__6671\ : InMux
    port map (
            O => \N__33709\,
            I => \N__33694\
        );

    \I__6670\ : Span4Mux_h
    port map (
            O => \N__33706\,
            I => \N__33688\
        );

    \I__6669\ : LocalMux
    port map (
            O => \N__33703\,
            I => \N__33688\
        );

    \I__6668\ : Span4Mux_h
    port map (
            O => \N__33700\,
            I => \N__33683\
        );

    \I__6667\ : Span4Mux_v
    port map (
            O => \N__33697\,
            I => \N__33683\
        );

    \I__6666\ : LocalMux
    port map (
            O => \N__33694\,
            I => \N__33680\
        );

    \I__6665\ : InMux
    port map (
            O => \N__33693\,
            I => \N__33677\
        );

    \I__6664\ : Span4Mux_v
    port map (
            O => \N__33688\,
            I => \N__33674\
        );

    \I__6663\ : Sp12to4
    port map (
            O => \N__33683\,
            I => \N__33671\
        );

    \I__6662\ : Span4Mux_h
    port map (
            O => \N__33680\,
            I => \N__33668\
        );

    \I__6661\ : LocalMux
    port map (
            O => \N__33677\,
            I => \N__33665\
        );

    \I__6660\ : Span4Mux_h
    port map (
            O => \N__33674\,
            I => \N__33662\
        );

    \I__6659\ : Span12Mux_v
    port map (
            O => \N__33671\,
            I => \N__33655\
        );

    \I__6658\ : Sp12to4
    port map (
            O => \N__33668\,
            I => \N__33655\
        );

    \I__6657\ : Sp12to4
    port map (
            O => \N__33665\,
            I => \N__33655\
        );

    \I__6656\ : Sp12to4
    port map (
            O => \N__33662\,
            I => \N__33652\
        );

    \I__6655\ : Span12Mux_v
    port map (
            O => \N__33655\,
            I => \N__33649\
        );

    \I__6654\ : Span12Mux_v
    port map (
            O => \N__33652\,
            I => \N__33644\
        );

    \I__6653\ : Span12Mux_h
    port map (
            O => \N__33649\,
            I => \N__33644\
        );

    \I__6652\ : Odrv12
    port map (
            O => \N__33644\,
            I => start_stop_c
        );

    \I__6651\ : IoInMux
    port map (
            O => \N__33641\,
            I => \N__33638\
        );

    \I__6650\ : LocalMux
    port map (
            O => \N__33638\,
            I => \N__33635\
        );

    \I__6649\ : Span4Mux_s3_v
    port map (
            O => \N__33635\,
            I => \N__33632\
        );

    \I__6648\ : Span4Mux_h
    port map (
            O => \N__33632\,
            I => \N__33629\
        );

    \I__6647\ : Span4Mux_v
    port map (
            O => \N__33629\,
            I => \N__33626\
        );

    \I__6646\ : Span4Mux_v
    port map (
            O => \N__33626\,
            I => \N__33622\
        );

    \I__6645\ : InMux
    port map (
            O => \N__33625\,
            I => \N__33619\
        );

    \I__6644\ : Odrv4
    port map (
            O => \N__33622\,
            I => s4_phy_c
        );

    \I__6643\ : LocalMux
    port map (
            O => \N__33619\,
            I => s4_phy_c
        );

    \I__6642\ : CascadeMux
    port map (
            O => \N__33614\,
            I => \N__33611\
        );

    \I__6641\ : InMux
    port map (
            O => \N__33611\,
            I => \N__33608\
        );

    \I__6640\ : LocalMux
    port map (
            O => \N__33608\,
            I => \N__33605\
        );

    \I__6639\ : Span4Mux_v
    port map (
            O => \N__33605\,
            I => \N__33602\
        );

    \I__6638\ : Odrv4
    port map (
            O => \N__33602\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\
        );

    \I__6637\ : CascadeMux
    port map (
            O => \N__33599\,
            I => \N__33596\
        );

    \I__6636\ : InMux
    port map (
            O => \N__33596\,
            I => \N__33593\
        );

    \I__6635\ : LocalMux
    port map (
            O => \N__33593\,
            I => \N__33590\
        );

    \I__6634\ : Odrv4
    port map (
            O => \N__33590\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\
        );

    \I__6633\ : CascadeMux
    port map (
            O => \N__33587\,
            I => \N__33584\
        );

    \I__6632\ : InMux
    port map (
            O => \N__33584\,
            I => \N__33581\
        );

    \I__6631\ : LocalMux
    port map (
            O => \N__33581\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\
        );

    \I__6630\ : CascadeMux
    port map (
            O => \N__33578\,
            I => \N__33575\
        );

    \I__6629\ : InMux
    port map (
            O => \N__33575\,
            I => \N__33572\
        );

    \I__6628\ : LocalMux
    port map (
            O => \N__33572\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\
        );

    \I__6627\ : CEMux
    port map (
            O => \N__33569\,
            I => \N__33566\
        );

    \I__6626\ : LocalMux
    port map (
            O => \N__33566\,
            I => \N__33562\
        );

    \I__6625\ : CEMux
    port map (
            O => \N__33565\,
            I => \N__33558\
        );

    \I__6624\ : Span4Mux_h
    port map (
            O => \N__33562\,
            I => \N__33553\
        );

    \I__6623\ : CEMux
    port map (
            O => \N__33561\,
            I => \N__33550\
        );

    \I__6622\ : LocalMux
    port map (
            O => \N__33558\,
            I => \N__33547\
        );

    \I__6621\ : CEMux
    port map (
            O => \N__33557\,
            I => \N__33544\
        );

    \I__6620\ : CEMux
    port map (
            O => \N__33556\,
            I => \N__33541\
        );

    \I__6619\ : Span4Mux_h
    port map (
            O => \N__33553\,
            I => \N__33537\
        );

    \I__6618\ : LocalMux
    port map (
            O => \N__33550\,
            I => \N__33534\
        );

    \I__6617\ : Span4Mux_v
    port map (
            O => \N__33547\,
            I => \N__33529\
        );

    \I__6616\ : LocalMux
    port map (
            O => \N__33544\,
            I => \N__33529\
        );

    \I__6615\ : LocalMux
    port map (
            O => \N__33541\,
            I => \N__33526\
        );

    \I__6614\ : CEMux
    port map (
            O => \N__33540\,
            I => \N__33523\
        );

    \I__6613\ : Span4Mux_h
    port map (
            O => \N__33537\,
            I => \N__33518\
        );

    \I__6612\ : Span4Mux_v
    port map (
            O => \N__33534\,
            I => \N__33518\
        );

    \I__6611\ : Span4Mux_h
    port map (
            O => \N__33529\,
            I => \N__33515\
        );

    \I__6610\ : Span4Mux_h
    port map (
            O => \N__33526\,
            I => \N__33512\
        );

    \I__6609\ : LocalMux
    port map (
            O => \N__33523\,
            I => \N__33509\
        );

    \I__6608\ : Span4Mux_v
    port map (
            O => \N__33518\,
            I => \N__33504\
        );

    \I__6607\ : Span4Mux_v
    port map (
            O => \N__33515\,
            I => \N__33504\
        );

    \I__6606\ : Span4Mux_v
    port map (
            O => \N__33512\,
            I => \N__33499\
        );

    \I__6605\ : Span4Mux_h
    port map (
            O => \N__33509\,
            I => \N__33499\
        );

    \I__6604\ : Odrv4
    port map (
            O => \N__33504\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__6603\ : Odrv4
    port map (
            O => \N__33499\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__6602\ : CascadeMux
    port map (
            O => \N__33494\,
            I => \N__33491\
        );

    \I__6601\ : InMux
    port map (
            O => \N__33491\,
            I => \N__33488\
        );

    \I__6600\ : LocalMux
    port map (
            O => \N__33488\,
            I => \N__33485\
        );

    \I__6599\ : Odrv4
    port map (
            O => \N__33485\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\
        );

    \I__6598\ : InMux
    port map (
            O => \N__33482\,
            I => \N__33479\
        );

    \I__6597\ : LocalMux
    port map (
            O => \N__33479\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_16\
        );

    \I__6596\ : InMux
    port map (
            O => \N__33476\,
            I => \N__33473\
        );

    \I__6595\ : LocalMux
    port map (
            O => \N__33473\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_17\
        );

    \I__6594\ : InMux
    port map (
            O => \N__33470\,
            I => \N__33467\
        );

    \I__6593\ : LocalMux
    port map (
            O => \N__33467\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_18\
        );

    \I__6592\ : CascadeMux
    port map (
            O => \N__33464\,
            I => \N__33461\
        );

    \I__6591\ : InMux
    port map (
            O => \N__33461\,
            I => \N__33458\
        );

    \I__6590\ : LocalMux
    port map (
            O => \N__33458\,
            I => \N__33455\
        );

    \I__6589\ : Span4Mux_h
    port map (
            O => \N__33455\,
            I => \N__33452\
        );

    \I__6588\ : Odrv4
    port map (
            O => \N__33452\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\
        );

    \I__6587\ : InMux
    port map (
            O => \N__33449\,
            I => \N__33446\
        );

    \I__6586\ : LocalMux
    port map (
            O => \N__33446\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_19\
        );

    \I__6585\ : InMux
    port map (
            O => \N__33443\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__6584\ : InMux
    port map (
            O => \N__33440\,
            I => \N__33437\
        );

    \I__6583\ : LocalMux
    port map (
            O => \N__33437\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0\
        );

    \I__6582\ : CascadeMux
    port map (
            O => \N__33434\,
            I => \N__33431\
        );

    \I__6581\ : InMux
    port map (
            O => \N__33431\,
            I => \N__33428\
        );

    \I__6580\ : LocalMux
    port map (
            O => \N__33428\,
            I => \N__33425\
        );

    \I__6579\ : Odrv4
    port map (
            O => \N__33425\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\
        );

    \I__6578\ : InMux
    port map (
            O => \N__33422\,
            I => \N__33419\
        );

    \I__6577\ : LocalMux
    port map (
            O => \N__33419\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\
        );

    \I__6576\ : CascadeMux
    port map (
            O => \N__33416\,
            I => \N__33413\
        );

    \I__6575\ : InMux
    port map (
            O => \N__33413\,
            I => \N__33410\
        );

    \I__6574\ : LocalMux
    port map (
            O => \N__33410\,
            I => \N__33407\
        );

    \I__6573\ : Span4Mux_v
    port map (
            O => \N__33407\,
            I => \N__33404\
        );

    \I__6572\ : Span4Mux_v
    port map (
            O => \N__33404\,
            I => \N__33401\
        );

    \I__6571\ : Span4Mux_h
    port map (
            O => \N__33401\,
            I => \N__33398\
        );

    \I__6570\ : Span4Mux_h
    port map (
            O => \N__33398\,
            I => \N__33395\
        );

    \I__6569\ : Odrv4
    port map (
            O => \N__33395\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\
        );

    \I__6568\ : InMux
    port map (
            O => \N__33392\,
            I => \N__33389\
        );

    \I__6567\ : LocalMux
    port map (
            O => \N__33389\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\
        );

    \I__6566\ : CascadeMux
    port map (
            O => \N__33386\,
            I => \N__33383\
        );

    \I__6565\ : InMux
    port map (
            O => \N__33383\,
            I => \N__33380\
        );

    \I__6564\ : LocalMux
    port map (
            O => \N__33380\,
            I => \N__33377\
        );

    \I__6563\ : Sp12to4
    port map (
            O => \N__33377\,
            I => \N__33374\
        );

    \I__6562\ : Span12Mux_h
    port map (
            O => \N__33374\,
            I => \N__33371\
        );

    \I__6561\ : Odrv12
    port map (
            O => \N__33371\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\
        );

    \I__6560\ : InMux
    port map (
            O => \N__33368\,
            I => \N__33365\
        );

    \I__6559\ : LocalMux
    port map (
            O => \N__33365\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\
        );

    \I__6558\ : CascadeMux
    port map (
            O => \N__33362\,
            I => \N__33359\
        );

    \I__6557\ : InMux
    port map (
            O => \N__33359\,
            I => \N__33356\
        );

    \I__6556\ : LocalMux
    port map (
            O => \N__33356\,
            I => \N__33353\
        );

    \I__6555\ : Odrv4
    port map (
            O => \N__33353\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\
        );

    \I__6554\ : InMux
    port map (
            O => \N__33350\,
            I => \N__33347\
        );

    \I__6553\ : LocalMux
    port map (
            O => \N__33347\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\
        );

    \I__6552\ : InMux
    port map (
            O => \N__33344\,
            I => \N__33341\
        );

    \I__6551\ : LocalMux
    port map (
            O => \N__33341\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\
        );

    \I__6550\ : CascadeMux
    port map (
            O => \N__33338\,
            I => \N__33335\
        );

    \I__6549\ : InMux
    port map (
            O => \N__33335\,
            I => \N__33332\
        );

    \I__6548\ : LocalMux
    port map (
            O => \N__33332\,
            I => \N__33329\
        );

    \I__6547\ : Span4Mux_v
    port map (
            O => \N__33329\,
            I => \N__33326\
        );

    \I__6546\ : Odrv4
    port map (
            O => \N__33326\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\
        );

    \I__6545\ : InMux
    port map (
            O => \N__33323\,
            I => \N__33320\
        );

    \I__6544\ : LocalMux
    port map (
            O => \N__33320\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\
        );

    \I__6543\ : CascadeMux
    port map (
            O => \N__33317\,
            I => \N__33314\
        );

    \I__6542\ : InMux
    port map (
            O => \N__33314\,
            I => \N__33311\
        );

    \I__6541\ : LocalMux
    port map (
            O => \N__33311\,
            I => \N__33308\
        );

    \I__6540\ : Odrv12
    port map (
            O => \N__33308\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\
        );

    \I__6539\ : InMux
    port map (
            O => \N__33305\,
            I => \N__33302\
        );

    \I__6538\ : LocalMux
    port map (
            O => \N__33302\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\
        );

    \I__6537\ : InMux
    port map (
            O => \N__33299\,
            I => \N__33296\
        );

    \I__6536\ : LocalMux
    port map (
            O => \N__33296\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\
        );

    \I__6535\ : InMux
    port map (
            O => \N__33293\,
            I => \N__33290\
        );

    \I__6534\ : LocalMux
    port map (
            O => \N__33290\,
            I => \N__33287\
        );

    \I__6533\ : Span4Mux_v
    port map (
            O => \N__33287\,
            I => \N__33284\
        );

    \I__6532\ : Span4Mux_v
    port map (
            O => \N__33284\,
            I => \N__33281\
        );

    \I__6531\ : Sp12to4
    port map (
            O => \N__33281\,
            I => \N__33278\
        );

    \I__6530\ : Odrv12
    port map (
            O => \N__33278\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_0\
        );

    \I__6529\ : CascadeMux
    port map (
            O => \N__33275\,
            I => \N__33272\
        );

    \I__6528\ : InMux
    port map (
            O => \N__33272\,
            I => \N__33269\
        );

    \I__6527\ : LocalMux
    port map (
            O => \N__33269\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\
        );

    \I__6526\ : InMux
    port map (
            O => \N__33266\,
            I => \N__33263\
        );

    \I__6525\ : LocalMux
    port map (
            O => \N__33263\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\
        );

    \I__6524\ : CascadeMux
    port map (
            O => \N__33260\,
            I => \N__33257\
        );

    \I__6523\ : InMux
    port map (
            O => \N__33257\,
            I => \N__33254\
        );

    \I__6522\ : LocalMux
    port map (
            O => \N__33254\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\
        );

    \I__6521\ : InMux
    port map (
            O => \N__33251\,
            I => \N__33248\
        );

    \I__6520\ : LocalMux
    port map (
            O => \N__33248\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\
        );

    \I__6519\ : CascadeMux
    port map (
            O => \N__33245\,
            I => \N__33242\
        );

    \I__6518\ : InMux
    port map (
            O => \N__33242\,
            I => \N__33239\
        );

    \I__6517\ : LocalMux
    port map (
            O => \N__33239\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\
        );

    \I__6516\ : InMux
    port map (
            O => \N__33236\,
            I => \N__33233\
        );

    \I__6515\ : LocalMux
    port map (
            O => \N__33233\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\
        );

    \I__6514\ : InMux
    port map (
            O => \N__33230\,
            I => \N__33227\
        );

    \I__6513\ : LocalMux
    port map (
            O => \N__33227\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\
        );

    \I__6512\ : CascadeMux
    port map (
            O => \N__33224\,
            I => \N__33221\
        );

    \I__6511\ : InMux
    port map (
            O => \N__33221\,
            I => \N__33218\
        );

    \I__6510\ : LocalMux
    port map (
            O => \N__33218\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\
        );

    \I__6509\ : CascadeMux
    port map (
            O => \N__33215\,
            I => \N__33212\
        );

    \I__6508\ : InMux
    port map (
            O => \N__33212\,
            I => \N__33209\
        );

    \I__6507\ : LocalMux
    port map (
            O => \N__33209\,
            I => \N__33206\
        );

    \I__6506\ : Span4Mux_h
    port map (
            O => \N__33206\,
            I => \N__33203\
        );

    \I__6505\ : Odrv4
    port map (
            O => \N__33203\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\
        );

    \I__6504\ : InMux
    port map (
            O => \N__33200\,
            I => \N__33197\
        );

    \I__6503\ : LocalMux
    port map (
            O => \N__33197\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\
        );

    \I__6502\ : CascadeMux
    port map (
            O => \N__33194\,
            I => \N__33191\
        );

    \I__6501\ : InMux
    port map (
            O => \N__33191\,
            I => \N__33188\
        );

    \I__6500\ : LocalMux
    port map (
            O => \N__33188\,
            I => \N__33185\
        );

    \I__6499\ : Span4Mux_h
    port map (
            O => \N__33185\,
            I => \N__33182\
        );

    \I__6498\ : Odrv4
    port map (
            O => \N__33182\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ1Z_6\
        );

    \I__6497\ : InMux
    port map (
            O => \N__33179\,
            I => \N__33176\
        );

    \I__6496\ : LocalMux
    port map (
            O => \N__33176\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\
        );

    \I__6495\ : CascadeMux
    port map (
            O => \N__33173\,
            I => \N__33170\
        );

    \I__6494\ : InMux
    port map (
            O => \N__33170\,
            I => \N__33167\
        );

    \I__6493\ : LocalMux
    port map (
            O => \N__33167\,
            I => \N__33164\
        );

    \I__6492\ : Odrv4
    port map (
            O => \N__33164\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\
        );

    \I__6491\ : InMux
    port map (
            O => \N__33161\,
            I => \N__33158\
        );

    \I__6490\ : LocalMux
    port map (
            O => \N__33158\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\
        );

    \I__6489\ : InMux
    port map (
            O => \N__33155\,
            I => \N__33152\
        );

    \I__6488\ : LocalMux
    port map (
            O => \N__33152\,
            I => \N__33149\
        );

    \I__6487\ : Odrv4
    port map (
            O => \N__33149\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9\
        );

    \I__6486\ : InMux
    port map (
            O => \N__33146\,
            I => \N__33143\
        );

    \I__6485\ : LocalMux
    port map (
            O => \N__33143\,
            I => \N__33139\
        );

    \I__6484\ : InMux
    port map (
            O => \N__33142\,
            I => \N__33136\
        );

    \I__6483\ : Span4Mux_h
    port map (
            O => \N__33139\,
            I => \N__33131\
        );

    \I__6482\ : LocalMux
    port map (
            O => \N__33136\,
            I => \N__33131\
        );

    \I__6481\ : Span4Mux_v
    port map (
            O => \N__33131\,
            I => \N__33127\
        );

    \I__6480\ : InMux
    port map (
            O => \N__33130\,
            I => \N__33124\
        );

    \I__6479\ : Odrv4
    port map (
            O => \N__33127\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto30_2\
        );

    \I__6478\ : LocalMux
    port map (
            O => \N__33124\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto30_2\
        );

    \I__6477\ : InMux
    port map (
            O => \N__33119\,
            I => \N__33116\
        );

    \I__6476\ : LocalMux
    port map (
            O => \N__33116\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto8Z0Z_0\
        );

    \I__6475\ : InMux
    port map (
            O => \N__33113\,
            I => \N__33110\
        );

    \I__6474\ : LocalMux
    port map (
            O => \N__33110\,
            I => \phase_controller_inst1.stoper_hc.un1_m2_eZ0\
        );

    \I__6473\ : InMux
    port map (
            O => \N__33107\,
            I => \N__33104\
        );

    \I__6472\ : LocalMux
    port map (
            O => \N__33104\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_12\
        );

    \I__6471\ : CascadeMux
    port map (
            O => \N__33101\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_11_cascade_\
        );

    \I__6470\ : CascadeMux
    port map (
            O => \N__33098\,
            I => \phase_controller_inst1.stoper_hc.un2_startlt31_cascade_\
        );

    \I__6469\ : InMux
    port map (
            O => \N__33095\,
            I => \N__33092\
        );

    \I__6468\ : LocalMux
    port map (
            O => \N__33092\,
            I => \N__33089\
        );

    \I__6467\ : Span4Mux_h
    port map (
            O => \N__33089\,
            I => \N__33086\
        );

    \I__6466\ : Odrv4
    port map (
            O => \N__33086\,
            I => \il_max_comp2_D1\
        );

    \I__6465\ : InMux
    port map (
            O => \N__33083\,
            I => \N__33070\
        );

    \I__6464\ : InMux
    port map (
            O => \N__33082\,
            I => \N__33045\
        );

    \I__6463\ : InMux
    port map (
            O => \N__33081\,
            I => \N__33045\
        );

    \I__6462\ : InMux
    port map (
            O => \N__33080\,
            I => \N__33045\
        );

    \I__6461\ : InMux
    port map (
            O => \N__33079\,
            I => \N__33045\
        );

    \I__6460\ : InMux
    port map (
            O => \N__33078\,
            I => \N__33045\
        );

    \I__6459\ : InMux
    port map (
            O => \N__33077\,
            I => \N__33045\
        );

    \I__6458\ : InMux
    port map (
            O => \N__33076\,
            I => \N__33045\
        );

    \I__6457\ : InMux
    port map (
            O => \N__33075\,
            I => \N__33045\
        );

    \I__6456\ : InMux
    port map (
            O => \N__33074\,
            I => \N__33042\
        );

    \I__6455\ : CascadeMux
    port map (
            O => \N__33073\,
            I => \N__33038\
        );

    \I__6454\ : LocalMux
    port map (
            O => \N__33070\,
            I => \N__33031\
        );

    \I__6453\ : InMux
    port map (
            O => \N__33069\,
            I => \N__33028\
        );

    \I__6452\ : InMux
    port map (
            O => \N__33068\,
            I => \N__33015\
        );

    \I__6451\ : InMux
    port map (
            O => \N__33067\,
            I => \N__33015\
        );

    \I__6450\ : InMux
    port map (
            O => \N__33066\,
            I => \N__33015\
        );

    \I__6449\ : InMux
    port map (
            O => \N__33065\,
            I => \N__33015\
        );

    \I__6448\ : InMux
    port map (
            O => \N__33064\,
            I => \N__33015\
        );

    \I__6447\ : InMux
    port map (
            O => \N__33063\,
            I => \N__33015\
        );

    \I__6446\ : InMux
    port map (
            O => \N__33062\,
            I => \N__33012\
        );

    \I__6445\ : LocalMux
    port map (
            O => \N__33045\,
            I => \N__33000\
        );

    \I__6444\ : LocalMux
    port map (
            O => \N__33042\,
            I => \N__32997\
        );

    \I__6443\ : InMux
    port map (
            O => \N__33041\,
            I => \N__32994\
        );

    \I__6442\ : InMux
    port map (
            O => \N__33038\,
            I => \N__32991\
        );

    \I__6441\ : InMux
    port map (
            O => \N__33037\,
            I => \N__32982\
        );

    \I__6440\ : InMux
    port map (
            O => \N__33036\,
            I => \N__32982\
        );

    \I__6439\ : InMux
    port map (
            O => \N__33035\,
            I => \N__32982\
        );

    \I__6438\ : InMux
    port map (
            O => \N__33034\,
            I => \N__32982\
        );

    \I__6437\ : Span4Mux_v
    port map (
            O => \N__33031\,
            I => \N__32979\
        );

    \I__6436\ : LocalMux
    port map (
            O => \N__33028\,
            I => \N__32976\
        );

    \I__6435\ : LocalMux
    port map (
            O => \N__33015\,
            I => \N__32971\
        );

    \I__6434\ : LocalMux
    port map (
            O => \N__33012\,
            I => \N__32971\
        );

    \I__6433\ : InMux
    port map (
            O => \N__33011\,
            I => \N__32968\
        );

    \I__6432\ : InMux
    port map (
            O => \N__33010\,
            I => \N__32963\
        );

    \I__6431\ : InMux
    port map (
            O => \N__33009\,
            I => \N__32963\
        );

    \I__6430\ : InMux
    port map (
            O => \N__33008\,
            I => \N__32958\
        );

    \I__6429\ : InMux
    port map (
            O => \N__33007\,
            I => \N__32958\
        );

    \I__6428\ : InMux
    port map (
            O => \N__33006\,
            I => \N__32955\
        );

    \I__6427\ : InMux
    port map (
            O => \N__33005\,
            I => \N__32950\
        );

    \I__6426\ : InMux
    port map (
            O => \N__33004\,
            I => \N__32950\
        );

    \I__6425\ : InMux
    port map (
            O => \N__33003\,
            I => \N__32947\
        );

    \I__6424\ : Span4Mux_h
    port map (
            O => \N__33000\,
            I => \N__32944\
        );

    \I__6423\ : Span4Mux_h
    port map (
            O => \N__32997\,
            I => \N__32939\
        );

    \I__6422\ : LocalMux
    port map (
            O => \N__32994\,
            I => \N__32939\
        );

    \I__6421\ : LocalMux
    port map (
            O => \N__32991\,
            I => \N__32926\
        );

    \I__6420\ : LocalMux
    port map (
            O => \N__32982\,
            I => \N__32926\
        );

    \I__6419\ : Span4Mux_h
    port map (
            O => \N__32979\,
            I => \N__32926\
        );

    \I__6418\ : Span4Mux_v
    port map (
            O => \N__32976\,
            I => \N__32926\
        );

    \I__6417\ : Span4Mux_v
    port map (
            O => \N__32971\,
            I => \N__32926\
        );

    \I__6416\ : LocalMux
    port map (
            O => \N__32968\,
            I => \N__32926\
        );

    \I__6415\ : LocalMux
    port map (
            O => \N__32963\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__6414\ : LocalMux
    port map (
            O => \N__32958\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__6413\ : LocalMux
    port map (
            O => \N__32955\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__6412\ : LocalMux
    port map (
            O => \N__32950\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__6411\ : LocalMux
    port map (
            O => \N__32947\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__6410\ : Odrv4
    port map (
            O => \N__32944\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__6409\ : Odrv4
    port map (
            O => \N__32939\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__6408\ : Odrv4
    port map (
            O => \N__32926\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__6407\ : InMux
    port map (
            O => \N__32909\,
            I => \N__32904\
        );

    \I__6406\ : InMux
    port map (
            O => \N__32908\,
            I => \N__32901\
        );

    \I__6405\ : CascadeMux
    port map (
            O => \N__32907\,
            I => \N__32892\
        );

    \I__6404\ : LocalMux
    port map (
            O => \N__32904\,
            I => \N__32888\
        );

    \I__6403\ : LocalMux
    port map (
            O => \N__32901\,
            I => \N__32885\
        );

    \I__6402\ : InMux
    port map (
            O => \N__32900\,
            I => \N__32882\
        );

    \I__6401\ : InMux
    port map (
            O => \N__32899\,
            I => \N__32870\
        );

    \I__6400\ : InMux
    port map (
            O => \N__32898\,
            I => \N__32870\
        );

    \I__6399\ : InMux
    port map (
            O => \N__32897\,
            I => \N__32870\
        );

    \I__6398\ : InMux
    port map (
            O => \N__32896\,
            I => \N__32870\
        );

    \I__6397\ : InMux
    port map (
            O => \N__32895\,
            I => \N__32870\
        );

    \I__6396\ : InMux
    port map (
            O => \N__32892\,
            I => \N__32865\
        );

    \I__6395\ : InMux
    port map (
            O => \N__32891\,
            I => \N__32865\
        );

    \I__6394\ : Span4Mux_v
    port map (
            O => \N__32888\,
            I => \N__32852\
        );

    \I__6393\ : Span4Mux_h
    port map (
            O => \N__32885\,
            I => \N__32852\
        );

    \I__6392\ : LocalMux
    port map (
            O => \N__32882\,
            I => \N__32852\
        );

    \I__6391\ : InMux
    port map (
            O => \N__32881\,
            I => \N__32849\
        );

    \I__6390\ : LocalMux
    port map (
            O => \N__32870\,
            I => \N__32846\
        );

    \I__6389\ : LocalMux
    port map (
            O => \N__32865\,
            I => \N__32843\
        );

    \I__6388\ : CascadeMux
    port map (
            O => \N__32864\,
            I => \N__32831\
        );

    \I__6387\ : CascadeMux
    port map (
            O => \N__32863\,
            I => \N__32827\
        );

    \I__6386\ : CascadeMux
    port map (
            O => \N__32862\,
            I => \N__32822\
        );

    \I__6385\ : CascadeMux
    port map (
            O => \N__32861\,
            I => \N__32819\
        );

    \I__6384\ : CascadeMux
    port map (
            O => \N__32860\,
            I => \N__32816\
        );

    \I__6383\ : CascadeMux
    port map (
            O => \N__32859\,
            I => \N__32812\
        );

    \I__6382\ : Span4Mux_h
    port map (
            O => \N__32852\,
            I => \N__32807\
        );

    \I__6381\ : LocalMux
    port map (
            O => \N__32849\,
            I => \N__32804\
        );

    \I__6380\ : Span4Mux_v
    port map (
            O => \N__32846\,
            I => \N__32799\
        );

    \I__6379\ : Span4Mux_h
    port map (
            O => \N__32843\,
            I => \N__32799\
        );

    \I__6378\ : InMux
    port map (
            O => \N__32842\,
            I => \N__32790\
        );

    \I__6377\ : InMux
    port map (
            O => \N__32841\,
            I => \N__32790\
        );

    \I__6376\ : InMux
    port map (
            O => \N__32840\,
            I => \N__32790\
        );

    \I__6375\ : InMux
    port map (
            O => \N__32839\,
            I => \N__32790\
        );

    \I__6374\ : InMux
    port map (
            O => \N__32838\,
            I => \N__32783\
        );

    \I__6373\ : InMux
    port map (
            O => \N__32837\,
            I => \N__32783\
        );

    \I__6372\ : InMux
    port map (
            O => \N__32836\,
            I => \N__32783\
        );

    \I__6371\ : InMux
    port map (
            O => \N__32835\,
            I => \N__32770\
        );

    \I__6370\ : InMux
    port map (
            O => \N__32834\,
            I => \N__32770\
        );

    \I__6369\ : InMux
    port map (
            O => \N__32831\,
            I => \N__32770\
        );

    \I__6368\ : InMux
    port map (
            O => \N__32830\,
            I => \N__32770\
        );

    \I__6367\ : InMux
    port map (
            O => \N__32827\,
            I => \N__32770\
        );

    \I__6366\ : InMux
    port map (
            O => \N__32826\,
            I => \N__32770\
        );

    \I__6365\ : InMux
    port map (
            O => \N__32825\,
            I => \N__32753\
        );

    \I__6364\ : InMux
    port map (
            O => \N__32822\,
            I => \N__32753\
        );

    \I__6363\ : InMux
    port map (
            O => \N__32819\,
            I => \N__32753\
        );

    \I__6362\ : InMux
    port map (
            O => \N__32816\,
            I => \N__32753\
        );

    \I__6361\ : InMux
    port map (
            O => \N__32815\,
            I => \N__32753\
        );

    \I__6360\ : InMux
    port map (
            O => \N__32812\,
            I => \N__32753\
        );

    \I__6359\ : InMux
    port map (
            O => \N__32811\,
            I => \N__32753\
        );

    \I__6358\ : InMux
    port map (
            O => \N__32810\,
            I => \N__32753\
        );

    \I__6357\ : Odrv4
    port map (
            O => \N__32807\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__6356\ : Odrv4
    port map (
            O => \N__32804\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__6355\ : Odrv4
    port map (
            O => \N__32799\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__6354\ : LocalMux
    port map (
            O => \N__32790\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__6353\ : LocalMux
    port map (
            O => \N__32783\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__6352\ : LocalMux
    port map (
            O => \N__32770\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__6351\ : LocalMux
    port map (
            O => \N__32753\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__6350\ : CascadeMux
    port map (
            O => \N__32738\,
            I => \N__32735\
        );

    \I__6349\ : InMux
    port map (
            O => \N__32735\,
            I => \N__32732\
        );

    \I__6348\ : LocalMux
    port map (
            O => \N__32732\,
            I => \N__32729\
        );

    \I__6347\ : Span4Mux_h
    port map (
            O => \N__32729\,
            I => \N__32726\
        );

    \I__6346\ : Odrv4
    port map (
            O => \N__32726\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\
        );

    \I__6345\ : InMux
    port map (
            O => \N__32723\,
            I => \N__32717\
        );

    \I__6344\ : InMux
    port map (
            O => \N__32722\,
            I => \N__32698\
        );

    \I__6343\ : InMux
    port map (
            O => \N__32721\,
            I => \N__32698\
        );

    \I__6342\ : InMux
    port map (
            O => \N__32720\,
            I => \N__32695\
        );

    \I__6341\ : LocalMux
    port map (
            O => \N__32717\,
            I => \N__32688\
        );

    \I__6340\ : InMux
    port map (
            O => \N__32716\,
            I => \N__32671\
        );

    \I__6339\ : InMux
    port map (
            O => \N__32715\,
            I => \N__32671\
        );

    \I__6338\ : InMux
    port map (
            O => \N__32714\,
            I => \N__32671\
        );

    \I__6337\ : InMux
    port map (
            O => \N__32713\,
            I => \N__32671\
        );

    \I__6336\ : InMux
    port map (
            O => \N__32712\,
            I => \N__32671\
        );

    \I__6335\ : InMux
    port map (
            O => \N__32711\,
            I => \N__32671\
        );

    \I__6334\ : InMux
    port map (
            O => \N__32710\,
            I => \N__32671\
        );

    \I__6333\ : InMux
    port map (
            O => \N__32709\,
            I => \N__32671\
        );

    \I__6332\ : InMux
    port map (
            O => \N__32708\,
            I => \N__32658\
        );

    \I__6331\ : InMux
    port map (
            O => \N__32707\,
            I => \N__32658\
        );

    \I__6330\ : InMux
    port map (
            O => \N__32706\,
            I => \N__32658\
        );

    \I__6329\ : InMux
    port map (
            O => \N__32705\,
            I => \N__32658\
        );

    \I__6328\ : InMux
    port map (
            O => \N__32704\,
            I => \N__32658\
        );

    \I__6327\ : InMux
    port map (
            O => \N__32703\,
            I => \N__32658\
        );

    \I__6326\ : LocalMux
    port map (
            O => \N__32698\,
            I => \N__32648\
        );

    \I__6325\ : LocalMux
    port map (
            O => \N__32695\,
            I => \N__32648\
        );

    \I__6324\ : InMux
    port map (
            O => \N__32694\,
            I => \N__32639\
        );

    \I__6323\ : InMux
    port map (
            O => \N__32693\,
            I => \N__32639\
        );

    \I__6322\ : InMux
    port map (
            O => \N__32692\,
            I => \N__32639\
        );

    \I__6321\ : InMux
    port map (
            O => \N__32691\,
            I => \N__32639\
        );

    \I__6320\ : Span4Mux_h
    port map (
            O => \N__32688\,
            I => \N__32635\
        );

    \I__6319\ : LocalMux
    port map (
            O => \N__32671\,
            I => \N__32632\
        );

    \I__6318\ : LocalMux
    port map (
            O => \N__32658\,
            I => \N__32629\
        );

    \I__6317\ : InMux
    port map (
            O => \N__32657\,
            I => \N__32618\
        );

    \I__6316\ : InMux
    port map (
            O => \N__32656\,
            I => \N__32618\
        );

    \I__6315\ : InMux
    port map (
            O => \N__32655\,
            I => \N__32618\
        );

    \I__6314\ : InMux
    port map (
            O => \N__32654\,
            I => \N__32618\
        );

    \I__6313\ : InMux
    port map (
            O => \N__32653\,
            I => \N__32618\
        );

    \I__6312\ : Span4Mux_v
    port map (
            O => \N__32648\,
            I => \N__32613\
        );

    \I__6311\ : LocalMux
    port map (
            O => \N__32639\,
            I => \N__32613\
        );

    \I__6310\ : InMux
    port map (
            O => \N__32638\,
            I => \N__32610\
        );

    \I__6309\ : Odrv4
    port map (
            O => \N__32635\,
            I => \current_shift_inst.PI_CTRL.N_79\
        );

    \I__6308\ : Odrv4
    port map (
            O => \N__32632\,
            I => \current_shift_inst.PI_CTRL.N_79\
        );

    \I__6307\ : Odrv4
    port map (
            O => \N__32629\,
            I => \current_shift_inst.PI_CTRL.N_79\
        );

    \I__6306\ : LocalMux
    port map (
            O => \N__32618\,
            I => \current_shift_inst.PI_CTRL.N_79\
        );

    \I__6305\ : Odrv4
    port map (
            O => \N__32613\,
            I => \current_shift_inst.PI_CTRL.N_79\
        );

    \I__6304\ : LocalMux
    port map (
            O => \N__32610\,
            I => \current_shift_inst.PI_CTRL.N_79\
        );

    \I__6303\ : InMux
    port map (
            O => \N__32597\,
            I => \N__32593\
        );

    \I__6302\ : InMux
    port map (
            O => \N__32596\,
            I => \N__32590\
        );

    \I__6301\ : LocalMux
    port map (
            O => \N__32593\,
            I => \N__32585\
        );

    \I__6300\ : LocalMux
    port map (
            O => \N__32590\,
            I => \N__32582\
        );

    \I__6299\ : InMux
    port map (
            O => \N__32589\,
            I => \N__32579\
        );

    \I__6298\ : InMux
    port map (
            O => \N__32588\,
            I => \N__32576\
        );

    \I__6297\ : Span4Mux_h
    port map (
            O => \N__32585\,
            I => \N__32573\
        );

    \I__6296\ : Span12Mux_v
    port map (
            O => \N__32582\,
            I => \N__32566\
        );

    \I__6295\ : LocalMux
    port map (
            O => \N__32579\,
            I => \N__32566\
        );

    \I__6294\ : LocalMux
    port map (
            O => \N__32576\,
            I => \N__32566\
        );

    \I__6293\ : Odrv4
    port map (
            O => \N__32573\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__6292\ : Odrv12
    port map (
            O => \N__32566\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__6291\ : CEMux
    port map (
            O => \N__32561\,
            I => \N__32556\
        );

    \I__6290\ : CEMux
    port map (
            O => \N__32560\,
            I => \N__32544\
        );

    \I__6289\ : CEMux
    port map (
            O => \N__32559\,
            I => \N__32541\
        );

    \I__6288\ : LocalMux
    port map (
            O => \N__32556\,
            I => \N__32537\
        );

    \I__6287\ : CEMux
    port map (
            O => \N__32555\,
            I => \N__32534\
        );

    \I__6286\ : CEMux
    port map (
            O => \N__32554\,
            I => \N__32531\
        );

    \I__6285\ : CEMux
    port map (
            O => \N__32553\,
            I => \N__32527\
        );

    \I__6284\ : CEMux
    port map (
            O => \N__32552\,
            I => \N__32524\
        );

    \I__6283\ : CEMux
    port map (
            O => \N__32551\,
            I => \N__32521\
        );

    \I__6282\ : CEMux
    port map (
            O => \N__32550\,
            I => \N__32518\
        );

    \I__6281\ : CEMux
    port map (
            O => \N__32549\,
            I => \N__32515\
        );

    \I__6280\ : CEMux
    port map (
            O => \N__32548\,
            I => \N__32510\
        );

    \I__6279\ : CEMux
    port map (
            O => \N__32547\,
            I => \N__32507\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__32544\,
            I => \N__32504\
        );

    \I__6277\ : LocalMux
    port map (
            O => \N__32541\,
            I => \N__32501\
        );

    \I__6276\ : CEMux
    port map (
            O => \N__32540\,
            I => \N__32498\
        );

    \I__6275\ : Span4Mux_h
    port map (
            O => \N__32537\,
            I => \N__32492\
        );

    \I__6274\ : LocalMux
    port map (
            O => \N__32534\,
            I => \N__32492\
        );

    \I__6273\ : LocalMux
    port map (
            O => \N__32531\,
            I => \N__32486\
        );

    \I__6272\ : CEMux
    port map (
            O => \N__32530\,
            I => \N__32481\
        );

    \I__6271\ : LocalMux
    port map (
            O => \N__32527\,
            I => \N__32477\
        );

    \I__6270\ : LocalMux
    port map (
            O => \N__32524\,
            I => \N__32470\
        );

    \I__6269\ : LocalMux
    port map (
            O => \N__32521\,
            I => \N__32470\
        );

    \I__6268\ : LocalMux
    port map (
            O => \N__32518\,
            I => \N__32470\
        );

    \I__6267\ : LocalMux
    port map (
            O => \N__32515\,
            I => \N__32467\
        );

    \I__6266\ : CEMux
    port map (
            O => \N__32514\,
            I => \N__32464\
        );

    \I__6265\ : CEMux
    port map (
            O => \N__32513\,
            I => \N__32461\
        );

    \I__6264\ : LocalMux
    port map (
            O => \N__32510\,
            I => \N__32456\
        );

    \I__6263\ : LocalMux
    port map (
            O => \N__32507\,
            I => \N__32456\
        );

    \I__6262\ : Span4Mux_v
    port map (
            O => \N__32504\,
            I => \N__32453\
        );

    \I__6261\ : Span4Mux_v
    port map (
            O => \N__32501\,
            I => \N__32448\
        );

    \I__6260\ : LocalMux
    port map (
            O => \N__32498\,
            I => \N__32448\
        );

    \I__6259\ : CEMux
    port map (
            O => \N__32497\,
            I => \N__32445\
        );

    \I__6258\ : Span4Mux_h
    port map (
            O => \N__32492\,
            I => \N__32442\
        );

    \I__6257\ : CEMux
    port map (
            O => \N__32491\,
            I => \N__32439\
        );

    \I__6256\ : CEMux
    port map (
            O => \N__32490\,
            I => \N__32436\
        );

    \I__6255\ : CEMux
    port map (
            O => \N__32489\,
            I => \N__32433\
        );

    \I__6254\ : Span4Mux_h
    port map (
            O => \N__32486\,
            I => \N__32429\
        );

    \I__6253\ : CEMux
    port map (
            O => \N__32485\,
            I => \N__32426\
        );

    \I__6252\ : CEMux
    port map (
            O => \N__32484\,
            I => \N__32423\
        );

    \I__6251\ : LocalMux
    port map (
            O => \N__32481\,
            I => \N__32420\
        );

    \I__6250\ : CEMux
    port map (
            O => \N__32480\,
            I => \N__32417\
        );

    \I__6249\ : Span4Mux_v
    port map (
            O => \N__32477\,
            I => \N__32414\
        );

    \I__6248\ : Span4Mux_v
    port map (
            O => \N__32470\,
            I => \N__32411\
        );

    \I__6247\ : Span4Mux_h
    port map (
            O => \N__32467\,
            I => \N__32404\
        );

    \I__6246\ : LocalMux
    port map (
            O => \N__32464\,
            I => \N__32404\
        );

    \I__6245\ : LocalMux
    port map (
            O => \N__32461\,
            I => \N__32404\
        );

    \I__6244\ : Span4Mux_v
    port map (
            O => \N__32456\,
            I => \N__32401\
        );

    \I__6243\ : Span4Mux_h
    port map (
            O => \N__32453\,
            I => \N__32396\
        );

    \I__6242\ : Span4Mux_h
    port map (
            O => \N__32448\,
            I => \N__32396\
        );

    \I__6241\ : LocalMux
    port map (
            O => \N__32445\,
            I => \N__32393\
        );

    \I__6240\ : Span4Mux_h
    port map (
            O => \N__32442\,
            I => \N__32384\
        );

    \I__6239\ : LocalMux
    port map (
            O => \N__32439\,
            I => \N__32384\
        );

    \I__6238\ : LocalMux
    port map (
            O => \N__32436\,
            I => \N__32384\
        );

    \I__6237\ : LocalMux
    port map (
            O => \N__32433\,
            I => \N__32384\
        );

    \I__6236\ : CEMux
    port map (
            O => \N__32432\,
            I => \N__32381\
        );

    \I__6235\ : Span4Mux_h
    port map (
            O => \N__32429\,
            I => \N__32376\
        );

    \I__6234\ : LocalMux
    port map (
            O => \N__32426\,
            I => \N__32376\
        );

    \I__6233\ : LocalMux
    port map (
            O => \N__32423\,
            I => \N__32373\
        );

    \I__6232\ : Span12Mux_v
    port map (
            O => \N__32420\,
            I => \N__32370\
        );

    \I__6231\ : LocalMux
    port map (
            O => \N__32417\,
            I => \N__32367\
        );

    \I__6230\ : Span4Mux_h
    port map (
            O => \N__32414\,
            I => \N__32358\
        );

    \I__6229\ : Span4Mux_h
    port map (
            O => \N__32411\,
            I => \N__32358\
        );

    \I__6228\ : Span4Mux_v
    port map (
            O => \N__32404\,
            I => \N__32358\
        );

    \I__6227\ : Span4Mux_s3_h
    port map (
            O => \N__32401\,
            I => \N__32358\
        );

    \I__6226\ : Span4Mux_h
    port map (
            O => \N__32396\,
            I => \N__32349\
        );

    \I__6225\ : Span4Mux_v
    port map (
            O => \N__32393\,
            I => \N__32349\
        );

    \I__6224\ : Span4Mux_v
    port map (
            O => \N__32384\,
            I => \N__32349\
        );

    \I__6223\ : LocalMux
    port map (
            O => \N__32381\,
            I => \N__32349\
        );

    \I__6222\ : Span4Mux_h
    port map (
            O => \N__32376\,
            I => \N__32344\
        );

    \I__6221\ : Span4Mux_h
    port map (
            O => \N__32373\,
            I => \N__32344\
        );

    \I__6220\ : Odrv12
    port map (
            O => \N__32370\,
            I => \N_605_g\
        );

    \I__6219\ : Odrv12
    port map (
            O => \N__32367\,
            I => \N_605_g\
        );

    \I__6218\ : Odrv4
    port map (
            O => \N__32358\,
            I => \N_605_g\
        );

    \I__6217\ : Odrv4
    port map (
            O => \N__32349\,
            I => \N_605_g\
        );

    \I__6216\ : Odrv4
    port map (
            O => \N__32344\,
            I => \N_605_g\
        );

    \I__6215\ : InMux
    port map (
            O => \N__32333\,
            I => \N__32330\
        );

    \I__6214\ : LocalMux
    port map (
            O => \N__32330\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto13_3Z0Z_1\
        );

    \I__6213\ : IoInMux
    port map (
            O => \N__32327\,
            I => \N__32324\
        );

    \I__6212\ : LocalMux
    port map (
            O => \N__32324\,
            I => \N__32321\
        );

    \I__6211\ : Span4Mux_s3_v
    port map (
            O => \N__32321\,
            I => \N__32318\
        );

    \I__6210\ : Span4Mux_h
    port map (
            O => \N__32318\,
            I => \N__32314\
        );

    \I__6209\ : InMux
    port map (
            O => \N__32317\,
            I => \N__32311\
        );

    \I__6208\ : Odrv4
    port map (
            O => \N__32314\,
            I => s1_phy_c
        );

    \I__6207\ : LocalMux
    port map (
            O => \N__32311\,
            I => s1_phy_c
        );

    \I__6206\ : CascadeMux
    port map (
            O => \N__32306\,
            I => \N__32302\
        );

    \I__6205\ : CascadeMux
    port map (
            O => \N__32305\,
            I => \N__32299\
        );

    \I__6204\ : InMux
    port map (
            O => \N__32302\,
            I => \N__32296\
        );

    \I__6203\ : InMux
    port map (
            O => \N__32299\,
            I => \N__32293\
        );

    \I__6202\ : LocalMux
    port map (
            O => \N__32296\,
            I => \N__32289\
        );

    \I__6201\ : LocalMux
    port map (
            O => \N__32293\,
            I => \N__32286\
        );

    \I__6200\ : CascadeMux
    port map (
            O => \N__32292\,
            I => \N__32283\
        );

    \I__6199\ : Span4Mux_v
    port map (
            O => \N__32289\,
            I => \N__32280\
        );

    \I__6198\ : Span4Mux_v
    port map (
            O => \N__32286\,
            I => \N__32277\
        );

    \I__6197\ : InMux
    port map (
            O => \N__32283\,
            I => \N__32274\
        );

    \I__6196\ : Odrv4
    port map (
            O => \N__32280\,
            I => \current_shift_inst.S3_riseZ0\
        );

    \I__6195\ : Odrv4
    port map (
            O => \N__32277\,
            I => \current_shift_inst.S3_riseZ0\
        );

    \I__6194\ : LocalMux
    port map (
            O => \N__32274\,
            I => \current_shift_inst.S3_riseZ0\
        );

    \I__6193\ : InMux
    port map (
            O => \N__32267\,
            I => \N__32264\
        );

    \I__6192\ : LocalMux
    port map (
            O => \N__32264\,
            I => \current_shift_inst.S3_sync_prevZ0\
        );

    \I__6191\ : InMux
    port map (
            O => \N__32261\,
            I => \N__32258\
        );

    \I__6190\ : LocalMux
    port map (
            O => \N__32258\,
            I => \current_shift_inst.S3_syncZ0Z0\
        );

    \I__6189\ : InMux
    port map (
            O => \N__32255\,
            I => \N__32249\
        );

    \I__6188\ : InMux
    port map (
            O => \N__32254\,
            I => \N__32249\
        );

    \I__6187\ : LocalMux
    port map (
            O => \N__32249\,
            I => \current_shift_inst.S3_syncZ0Z1\
        );

    \I__6186\ : InMux
    port map (
            O => \N__32246\,
            I => \N__32240\
        );

    \I__6185\ : InMux
    port map (
            O => \N__32245\,
            I => \N__32240\
        );

    \I__6184\ : LocalMux
    port map (
            O => \N__32240\,
            I => \N__32236\
        );

    \I__6183\ : InMux
    port map (
            O => \N__32239\,
            I => \N__32233\
        );

    \I__6182\ : Span4Mux_h
    port map (
            O => \N__32236\,
            I => \N__32230\
        );

    \I__6181\ : LocalMux
    port map (
            O => \N__32233\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__6180\ : Odrv4
    port map (
            O => \N__32230\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__6179\ : InMux
    port map (
            O => \N__32225\,
            I => \N__32222\
        );

    \I__6178\ : LocalMux
    port map (
            O => \N__32222\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_24\
        );

    \I__6177\ : InMux
    port map (
            O => \N__32219\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\
        );

    \I__6176\ : CascadeMux
    port map (
            O => \N__32216\,
            I => \N__32212\
        );

    \I__6175\ : CascadeMux
    port map (
            O => \N__32215\,
            I => \N__32209\
        );

    \I__6174\ : InMux
    port map (
            O => \N__32212\,
            I => \N__32204\
        );

    \I__6173\ : InMux
    port map (
            O => \N__32209\,
            I => \N__32204\
        );

    \I__6172\ : LocalMux
    port map (
            O => \N__32204\,
            I => \N__32200\
        );

    \I__6171\ : InMux
    port map (
            O => \N__32203\,
            I => \N__32197\
        );

    \I__6170\ : Span4Mux_h
    port map (
            O => \N__32200\,
            I => \N__32194\
        );

    \I__6169\ : LocalMux
    port map (
            O => \N__32197\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__6168\ : Odrv4
    port map (
            O => \N__32194\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__6167\ : InMux
    port map (
            O => \N__32189\,
            I => \N__32186\
        );

    \I__6166\ : LocalMux
    port map (
            O => \N__32186\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_25\
        );

    \I__6165\ : InMux
    port map (
            O => \N__32183\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\
        );

    \I__6164\ : CascadeMux
    port map (
            O => \N__32180\,
            I => \N__32176\
        );

    \I__6163\ : CascadeMux
    port map (
            O => \N__32179\,
            I => \N__32173\
        );

    \I__6162\ : InMux
    port map (
            O => \N__32176\,
            I => \N__32168\
        );

    \I__6161\ : InMux
    port map (
            O => \N__32173\,
            I => \N__32168\
        );

    \I__6160\ : LocalMux
    port map (
            O => \N__32168\,
            I => \N__32164\
        );

    \I__6159\ : InMux
    port map (
            O => \N__32167\,
            I => \N__32161\
        );

    \I__6158\ : Span4Mux_h
    port map (
            O => \N__32164\,
            I => \N__32158\
        );

    \I__6157\ : LocalMux
    port map (
            O => \N__32161\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__6156\ : Odrv4
    port map (
            O => \N__32158\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__6155\ : InMux
    port map (
            O => \N__32153\,
            I => \N__32150\
        );

    \I__6154\ : LocalMux
    port map (
            O => \N__32150\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_26\
        );

    \I__6153\ : InMux
    port map (
            O => \N__32147\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\
        );

    \I__6152\ : InMux
    port map (
            O => \N__32144\,
            I => \N__32140\
        );

    \I__6151\ : InMux
    port map (
            O => \N__32143\,
            I => \N__32137\
        );

    \I__6150\ : LocalMux
    port map (
            O => \N__32140\,
            I => \N__32133\
        );

    \I__6149\ : LocalMux
    port map (
            O => \N__32137\,
            I => \N__32130\
        );

    \I__6148\ : InMux
    port map (
            O => \N__32136\,
            I => \N__32127\
        );

    \I__6147\ : Span4Mux_h
    port map (
            O => \N__32133\,
            I => \N__32124\
        );

    \I__6146\ : Span4Mux_h
    port map (
            O => \N__32130\,
            I => \N__32121\
        );

    \I__6145\ : LocalMux
    port map (
            O => \N__32127\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__6144\ : Odrv4
    port map (
            O => \N__32124\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__6143\ : Odrv4
    port map (
            O => \N__32121\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__6142\ : InMux
    port map (
            O => \N__32114\,
            I => \N__32111\
        );

    \I__6141\ : LocalMux
    port map (
            O => \N__32111\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_27\
        );

    \I__6140\ : InMux
    port map (
            O => \N__32108\,
            I => \bfn_12_22_0_\
        );

    \I__6139\ : InMux
    port map (
            O => \N__32105\,
            I => \N__32101\
        );

    \I__6138\ : InMux
    port map (
            O => \N__32104\,
            I => \N__32098\
        );

    \I__6137\ : LocalMux
    port map (
            O => \N__32101\,
            I => \N__32094\
        );

    \I__6136\ : LocalMux
    port map (
            O => \N__32098\,
            I => \N__32091\
        );

    \I__6135\ : InMux
    port map (
            O => \N__32097\,
            I => \N__32088\
        );

    \I__6134\ : Span4Mux_h
    port map (
            O => \N__32094\,
            I => \N__32085\
        );

    \I__6133\ : Span4Mux_h
    port map (
            O => \N__32091\,
            I => \N__32082\
        );

    \I__6132\ : LocalMux
    port map (
            O => \N__32088\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__6131\ : Odrv4
    port map (
            O => \N__32085\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__6130\ : Odrv4
    port map (
            O => \N__32082\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__6129\ : InMux
    port map (
            O => \N__32075\,
            I => \N__32072\
        );

    \I__6128\ : LocalMux
    port map (
            O => \N__32072\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_28\
        );

    \I__6127\ : InMux
    port map (
            O => \N__32069\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\
        );

    \I__6126\ : InMux
    port map (
            O => \N__32066\,
            I => \N__32063\
        );

    \I__6125\ : LocalMux
    port map (
            O => \N__32063\,
            I => \N__32059\
        );

    \I__6124\ : InMux
    port map (
            O => \N__32062\,
            I => \N__32056\
        );

    \I__6123\ : Span4Mux_h
    port map (
            O => \N__32059\,
            I => \N__32053\
        );

    \I__6122\ : LocalMux
    port map (
            O => \N__32056\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__6121\ : Odrv4
    port map (
            O => \N__32053\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__6120\ : CascadeMux
    port map (
            O => \N__32048\,
            I => \N__32044\
        );

    \I__6119\ : CascadeMux
    port map (
            O => \N__32047\,
            I => \N__32041\
        );

    \I__6118\ : InMux
    port map (
            O => \N__32044\,
            I => \N__32035\
        );

    \I__6117\ : InMux
    port map (
            O => \N__32041\,
            I => \N__32035\
        );

    \I__6116\ : InMux
    port map (
            O => \N__32040\,
            I => \N__32032\
        );

    \I__6115\ : LocalMux
    port map (
            O => \N__32035\,
            I => \N__32029\
        );

    \I__6114\ : LocalMux
    port map (
            O => \N__32032\,
            I => \N__32024\
        );

    \I__6113\ : Span4Mux_v
    port map (
            O => \N__32029\,
            I => \N__32024\
        );

    \I__6112\ : Odrv4
    port map (
            O => \N__32024\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__6111\ : InMux
    port map (
            O => \N__32021\,
            I => \N__32018\
        );

    \I__6110\ : LocalMux
    port map (
            O => \N__32018\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_29\
        );

    \I__6109\ : InMux
    port map (
            O => \N__32015\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\
        );

    \I__6108\ : InMux
    port map (
            O => \N__32012\,
            I => \N__32009\
        );

    \I__6107\ : LocalMux
    port map (
            O => \N__32009\,
            I => \N__32005\
        );

    \I__6106\ : InMux
    port map (
            O => \N__32008\,
            I => \N__32002\
        );

    \I__6105\ : Span4Mux_h
    port map (
            O => \N__32005\,
            I => \N__31999\
        );

    \I__6104\ : LocalMux
    port map (
            O => \N__32002\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__6103\ : Odrv4
    port map (
            O => \N__31999\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__6102\ : CascadeMux
    port map (
            O => \N__31994\,
            I => \N__31990\
        );

    \I__6101\ : CascadeMux
    port map (
            O => \N__31993\,
            I => \N__31987\
        );

    \I__6100\ : InMux
    port map (
            O => \N__31990\,
            I => \N__31981\
        );

    \I__6099\ : InMux
    port map (
            O => \N__31987\,
            I => \N__31981\
        );

    \I__6098\ : InMux
    port map (
            O => \N__31986\,
            I => \N__31978\
        );

    \I__6097\ : LocalMux
    port map (
            O => \N__31981\,
            I => \N__31975\
        );

    \I__6096\ : LocalMux
    port map (
            O => \N__31978\,
            I => \N__31970\
        );

    \I__6095\ : Span4Mux_v
    port map (
            O => \N__31975\,
            I => \N__31970\
        );

    \I__6094\ : Odrv4
    port map (
            O => \N__31970\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__6093\ : InMux
    port map (
            O => \N__31967\,
            I => \N__31964\
        );

    \I__6092\ : LocalMux
    port map (
            O => \N__31964\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_30\
        );

    \I__6091\ : InMux
    port map (
            O => \N__31961\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\
        );

    \I__6090\ : CEMux
    port map (
            O => \N__31958\,
            I => \N__31940\
        );

    \I__6089\ : CEMux
    port map (
            O => \N__31957\,
            I => \N__31940\
        );

    \I__6088\ : CEMux
    port map (
            O => \N__31956\,
            I => \N__31940\
        );

    \I__6087\ : CEMux
    port map (
            O => \N__31955\,
            I => \N__31940\
        );

    \I__6086\ : CEMux
    port map (
            O => \N__31954\,
            I => \N__31940\
        );

    \I__6085\ : CEMux
    port map (
            O => \N__31953\,
            I => \N__31940\
        );

    \I__6084\ : GlobalMux
    port map (
            O => \N__31940\,
            I => \N__31937\
        );

    \I__6083\ : gio2CtrlBuf
    port map (
            O => \N__31937\,
            I => \current_shift_inst.timer_s1.N_187_i_g\
        );

    \I__6082\ : InMux
    port map (
            O => \N__31934\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\
        );

    \I__6081\ : InMux
    port map (
            O => \N__31931\,
            I => \N__31928\
        );

    \I__6080\ : LocalMux
    port map (
            O => \N__31928\,
            I => \N__31924\
        );

    \I__6079\ : InMux
    port map (
            O => \N__31927\,
            I => \N__31921\
        );

    \I__6078\ : Span4Mux_h
    port map (
            O => \N__31924\,
            I => \N__31918\
        );

    \I__6077\ : LocalMux
    port map (
            O => \N__31921\,
            I => \N__31915\
        );

    \I__6076\ : Span4Mux_h
    port map (
            O => \N__31918\,
            I => \N__31910\
        );

    \I__6075\ : Span4Mux_v
    port map (
            O => \N__31915\,
            I => \N__31910\
        );

    \I__6074\ : Odrv4
    port map (
            O => \N__31910\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__6073\ : InMux
    port map (
            O => \N__31907\,
            I => \N__31901\
        );

    \I__6072\ : InMux
    port map (
            O => \N__31906\,
            I => \N__31901\
        );

    \I__6071\ : LocalMux
    port map (
            O => \N__31901\,
            I => \N__31897\
        );

    \I__6070\ : InMux
    port map (
            O => \N__31900\,
            I => \N__31894\
        );

    \I__6069\ : Span4Mux_h
    port map (
            O => \N__31897\,
            I => \N__31891\
        );

    \I__6068\ : LocalMux
    port map (
            O => \N__31894\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__6067\ : Odrv4
    port map (
            O => \N__31891\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__6066\ : InMux
    port map (
            O => \N__31886\,
            I => \N__31883\
        );

    \I__6065\ : LocalMux
    port map (
            O => \N__31883\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_16\
        );

    \I__6064\ : InMux
    port map (
            O => \N__31880\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\
        );

    \I__6063\ : CascadeMux
    port map (
            O => \N__31877\,
            I => \N__31873\
        );

    \I__6062\ : CascadeMux
    port map (
            O => \N__31876\,
            I => \N__31870\
        );

    \I__6061\ : InMux
    port map (
            O => \N__31873\,
            I => \N__31865\
        );

    \I__6060\ : InMux
    port map (
            O => \N__31870\,
            I => \N__31865\
        );

    \I__6059\ : LocalMux
    port map (
            O => \N__31865\,
            I => \N__31861\
        );

    \I__6058\ : InMux
    port map (
            O => \N__31864\,
            I => \N__31858\
        );

    \I__6057\ : Span4Mux_h
    port map (
            O => \N__31861\,
            I => \N__31855\
        );

    \I__6056\ : LocalMux
    port map (
            O => \N__31858\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__6055\ : Odrv4
    port map (
            O => \N__31855\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__6054\ : InMux
    port map (
            O => \N__31850\,
            I => \N__31847\
        );

    \I__6053\ : LocalMux
    port map (
            O => \N__31847\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_17\
        );

    \I__6052\ : InMux
    port map (
            O => \N__31844\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\
        );

    \I__6051\ : CascadeMux
    port map (
            O => \N__31841\,
            I => \N__31837\
        );

    \I__6050\ : CascadeMux
    port map (
            O => \N__31840\,
            I => \N__31834\
        );

    \I__6049\ : InMux
    port map (
            O => \N__31837\,
            I => \N__31829\
        );

    \I__6048\ : InMux
    port map (
            O => \N__31834\,
            I => \N__31829\
        );

    \I__6047\ : LocalMux
    port map (
            O => \N__31829\,
            I => \N__31825\
        );

    \I__6046\ : InMux
    port map (
            O => \N__31828\,
            I => \N__31822\
        );

    \I__6045\ : Span4Mux_h
    port map (
            O => \N__31825\,
            I => \N__31819\
        );

    \I__6044\ : LocalMux
    port map (
            O => \N__31822\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__6043\ : Odrv4
    port map (
            O => \N__31819\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__6042\ : InMux
    port map (
            O => \N__31814\,
            I => \N__31811\
        );

    \I__6041\ : LocalMux
    port map (
            O => \N__31811\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_18\
        );

    \I__6040\ : InMux
    port map (
            O => \N__31808\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\
        );

    \I__6039\ : InMux
    port map (
            O => \N__31805\,
            I => \N__31801\
        );

    \I__6038\ : InMux
    port map (
            O => \N__31804\,
            I => \N__31798\
        );

    \I__6037\ : LocalMux
    port map (
            O => \N__31801\,
            I => \N__31794\
        );

    \I__6036\ : LocalMux
    port map (
            O => \N__31798\,
            I => \N__31791\
        );

    \I__6035\ : InMux
    port map (
            O => \N__31797\,
            I => \N__31788\
        );

    \I__6034\ : Span4Mux_h
    port map (
            O => \N__31794\,
            I => \N__31785\
        );

    \I__6033\ : Span4Mux_h
    port map (
            O => \N__31791\,
            I => \N__31782\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__31788\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__6031\ : Odrv4
    port map (
            O => \N__31785\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__6030\ : Odrv4
    port map (
            O => \N__31782\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__6029\ : InMux
    port map (
            O => \N__31775\,
            I => \N__31772\
        );

    \I__6028\ : LocalMux
    port map (
            O => \N__31772\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_19\
        );

    \I__6027\ : InMux
    port map (
            O => \N__31769\,
            I => \bfn_12_21_0_\
        );

    \I__6026\ : InMux
    port map (
            O => \N__31766\,
            I => \N__31762\
        );

    \I__6025\ : InMux
    port map (
            O => \N__31765\,
            I => \N__31759\
        );

    \I__6024\ : LocalMux
    port map (
            O => \N__31762\,
            I => \N__31755\
        );

    \I__6023\ : LocalMux
    port map (
            O => \N__31759\,
            I => \N__31752\
        );

    \I__6022\ : InMux
    port map (
            O => \N__31758\,
            I => \N__31749\
        );

    \I__6021\ : Span4Mux_h
    port map (
            O => \N__31755\,
            I => \N__31746\
        );

    \I__6020\ : Span4Mux_h
    port map (
            O => \N__31752\,
            I => \N__31743\
        );

    \I__6019\ : LocalMux
    port map (
            O => \N__31749\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__6018\ : Odrv4
    port map (
            O => \N__31746\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__6017\ : Odrv4
    port map (
            O => \N__31743\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__6016\ : InMux
    port map (
            O => \N__31736\,
            I => \N__31733\
        );

    \I__6015\ : LocalMux
    port map (
            O => \N__31733\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_20\
        );

    \I__6014\ : InMux
    port map (
            O => \N__31730\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\
        );

    \I__6013\ : CascadeMux
    port map (
            O => \N__31727\,
            I => \N__31723\
        );

    \I__6012\ : CascadeMux
    port map (
            O => \N__31726\,
            I => \N__31720\
        );

    \I__6011\ : InMux
    port map (
            O => \N__31723\,
            I => \N__31714\
        );

    \I__6010\ : InMux
    port map (
            O => \N__31720\,
            I => \N__31714\
        );

    \I__6009\ : InMux
    port map (
            O => \N__31719\,
            I => \N__31711\
        );

    \I__6008\ : LocalMux
    port map (
            O => \N__31714\,
            I => \N__31708\
        );

    \I__6007\ : LocalMux
    port map (
            O => \N__31711\,
            I => \N__31703\
        );

    \I__6006\ : Span4Mux_v
    port map (
            O => \N__31708\,
            I => \N__31703\
        );

    \I__6005\ : Odrv4
    port map (
            O => \N__31703\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__6004\ : InMux
    port map (
            O => \N__31700\,
            I => \N__31697\
        );

    \I__6003\ : LocalMux
    port map (
            O => \N__31697\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_21\
        );

    \I__6002\ : InMux
    port map (
            O => \N__31694\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\
        );

    \I__6001\ : CascadeMux
    port map (
            O => \N__31691\,
            I => \N__31687\
        );

    \I__6000\ : CascadeMux
    port map (
            O => \N__31690\,
            I => \N__31684\
        );

    \I__5999\ : InMux
    port map (
            O => \N__31687\,
            I => \N__31678\
        );

    \I__5998\ : InMux
    port map (
            O => \N__31684\,
            I => \N__31678\
        );

    \I__5997\ : InMux
    port map (
            O => \N__31683\,
            I => \N__31675\
        );

    \I__5996\ : LocalMux
    port map (
            O => \N__31678\,
            I => \N__31672\
        );

    \I__5995\ : LocalMux
    port map (
            O => \N__31675\,
            I => \N__31667\
        );

    \I__5994\ : Span4Mux_v
    port map (
            O => \N__31672\,
            I => \N__31667\
        );

    \I__5993\ : Odrv4
    port map (
            O => \N__31667\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__5992\ : InMux
    port map (
            O => \N__31664\,
            I => \N__31661\
        );

    \I__5991\ : LocalMux
    port map (
            O => \N__31661\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_22\
        );

    \I__5990\ : InMux
    port map (
            O => \N__31658\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\
        );

    \I__5989\ : InMux
    port map (
            O => \N__31655\,
            I => \N__31649\
        );

    \I__5988\ : InMux
    port map (
            O => \N__31654\,
            I => \N__31649\
        );

    \I__5987\ : LocalMux
    port map (
            O => \N__31649\,
            I => \N__31645\
        );

    \I__5986\ : InMux
    port map (
            O => \N__31648\,
            I => \N__31642\
        );

    \I__5985\ : Span4Mux_h
    port map (
            O => \N__31645\,
            I => \N__31639\
        );

    \I__5984\ : LocalMux
    port map (
            O => \N__31642\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__5983\ : Odrv4
    port map (
            O => \N__31639\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__5982\ : InMux
    port map (
            O => \N__31634\,
            I => \N__31631\
        );

    \I__5981\ : LocalMux
    port map (
            O => \N__31631\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_23\
        );

    \I__5980\ : InMux
    port map (
            O => \N__31628\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\
        );

    \I__5979\ : InMux
    port map (
            O => \N__31625\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\
        );

    \I__5978\ : InMux
    port map (
            O => \N__31622\,
            I => \N__31616\
        );

    \I__5977\ : InMux
    port map (
            O => \N__31621\,
            I => \N__31616\
        );

    \I__5976\ : LocalMux
    port map (
            O => \N__31616\,
            I => \N__31612\
        );

    \I__5975\ : InMux
    port map (
            O => \N__31615\,
            I => \N__31609\
        );

    \I__5974\ : Span4Mux_h
    port map (
            O => \N__31612\,
            I => \N__31606\
        );

    \I__5973\ : LocalMux
    port map (
            O => \N__31609\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__5972\ : Odrv4
    port map (
            O => \N__31606\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__5971\ : InMux
    port map (
            O => \N__31601\,
            I => \N__31598\
        );

    \I__5970\ : LocalMux
    port map (
            O => \N__31598\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_9\
        );

    \I__5969\ : InMux
    port map (
            O => \N__31595\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\
        );

    \I__5968\ : InMux
    port map (
            O => \N__31592\,
            I => \N__31586\
        );

    \I__5967\ : InMux
    port map (
            O => \N__31591\,
            I => \N__31586\
        );

    \I__5966\ : LocalMux
    port map (
            O => \N__31586\,
            I => \N__31582\
        );

    \I__5965\ : InMux
    port map (
            O => \N__31585\,
            I => \N__31579\
        );

    \I__5964\ : Span4Mux_h
    port map (
            O => \N__31582\,
            I => \N__31576\
        );

    \I__5963\ : LocalMux
    port map (
            O => \N__31579\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__5962\ : Odrv4
    port map (
            O => \N__31576\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__5961\ : InMux
    port map (
            O => \N__31571\,
            I => \N__31568\
        );

    \I__5960\ : LocalMux
    port map (
            O => \N__31568\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_10\
        );

    \I__5959\ : InMux
    port map (
            O => \N__31565\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\
        );

    \I__5958\ : CascadeMux
    port map (
            O => \N__31562\,
            I => \N__31558\
        );

    \I__5957\ : InMux
    port map (
            O => \N__31561\,
            I => \N__31555\
        );

    \I__5956\ : InMux
    port map (
            O => \N__31558\,
            I => \N__31552\
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__31555\,
            I => \N__31548\
        );

    \I__5954\ : LocalMux
    port map (
            O => \N__31552\,
            I => \N__31545\
        );

    \I__5953\ : InMux
    port map (
            O => \N__31551\,
            I => \N__31542\
        );

    \I__5952\ : Span4Mux_h
    port map (
            O => \N__31548\,
            I => \N__31539\
        );

    \I__5951\ : Span4Mux_h
    port map (
            O => \N__31545\,
            I => \N__31536\
        );

    \I__5950\ : LocalMux
    port map (
            O => \N__31542\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__5949\ : Odrv4
    port map (
            O => \N__31539\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__5948\ : Odrv4
    port map (
            O => \N__31536\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__5947\ : InMux
    port map (
            O => \N__31529\,
            I => \N__31526\
        );

    \I__5946\ : LocalMux
    port map (
            O => \N__31526\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_11\
        );

    \I__5945\ : InMux
    port map (
            O => \N__31523\,
            I => \bfn_12_20_0_\
        );

    \I__5944\ : CascadeMux
    port map (
            O => \N__31520\,
            I => \N__31516\
        );

    \I__5943\ : InMux
    port map (
            O => \N__31519\,
            I => \N__31513\
        );

    \I__5942\ : InMux
    port map (
            O => \N__31516\,
            I => \N__31510\
        );

    \I__5941\ : LocalMux
    port map (
            O => \N__31513\,
            I => \N__31506\
        );

    \I__5940\ : LocalMux
    port map (
            O => \N__31510\,
            I => \N__31503\
        );

    \I__5939\ : InMux
    port map (
            O => \N__31509\,
            I => \N__31500\
        );

    \I__5938\ : Span4Mux_h
    port map (
            O => \N__31506\,
            I => \N__31497\
        );

    \I__5937\ : Span4Mux_h
    port map (
            O => \N__31503\,
            I => \N__31494\
        );

    \I__5936\ : LocalMux
    port map (
            O => \N__31500\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__5935\ : Odrv4
    port map (
            O => \N__31497\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__5934\ : Odrv4
    port map (
            O => \N__31494\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__5933\ : InMux
    port map (
            O => \N__31487\,
            I => \N__31484\
        );

    \I__5932\ : LocalMux
    port map (
            O => \N__31484\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_12\
        );

    \I__5931\ : InMux
    port map (
            O => \N__31481\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\
        );

    \I__5930\ : CascadeMux
    port map (
            O => \N__31478\,
            I => \N__31474\
        );

    \I__5929\ : CascadeMux
    port map (
            O => \N__31477\,
            I => \N__31471\
        );

    \I__5928\ : InMux
    port map (
            O => \N__31474\,
            I => \N__31465\
        );

    \I__5927\ : InMux
    port map (
            O => \N__31471\,
            I => \N__31465\
        );

    \I__5926\ : InMux
    port map (
            O => \N__31470\,
            I => \N__31462\
        );

    \I__5925\ : LocalMux
    port map (
            O => \N__31465\,
            I => \N__31459\
        );

    \I__5924\ : LocalMux
    port map (
            O => \N__31462\,
            I => \N__31454\
        );

    \I__5923\ : Span4Mux_v
    port map (
            O => \N__31459\,
            I => \N__31454\
        );

    \I__5922\ : Odrv4
    port map (
            O => \N__31454\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__5921\ : InMux
    port map (
            O => \N__31451\,
            I => \N__31448\
        );

    \I__5920\ : LocalMux
    port map (
            O => \N__31448\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_13\
        );

    \I__5919\ : InMux
    port map (
            O => \N__31445\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\
        );

    \I__5918\ : CascadeMux
    port map (
            O => \N__31442\,
            I => \N__31438\
        );

    \I__5917\ : CascadeMux
    port map (
            O => \N__31441\,
            I => \N__31435\
        );

    \I__5916\ : InMux
    port map (
            O => \N__31438\,
            I => \N__31429\
        );

    \I__5915\ : InMux
    port map (
            O => \N__31435\,
            I => \N__31429\
        );

    \I__5914\ : InMux
    port map (
            O => \N__31434\,
            I => \N__31426\
        );

    \I__5913\ : LocalMux
    port map (
            O => \N__31429\,
            I => \N__31423\
        );

    \I__5912\ : LocalMux
    port map (
            O => \N__31426\,
            I => \N__31418\
        );

    \I__5911\ : Span4Mux_v
    port map (
            O => \N__31423\,
            I => \N__31418\
        );

    \I__5910\ : Odrv4
    port map (
            O => \N__31418\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__5909\ : InMux
    port map (
            O => \N__31415\,
            I => \N__31412\
        );

    \I__5908\ : LocalMux
    port map (
            O => \N__31412\,
            I => \N__31409\
        );

    \I__5907\ : Odrv4
    port map (
            O => \N__31409\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_14\
        );

    \I__5906\ : InMux
    port map (
            O => \N__31406\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\
        );

    \I__5905\ : InMux
    port map (
            O => \N__31403\,
            I => \N__31397\
        );

    \I__5904\ : InMux
    port map (
            O => \N__31402\,
            I => \N__31397\
        );

    \I__5903\ : LocalMux
    port map (
            O => \N__31397\,
            I => \N__31393\
        );

    \I__5902\ : InMux
    port map (
            O => \N__31396\,
            I => \N__31390\
        );

    \I__5901\ : Span4Mux_h
    port map (
            O => \N__31393\,
            I => \N__31387\
        );

    \I__5900\ : LocalMux
    port map (
            O => \N__31390\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__5899\ : Odrv4
    port map (
            O => \N__31387\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__5898\ : InMux
    port map (
            O => \N__31382\,
            I => \N__31379\
        );

    \I__5897\ : LocalMux
    port map (
            O => \N__31379\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_15\
        );

    \I__5896\ : InMux
    port map (
            O => \N__31376\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\
        );

    \I__5895\ : InMux
    port map (
            O => \N__31373\,
            I => \N__31367\
        );

    \I__5894\ : InMux
    port map (
            O => \N__31372\,
            I => \N__31367\
        );

    \I__5893\ : LocalMux
    port map (
            O => \N__31367\,
            I => \N__31363\
        );

    \I__5892\ : InMux
    port map (
            O => \N__31366\,
            I => \N__31360\
        );

    \I__5891\ : Span4Mux_h
    port map (
            O => \N__31363\,
            I => \N__31357\
        );

    \I__5890\ : LocalMux
    port map (
            O => \N__31360\,
            I => \N__31354\
        );

    \I__5889\ : Span4Mux_v
    port map (
            O => \N__31357\,
            I => \N__31350\
        );

    \I__5888\ : Span4Mux_v
    port map (
            O => \N__31354\,
            I => \N__31347\
        );

    \I__5887\ : InMux
    port map (
            O => \N__31353\,
            I => \N__31344\
        );

    \I__5886\ : Odrv4
    port map (
            O => \N__31350\,
            I => \current_shift_inst.elapsed_time_ns_phase_26\
        );

    \I__5885\ : Odrv4
    port map (
            O => \N__31347\,
            I => \current_shift_inst.elapsed_time_ns_phase_26\
        );

    \I__5884\ : LocalMux
    port map (
            O => \N__31344\,
            I => \current_shift_inst.elapsed_time_ns_phase_26\
        );

    \I__5883\ : CascadeMux
    port map (
            O => \N__31337\,
            I => \N__31333\
        );

    \I__5882\ : InMux
    port map (
            O => \N__31336\,
            I => \N__31329\
        );

    \I__5881\ : InMux
    port map (
            O => \N__31333\,
            I => \N__31324\
        );

    \I__5880\ : InMux
    port map (
            O => \N__31332\,
            I => \N__31324\
        );

    \I__5879\ : LocalMux
    port map (
            O => \N__31329\,
            I => \N__31320\
        );

    \I__5878\ : LocalMux
    port map (
            O => \N__31324\,
            I => \N__31317\
        );

    \I__5877\ : CascadeMux
    port map (
            O => \N__31323\,
            I => \N__31314\
        );

    \I__5876\ : Span4Mux_h
    port map (
            O => \N__31320\,
            I => \N__31311\
        );

    \I__5875\ : Span4Mux_h
    port map (
            O => \N__31317\,
            I => \N__31308\
        );

    \I__5874\ : InMux
    port map (
            O => \N__31314\,
            I => \N__31305\
        );

    \I__5873\ : Odrv4
    port map (
            O => \N__31311\,
            I => \current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0\
        );

    \I__5872\ : Odrv4
    port map (
            O => \N__31308\,
            I => \current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0\
        );

    \I__5871\ : LocalMux
    port map (
            O => \N__31305\,
            I => \current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0\
        );

    \I__5870\ : CascadeMux
    port map (
            O => \N__31298\,
            I => \N__31295\
        );

    \I__5869\ : InMux
    port map (
            O => \N__31295\,
            I => \N__31292\
        );

    \I__5868\ : LocalMux
    port map (
            O => \N__31292\,
            I => \N__31289\
        );

    \I__5867\ : Span4Mux_h
    port map (
            O => \N__31289\,
            I => \N__31286\
        );

    \I__5866\ : Odrv4
    port map (
            O => \N__31286\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI7K6K_26\
        );

    \I__5865\ : InMux
    port map (
            O => \N__31283\,
            I => \N__31279\
        );

    \I__5864\ : InMux
    port map (
            O => \N__31282\,
            I => \N__31276\
        );

    \I__5863\ : LocalMux
    port map (
            O => \N__31279\,
            I => \N__31272\
        );

    \I__5862\ : LocalMux
    port map (
            O => \N__31276\,
            I => \N__31268\
        );

    \I__5861\ : CascadeMux
    port map (
            O => \N__31275\,
            I => \N__31265\
        );

    \I__5860\ : Span4Mux_h
    port map (
            O => \N__31272\,
            I => \N__31262\
        );

    \I__5859\ : InMux
    port map (
            O => \N__31271\,
            I => \N__31259\
        );

    \I__5858\ : Span4Mux_v
    port map (
            O => \N__31268\,
            I => \N__31256\
        );

    \I__5857\ : InMux
    port map (
            O => \N__31265\,
            I => \N__31253\
        );

    \I__5856\ : Span4Mux_h
    port map (
            O => \N__31262\,
            I => \N__31250\
        );

    \I__5855\ : LocalMux
    port map (
            O => \N__31259\,
            I => \N__31247\
        );

    \I__5854\ : Span4Mux_h
    port map (
            O => \N__31256\,
            I => \N__31242\
        );

    \I__5853\ : LocalMux
    port map (
            O => \N__31253\,
            I => \N__31242\
        );

    \I__5852\ : Odrv4
    port map (
            O => \N__31250\,
            I => \current_shift_inst.elapsed_time_ns_phase_24\
        );

    \I__5851\ : Odrv12
    port map (
            O => \N__31247\,
            I => \current_shift_inst.elapsed_time_ns_phase_24\
        );

    \I__5850\ : Odrv4
    port map (
            O => \N__31242\,
            I => \current_shift_inst.elapsed_time_ns_phase_24\
        );

    \I__5849\ : CascadeMux
    port map (
            O => \N__31235\,
            I => \N__31232\
        );

    \I__5848\ : InMux
    port map (
            O => \N__31232\,
            I => \N__31227\
        );

    \I__5847\ : InMux
    port map (
            O => \N__31231\,
            I => \N__31224\
        );

    \I__5846\ : InMux
    port map (
            O => \N__31230\,
            I => \N__31221\
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__31227\,
            I => \N__31215\
        );

    \I__5844\ : LocalMux
    port map (
            O => \N__31224\,
            I => \N__31215\
        );

    \I__5843\ : LocalMux
    port map (
            O => \N__31221\,
            I => \N__31212\
        );

    \I__5842\ : CascadeMux
    port map (
            O => \N__31220\,
            I => \N__31209\
        );

    \I__5841\ : Span4Mux_h
    port map (
            O => \N__31215\,
            I => \N__31206\
        );

    \I__5840\ : Span4Mux_h
    port map (
            O => \N__31212\,
            I => \N__31203\
        );

    \I__5839\ : InMux
    port map (
            O => \N__31209\,
            I => \N__31200\
        );

    \I__5838\ : Odrv4
    port map (
            O => \N__31206\,
            I => \current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0\
        );

    \I__5837\ : Odrv4
    port map (
            O => \N__31203\,
            I => \current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0\
        );

    \I__5836\ : LocalMux
    port map (
            O => \N__31200\,
            I => \current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0\
        );

    \I__5835\ : CascadeMux
    port map (
            O => \N__31193\,
            I => \N__31190\
        );

    \I__5834\ : InMux
    port map (
            O => \N__31190\,
            I => \N__31185\
        );

    \I__5833\ : InMux
    port map (
            O => \N__31189\,
            I => \N__31182\
        );

    \I__5832\ : InMux
    port map (
            O => \N__31188\,
            I => \N__31179\
        );

    \I__5831\ : LocalMux
    port map (
            O => \N__31185\,
            I => \N__31175\
        );

    \I__5830\ : LocalMux
    port map (
            O => \N__31182\,
            I => \N__31172\
        );

    \I__5829\ : LocalMux
    port map (
            O => \N__31179\,
            I => \N__31169\
        );

    \I__5828\ : CascadeMux
    port map (
            O => \N__31178\,
            I => \N__31166\
        );

    \I__5827\ : Span4Mux_v
    port map (
            O => \N__31175\,
            I => \N__31163\
        );

    \I__5826\ : Span4Mux_h
    port map (
            O => \N__31172\,
            I => \N__31160\
        );

    \I__5825\ : Span4Mux_h
    port map (
            O => \N__31169\,
            I => \N__31157\
        );

    \I__5824\ : InMux
    port map (
            O => \N__31166\,
            I => \N__31154\
        );

    \I__5823\ : Odrv4
    port map (
            O => \N__31163\,
            I => \current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0\
        );

    \I__5822\ : Odrv4
    port map (
            O => \N__31160\,
            I => \current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0\
        );

    \I__5821\ : Odrv4
    port map (
            O => \N__31157\,
            I => \current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0\
        );

    \I__5820\ : LocalMux
    port map (
            O => \N__31154\,
            I => \current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0\
        );

    \I__5819\ : InMux
    port map (
            O => \N__31145\,
            I => \N__31142\
        );

    \I__5818\ : LocalMux
    port map (
            O => \N__31142\,
            I => \N__31137\
        );

    \I__5817\ : InMux
    port map (
            O => \N__31141\,
            I => \N__31132\
        );

    \I__5816\ : InMux
    port map (
            O => \N__31140\,
            I => \N__31132\
        );

    \I__5815\ : Span4Mux_h
    port map (
            O => \N__31137\,
            I => \N__31129\
        );

    \I__5814\ : LocalMux
    port map (
            O => \N__31132\,
            I => \N__31125\
        );

    \I__5813\ : Span4Mux_h
    port map (
            O => \N__31129\,
            I => \N__31122\
        );

    \I__5812\ : InMux
    port map (
            O => \N__31128\,
            I => \N__31119\
        );

    \I__5811\ : Odrv12
    port map (
            O => \N__31125\,
            I => \current_shift_inst.elapsed_time_ns_phase_25\
        );

    \I__5810\ : Odrv4
    port map (
            O => \N__31122\,
            I => \current_shift_inst.elapsed_time_ns_phase_25\
        );

    \I__5809\ : LocalMux
    port map (
            O => \N__31119\,
            I => \current_shift_inst.elapsed_time_ns_phase_25\
        );

    \I__5808\ : InMux
    port map (
            O => \N__31112\,
            I => \N__31109\
        );

    \I__5807\ : LocalMux
    port map (
            O => \N__31109\,
            I => \N__31106\
        );

    \I__5806\ : Span4Mux_h
    port map (
            O => \N__31106\,
            I => \N__31103\
        );

    \I__5805\ : Odrv4
    port map (
            O => \N__31103\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5S981_24\
        );

    \I__5804\ : CascadeMux
    port map (
            O => \N__31100\,
            I => \N__31096\
        );

    \I__5803\ : InMux
    port map (
            O => \N__31099\,
            I => \N__31093\
        );

    \I__5802\ : InMux
    port map (
            O => \N__31096\,
            I => \N__31090\
        );

    \I__5801\ : LocalMux
    port map (
            O => \N__31093\,
            I => \N__31087\
        );

    \I__5800\ : LocalMux
    port map (
            O => \N__31090\,
            I => \N__31083\
        );

    \I__5799\ : Span4Mux_v
    port map (
            O => \N__31087\,
            I => \N__31080\
        );

    \I__5798\ : InMux
    port map (
            O => \N__31086\,
            I => \N__31077\
        );

    \I__5797\ : Span4Mux_h
    port map (
            O => \N__31083\,
            I => \N__31074\
        );

    \I__5796\ : Odrv4
    port map (
            O => \N__31080\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__5795\ : LocalMux
    port map (
            O => \N__31077\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__5794\ : Odrv4
    port map (
            O => \N__31074\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__5793\ : InMux
    port map (
            O => \N__31067\,
            I => \N__31064\
        );

    \I__5792\ : LocalMux
    port map (
            O => \N__31064\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_3\
        );

    \I__5791\ : CascadeMux
    port map (
            O => \N__31061\,
            I => \N__31057\
        );

    \I__5790\ : InMux
    port map (
            O => \N__31060\,
            I => \N__31054\
        );

    \I__5789\ : InMux
    port map (
            O => \N__31057\,
            I => \N__31051\
        );

    \I__5788\ : LocalMux
    port map (
            O => \N__31054\,
            I => \N__31048\
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__31051\,
            I => \N__31044\
        );

    \I__5786\ : Span4Mux_v
    port map (
            O => \N__31048\,
            I => \N__31041\
        );

    \I__5785\ : InMux
    port map (
            O => \N__31047\,
            I => \N__31038\
        );

    \I__5784\ : Span4Mux_h
    port map (
            O => \N__31044\,
            I => \N__31035\
        );

    \I__5783\ : Odrv4
    port map (
            O => \N__31041\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__5782\ : LocalMux
    port map (
            O => \N__31038\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__5781\ : Odrv4
    port map (
            O => \N__31035\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__5780\ : InMux
    port map (
            O => \N__31028\,
            I => \N__31025\
        );

    \I__5779\ : LocalMux
    port map (
            O => \N__31025\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_4\
        );

    \I__5778\ : InMux
    port map (
            O => \N__31022\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\
        );

    \I__5777\ : InMux
    port map (
            O => \N__31019\,
            I => \N__31012\
        );

    \I__5776\ : InMux
    port map (
            O => \N__31018\,
            I => \N__31012\
        );

    \I__5775\ : InMux
    port map (
            O => \N__31017\,
            I => \N__31009\
        );

    \I__5774\ : LocalMux
    port map (
            O => \N__31012\,
            I => \N__31006\
        );

    \I__5773\ : LocalMux
    port map (
            O => \N__31009\,
            I => \N__31001\
        );

    \I__5772\ : Span4Mux_v
    port map (
            O => \N__31006\,
            I => \N__31001\
        );

    \I__5771\ : Odrv4
    port map (
            O => \N__31001\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__5770\ : InMux
    port map (
            O => \N__30998\,
            I => \N__30995\
        );

    \I__5769\ : LocalMux
    port map (
            O => \N__30995\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_5\
        );

    \I__5768\ : InMux
    port map (
            O => \N__30992\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\
        );

    \I__5767\ : InMux
    port map (
            O => \N__30989\,
            I => \N__30982\
        );

    \I__5766\ : InMux
    port map (
            O => \N__30988\,
            I => \N__30982\
        );

    \I__5765\ : InMux
    port map (
            O => \N__30987\,
            I => \N__30979\
        );

    \I__5764\ : LocalMux
    port map (
            O => \N__30982\,
            I => \N__30976\
        );

    \I__5763\ : LocalMux
    port map (
            O => \N__30979\,
            I => \N__30971\
        );

    \I__5762\ : Span4Mux_v
    port map (
            O => \N__30976\,
            I => \N__30971\
        );

    \I__5761\ : Odrv4
    port map (
            O => \N__30971\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__5760\ : InMux
    port map (
            O => \N__30968\,
            I => \N__30965\
        );

    \I__5759\ : LocalMux
    port map (
            O => \N__30965\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_6\
        );

    \I__5758\ : InMux
    port map (
            O => \N__30962\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\
        );

    \I__5757\ : CascadeMux
    port map (
            O => \N__30959\,
            I => \N__30955\
        );

    \I__5756\ : CascadeMux
    port map (
            O => \N__30958\,
            I => \N__30952\
        );

    \I__5755\ : InMux
    port map (
            O => \N__30955\,
            I => \N__30947\
        );

    \I__5754\ : InMux
    port map (
            O => \N__30952\,
            I => \N__30947\
        );

    \I__5753\ : LocalMux
    port map (
            O => \N__30947\,
            I => \N__30943\
        );

    \I__5752\ : InMux
    port map (
            O => \N__30946\,
            I => \N__30940\
        );

    \I__5751\ : Span4Mux_h
    port map (
            O => \N__30943\,
            I => \N__30937\
        );

    \I__5750\ : LocalMux
    port map (
            O => \N__30940\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__5749\ : Odrv4
    port map (
            O => \N__30937\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__5748\ : InMux
    port map (
            O => \N__30932\,
            I => \N__30929\
        );

    \I__5747\ : LocalMux
    port map (
            O => \N__30929\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_7\
        );

    \I__5746\ : InMux
    port map (
            O => \N__30926\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\
        );

    \I__5745\ : CascadeMux
    port map (
            O => \N__30923\,
            I => \N__30919\
        );

    \I__5744\ : CascadeMux
    port map (
            O => \N__30922\,
            I => \N__30916\
        );

    \I__5743\ : InMux
    port map (
            O => \N__30919\,
            I => \N__30911\
        );

    \I__5742\ : InMux
    port map (
            O => \N__30916\,
            I => \N__30911\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__30911\,
            I => \N__30907\
        );

    \I__5740\ : InMux
    port map (
            O => \N__30910\,
            I => \N__30904\
        );

    \I__5739\ : Span4Mux_h
    port map (
            O => \N__30907\,
            I => \N__30901\
        );

    \I__5738\ : LocalMux
    port map (
            O => \N__30904\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__5737\ : Odrv4
    port map (
            O => \N__30901\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__5736\ : InMux
    port map (
            O => \N__30896\,
            I => \N__30893\
        );

    \I__5735\ : LocalMux
    port map (
            O => \N__30893\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_8\
        );

    \I__5734\ : InMux
    port map (
            O => \N__30890\,
            I => \N__30887\
        );

    \I__5733\ : LocalMux
    port map (
            O => \N__30887\,
            I => \N__30882\
        );

    \I__5732\ : InMux
    port map (
            O => \N__30886\,
            I => \N__30879\
        );

    \I__5731\ : InMux
    port map (
            O => \N__30885\,
            I => \N__30876\
        );

    \I__5730\ : Span4Mux_v
    port map (
            O => \N__30882\,
            I => \N__30871\
        );

    \I__5729\ : LocalMux
    port map (
            O => \N__30879\,
            I => \N__30871\
        );

    \I__5728\ : LocalMux
    port map (
            O => \N__30876\,
            I => \N__30868\
        );

    \I__5727\ : Span4Mux_h
    port map (
            O => \N__30871\,
            I => \N__30864\
        );

    \I__5726\ : Span4Mux_h
    port map (
            O => \N__30868\,
            I => \N__30861\
        );

    \I__5725\ : InMux
    port map (
            O => \N__30867\,
            I => \N__30858\
        );

    \I__5724\ : Span4Mux_v
    port map (
            O => \N__30864\,
            I => \N__30855\
        );

    \I__5723\ : Span4Mux_h
    port map (
            O => \N__30861\,
            I => \N__30850\
        );

    \I__5722\ : LocalMux
    port map (
            O => \N__30858\,
            I => \N__30850\
        );

    \I__5721\ : Odrv4
    port map (
            O => \N__30855\,
            I => \current_shift_inst.elapsed_time_ns_phase_11\
        );

    \I__5720\ : Odrv4
    port map (
            O => \N__30850\,
            I => \current_shift_inst.elapsed_time_ns_phase_11\
        );

    \I__5719\ : InMux
    port map (
            O => \N__30845\,
            I => \N__30840\
        );

    \I__5718\ : InMux
    port map (
            O => \N__30844\,
            I => \N__30837\
        );

    \I__5717\ : InMux
    port map (
            O => \N__30843\,
            I => \N__30834\
        );

    \I__5716\ : LocalMux
    port map (
            O => \N__30840\,
            I => \N__30831\
        );

    \I__5715\ : LocalMux
    port map (
            O => \N__30837\,
            I => \N__30828\
        );

    \I__5714\ : LocalMux
    port map (
            O => \N__30834\,
            I => \N__30824\
        );

    \I__5713\ : Span4Mux_h
    port map (
            O => \N__30831\,
            I => \N__30819\
        );

    \I__5712\ : Span4Mux_h
    port map (
            O => \N__30828\,
            I => \N__30819\
        );

    \I__5711\ : InMux
    port map (
            O => \N__30827\,
            I => \N__30816\
        );

    \I__5710\ : Odrv12
    port map (
            O => \N__30824\,
            I => \current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0\
        );

    \I__5709\ : Odrv4
    port map (
            O => \N__30819\,
            I => \current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0\
        );

    \I__5708\ : LocalMux
    port map (
            O => \N__30816\,
            I => \current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0\
        );

    \I__5707\ : CascadeMux
    port map (
            O => \N__30809\,
            I => \N__30806\
        );

    \I__5706\ : InMux
    port map (
            O => \N__30806\,
            I => \N__30802\
        );

    \I__5705\ : InMux
    port map (
            O => \N__30805\,
            I => \N__30798\
        );

    \I__5704\ : LocalMux
    port map (
            O => \N__30802\,
            I => \N__30794\
        );

    \I__5703\ : InMux
    port map (
            O => \N__30801\,
            I => \N__30791\
        );

    \I__5702\ : LocalMux
    port map (
            O => \N__30798\,
            I => \N__30788\
        );

    \I__5701\ : CascadeMux
    port map (
            O => \N__30797\,
            I => \N__30785\
        );

    \I__5700\ : Span4Mux_h
    port map (
            O => \N__30794\,
            I => \N__30782\
        );

    \I__5699\ : LocalMux
    port map (
            O => \N__30791\,
            I => \N__30779\
        );

    \I__5698\ : Span4Mux_h
    port map (
            O => \N__30788\,
            I => \N__30776\
        );

    \I__5697\ : InMux
    port map (
            O => \N__30785\,
            I => \N__30773\
        );

    \I__5696\ : Odrv4
    port map (
            O => \N__30782\,
            I => \current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0\
        );

    \I__5695\ : Odrv12
    port map (
            O => \N__30779\,
            I => \current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0\
        );

    \I__5694\ : Odrv4
    port map (
            O => \N__30776\,
            I => \current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0\
        );

    \I__5693\ : LocalMux
    port map (
            O => \N__30773\,
            I => \current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0\
        );

    \I__5692\ : InMux
    port map (
            O => \N__30764\,
            I => \N__30759\
        );

    \I__5691\ : InMux
    port map (
            O => \N__30763\,
            I => \N__30756\
        );

    \I__5690\ : InMux
    port map (
            O => \N__30762\,
            I => \N__30753\
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__30759\,
            I => \N__30750\
        );

    \I__5688\ : LocalMux
    port map (
            O => \N__30756\,
            I => \N__30747\
        );

    \I__5687\ : LocalMux
    port map (
            O => \N__30753\,
            I => \N__30741\
        );

    \I__5686\ : Span4Mux_h
    port map (
            O => \N__30750\,
            I => \N__30741\
        );

    \I__5685\ : Span4Mux_h
    port map (
            O => \N__30747\,
            I => \N__30738\
        );

    \I__5684\ : InMux
    port map (
            O => \N__30746\,
            I => \N__30735\
        );

    \I__5683\ : Span4Mux_v
    port map (
            O => \N__30741\,
            I => \N__30728\
        );

    \I__5682\ : Span4Mux_h
    port map (
            O => \N__30738\,
            I => \N__30728\
        );

    \I__5681\ : LocalMux
    port map (
            O => \N__30735\,
            I => \N__30728\
        );

    \I__5680\ : Odrv4
    port map (
            O => \N__30728\,
            I => \current_shift_inst.elapsed_time_ns_phase_12\
        );

    \I__5679\ : InMux
    port map (
            O => \N__30725\,
            I => \N__30722\
        );

    \I__5678\ : LocalMux
    port map (
            O => \N__30722\,
            I => \N__30719\
        );

    \I__5677\ : Span4Mux_h
    port map (
            O => \N__30719\,
            I => \N__30716\
        );

    \I__5676\ : Odrv4
    port map (
            O => \N__30716\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIDLO51_11\
        );

    \I__5675\ : CascadeMux
    port map (
            O => \N__30713\,
            I => \N__30710\
        );

    \I__5674\ : InMux
    port map (
            O => \N__30710\,
            I => \N__30707\
        );

    \I__5673\ : LocalMux
    port map (
            O => \N__30707\,
            I => \N__30704\
        );

    \I__5672\ : Span4Mux_h
    port map (
            O => \N__30704\,
            I => \N__30701\
        );

    \I__5671\ : Odrv4
    port map (
            O => \N__30701\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI1C4K_24\
        );

    \I__5670\ : InMux
    port map (
            O => \N__30698\,
            I => \N__30693\
        );

    \I__5669\ : InMux
    port map (
            O => \N__30697\,
            I => \N__30690\
        );

    \I__5668\ : InMux
    port map (
            O => \N__30696\,
            I => \N__30687\
        );

    \I__5667\ : LocalMux
    port map (
            O => \N__30693\,
            I => \N__30684\
        );

    \I__5666\ : LocalMux
    port map (
            O => \N__30690\,
            I => \N__30680\
        );

    \I__5665\ : LocalMux
    port map (
            O => \N__30687\,
            I => \N__30677\
        );

    \I__5664\ : Span4Mux_v
    port map (
            O => \N__30684\,
            I => \N__30674\
        );

    \I__5663\ : InMux
    port map (
            O => \N__30683\,
            I => \N__30671\
        );

    \I__5662\ : Span4Mux_v
    port map (
            O => \N__30680\,
            I => \N__30668\
        );

    \I__5661\ : Span4Mux_v
    port map (
            O => \N__30677\,
            I => \N__30661\
        );

    \I__5660\ : Span4Mux_h
    port map (
            O => \N__30674\,
            I => \N__30661\
        );

    \I__5659\ : LocalMux
    port map (
            O => \N__30671\,
            I => \N__30661\
        );

    \I__5658\ : Odrv4
    port map (
            O => \N__30668\,
            I => \current_shift_inst.elapsed_time_ns_phase_27\
        );

    \I__5657\ : Odrv4
    port map (
            O => \N__30661\,
            I => \current_shift_inst.elapsed_time_ns_phase_27\
        );

    \I__5656\ : InMux
    port map (
            O => \N__30656\,
            I => \N__30651\
        );

    \I__5655\ : CascadeMux
    port map (
            O => \N__30655\,
            I => \N__30648\
        );

    \I__5654\ : InMux
    port map (
            O => \N__30654\,
            I => \N__30645\
        );

    \I__5653\ : LocalMux
    port map (
            O => \N__30651\,
            I => \N__30641\
        );

    \I__5652\ : InMux
    port map (
            O => \N__30648\,
            I => \N__30638\
        );

    \I__5651\ : LocalMux
    port map (
            O => \N__30645\,
            I => \N__30635\
        );

    \I__5650\ : CascadeMux
    port map (
            O => \N__30644\,
            I => \N__30632\
        );

    \I__5649\ : Span4Mux_h
    port map (
            O => \N__30641\,
            I => \N__30629\
        );

    \I__5648\ : LocalMux
    port map (
            O => \N__30638\,
            I => \N__30624\
        );

    \I__5647\ : Span4Mux_h
    port map (
            O => \N__30635\,
            I => \N__30624\
        );

    \I__5646\ : InMux
    port map (
            O => \N__30632\,
            I => \N__30621\
        );

    \I__5645\ : Odrv4
    port map (
            O => \N__30629\,
            I => \current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0\
        );

    \I__5644\ : Odrv4
    port map (
            O => \N__30624\,
            I => \current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0\
        );

    \I__5643\ : LocalMux
    port map (
            O => \N__30621\,
            I => \current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0\
        );

    \I__5642\ : InMux
    port map (
            O => \N__30614\,
            I => \N__30611\
        );

    \I__5641\ : LocalMux
    port map (
            O => \N__30611\,
            I => \N__30608\
        );

    \I__5640\ : Span4Mux_h
    port map (
            O => \N__30608\,
            I => \N__30605\
        );

    \I__5639\ : Odrv4
    port map (
            O => \N__30605\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIHCE81_26\
        );

    \I__5638\ : InMux
    port map (
            O => \N__30602\,
            I => \N__30599\
        );

    \I__5637\ : LocalMux
    port map (
            O => \N__30599\,
            I => \N__30593\
        );

    \I__5636\ : CascadeMux
    port map (
            O => \N__30598\,
            I => \N__30590\
        );

    \I__5635\ : InMux
    port map (
            O => \N__30597\,
            I => \N__30585\
        );

    \I__5634\ : InMux
    port map (
            O => \N__30596\,
            I => \N__30585\
        );

    \I__5633\ : Span4Mux_h
    port map (
            O => \N__30593\,
            I => \N__30582\
        );

    \I__5632\ : InMux
    port map (
            O => \N__30590\,
            I => \N__30579\
        );

    \I__5631\ : LocalMux
    port map (
            O => \N__30585\,
            I => \N__30576\
        );

    \I__5630\ : Span4Mux_h
    port map (
            O => \N__30582\,
            I => \N__30571\
        );

    \I__5629\ : LocalMux
    port map (
            O => \N__30579\,
            I => \N__30571\
        );

    \I__5628\ : Odrv12
    port map (
            O => \N__30576\,
            I => \current_shift_inst.elapsed_time_ns_phase_23\
        );

    \I__5627\ : Odrv4
    port map (
            O => \N__30571\,
            I => \current_shift_inst.elapsed_time_ns_phase_23\
        );

    \I__5626\ : CascadeMux
    port map (
            O => \N__30566\,
            I => \N__30563\
        );

    \I__5625\ : InMux
    port map (
            O => \N__30563\,
            I => \N__30556\
        );

    \I__5624\ : InMux
    port map (
            O => \N__30562\,
            I => \N__30556\
        );

    \I__5623\ : InMux
    port map (
            O => \N__30561\,
            I => \N__30553\
        );

    \I__5622\ : LocalMux
    port map (
            O => \N__30556\,
            I => \N__30549\
        );

    \I__5621\ : LocalMux
    port map (
            O => \N__30553\,
            I => \N__30546\
        );

    \I__5620\ : CascadeMux
    port map (
            O => \N__30552\,
            I => \N__30543\
        );

    \I__5619\ : Span4Mux_h
    port map (
            O => \N__30549\,
            I => \N__30540\
        );

    \I__5618\ : Span4Mux_h
    port map (
            O => \N__30546\,
            I => \N__30537\
        );

    \I__5617\ : InMux
    port map (
            O => \N__30543\,
            I => \N__30534\
        );

    \I__5616\ : Odrv4
    port map (
            O => \N__30540\,
            I => \current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0\
        );

    \I__5615\ : Odrv4
    port map (
            O => \N__30537\,
            I => \current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0\
        );

    \I__5614\ : LocalMux
    port map (
            O => \N__30534\,
            I => \current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0\
        );

    \I__5613\ : InMux
    port map (
            O => \N__30527\,
            I => \N__30524\
        );

    \I__5612\ : LocalMux
    port map (
            O => \N__30524\,
            I => \N__30521\
        );

    \I__5611\ : Span4Mux_h
    port map (
            O => \N__30521\,
            I => \N__30518\
        );

    \I__5610\ : Odrv4
    port map (
            O => \N__30518\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPB581_22\
        );

    \I__5609\ : CascadeMux
    port map (
            O => \N__30515\,
            I => \N__30512\
        );

    \I__5608\ : InMux
    port map (
            O => \N__30512\,
            I => \N__30509\
        );

    \I__5607\ : LocalMux
    port map (
            O => \N__30509\,
            I => \N__30503\
        );

    \I__5606\ : InMux
    port map (
            O => \N__30508\,
            I => \N__30498\
        );

    \I__5605\ : InMux
    port map (
            O => \N__30507\,
            I => \N__30498\
        );

    \I__5604\ : CascadeMux
    port map (
            O => \N__30506\,
            I => \N__30495\
        );

    \I__5603\ : Span4Mux_v
    port map (
            O => \N__30503\,
            I => \N__30492\
        );

    \I__5602\ : LocalMux
    port map (
            O => \N__30498\,
            I => \N__30489\
        );

    \I__5601\ : InMux
    port map (
            O => \N__30495\,
            I => \N__30486\
        );

    \I__5600\ : Span4Mux_h
    port map (
            O => \N__30492\,
            I => \N__30483\
        );

    \I__5599\ : Span12Mux_v
    port map (
            O => \N__30489\,
            I => \N__30480\
        );

    \I__5598\ : LocalMux
    port map (
            O => \N__30486\,
            I => \N__30477\
        );

    \I__5597\ : Odrv4
    port map (
            O => \N__30483\,
            I => \current_shift_inst.elapsed_time_ns_phase_22\
        );

    \I__5596\ : Odrv12
    port map (
            O => \N__30480\,
            I => \current_shift_inst.elapsed_time_ns_phase_22\
        );

    \I__5595\ : Odrv4
    port map (
            O => \N__30477\,
            I => \current_shift_inst.elapsed_time_ns_phase_22\
        );

    \I__5594\ : CascadeMux
    port map (
            O => \N__30470\,
            I => \N__30467\
        );

    \I__5593\ : InMux
    port map (
            O => \N__30467\,
            I => \N__30460\
        );

    \I__5592\ : InMux
    port map (
            O => \N__30466\,
            I => \N__30460\
        );

    \I__5591\ : InMux
    port map (
            O => \N__30465\,
            I => \N__30456\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__30460\,
            I => \N__30453\
        );

    \I__5589\ : CascadeMux
    port map (
            O => \N__30459\,
            I => \N__30450\
        );

    \I__5588\ : LocalMux
    port map (
            O => \N__30456\,
            I => \N__30447\
        );

    \I__5587\ : Span4Mux_h
    port map (
            O => \N__30453\,
            I => \N__30444\
        );

    \I__5586\ : InMux
    port map (
            O => \N__30450\,
            I => \N__30441\
        );

    \I__5585\ : Odrv12
    port map (
            O => \N__30447\,
            I => \current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0\
        );

    \I__5584\ : Odrv4
    port map (
            O => \N__30444\,
            I => \current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0\
        );

    \I__5583\ : LocalMux
    port map (
            O => \N__30441\,
            I => \current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0\
        );

    \I__5582\ : CascadeMux
    port map (
            O => \N__30434\,
            I => \N__30431\
        );

    \I__5581\ : InMux
    port map (
            O => \N__30431\,
            I => \N__30428\
        );

    \I__5580\ : LocalMux
    port map (
            O => \N__30428\,
            I => \N__30425\
        );

    \I__5579\ : Span4Mux_v
    port map (
            O => \N__30425\,
            I => \N__30422\
        );

    \I__5578\ : Odrv4
    port map (
            O => \N__30422\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIR32K_22\
        );

    \I__5577\ : CascadeMux
    port map (
            O => \N__30419\,
            I => \N__30416\
        );

    \I__5576\ : InMux
    port map (
            O => \N__30416\,
            I => \N__30413\
        );

    \I__5575\ : LocalMux
    port map (
            O => \N__30413\,
            I => \N__30410\
        );

    \I__5574\ : Odrv4
    port map (
            O => \N__30410\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\
        );

    \I__5573\ : CascadeMux
    port map (
            O => \N__30407\,
            I => \N__30404\
        );

    \I__5572\ : InMux
    port map (
            O => \N__30404\,
            I => \N__30399\
        );

    \I__5571\ : InMux
    port map (
            O => \N__30403\,
            I => \N__30396\
        );

    \I__5570\ : CascadeMux
    port map (
            O => \N__30402\,
            I => \N__30393\
        );

    \I__5569\ : LocalMux
    port map (
            O => \N__30399\,
            I => \N__30389\
        );

    \I__5568\ : LocalMux
    port map (
            O => \N__30396\,
            I => \N__30386\
        );

    \I__5567\ : InMux
    port map (
            O => \N__30393\,
            I => \N__30381\
        );

    \I__5566\ : InMux
    port map (
            O => \N__30392\,
            I => \N__30381\
        );

    \I__5565\ : Span12Mux_h
    port map (
            O => \N__30389\,
            I => \N__30378\
        );

    \I__5564\ : Span4Mux_h
    port map (
            O => \N__30386\,
            I => \N__30375\
        );

    \I__5563\ : LocalMux
    port map (
            O => \N__30381\,
            I => \N__30372\
        );

    \I__5562\ : Odrv12
    port map (
            O => \N__30378\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__5561\ : Odrv4
    port map (
            O => \N__30375\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__5560\ : Odrv12
    port map (
            O => \N__30372\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__5559\ : InMux
    port map (
            O => \N__30365\,
            I => \N__30362\
        );

    \I__5558\ : LocalMux
    port map (
            O => \N__30362\,
            I => \N__30359\
        );

    \I__5557\ : Odrv4
    port map (
            O => \N__30359\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\
        );

    \I__5556\ : InMux
    port map (
            O => \N__30356\,
            I => \N__30353\
        );

    \I__5555\ : LocalMux
    port map (
            O => \N__30353\,
            I => \N__30350\
        );

    \I__5554\ : Span4Mux_h
    port map (
            O => \N__30350\,
            I => \N__30344\
        );

    \I__5553\ : InMux
    port map (
            O => \N__30349\,
            I => \N__30341\
        );

    \I__5552\ : InMux
    port map (
            O => \N__30348\,
            I => \N__30336\
        );

    \I__5551\ : InMux
    port map (
            O => \N__30347\,
            I => \N__30336\
        );

    \I__5550\ : Span4Mux_h
    port map (
            O => \N__30344\,
            I => \N__30333\
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__30341\,
            I => \N__30330\
        );

    \I__5548\ : LocalMux
    port map (
            O => \N__30336\,
            I => \N__30327\
        );

    \I__5547\ : Odrv4
    port map (
            O => \N__30333\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__5546\ : Odrv4
    port map (
            O => \N__30330\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__5545\ : Odrv4
    port map (
            O => \N__30327\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__5544\ : CascadeMux
    port map (
            O => \N__30320\,
            I => \phase_controller_inst1.stoper_hc.un1_m5_iZ0Z_1_cascade_\
        );

    \I__5543\ : CascadeMux
    port map (
            O => \N__30317\,
            I => \phase_controller_inst1.stoper_hc.un1_N_4_cascade_\
        );

    \I__5542\ : InMux
    port map (
            O => \N__30314\,
            I => \N__30311\
        );

    \I__5541\ : LocalMux
    port map (
            O => \N__30311\,
            I => \current_shift_inst.S1_sync_prevZ0\
        );

    \I__5540\ : InMux
    port map (
            O => \N__30308\,
            I => \N__30305\
        );

    \I__5539\ : LocalMux
    port map (
            O => \N__30305\,
            I => \current_shift_inst.S1_syncZ0Z0\
        );

    \I__5538\ : InMux
    port map (
            O => \N__30302\,
            I => \N__30296\
        );

    \I__5537\ : InMux
    port map (
            O => \N__30301\,
            I => \N__30296\
        );

    \I__5536\ : LocalMux
    port map (
            O => \N__30296\,
            I => \current_shift_inst.S1_syncZ0Z1\
        );

    \I__5535\ : InMux
    port map (
            O => \N__30293\,
            I => \N__30290\
        );

    \I__5534\ : LocalMux
    port map (
            O => \N__30290\,
            I => \N__30286\
        );

    \I__5533\ : CascadeMux
    port map (
            O => \N__30289\,
            I => \N__30282\
        );

    \I__5532\ : Span4Mux_h
    port map (
            O => \N__30286\,
            I => \N__30275\
        );

    \I__5531\ : InMux
    port map (
            O => \N__30285\,
            I => \N__30272\
        );

    \I__5530\ : InMux
    port map (
            O => \N__30282\,
            I => \N__30265\
        );

    \I__5529\ : InMux
    port map (
            O => \N__30281\,
            I => \N__30265\
        );

    \I__5528\ : InMux
    port map (
            O => \N__30280\,
            I => \N__30265\
        );

    \I__5527\ : InMux
    port map (
            O => \N__30279\,
            I => \N__30262\
        );

    \I__5526\ : InMux
    port map (
            O => \N__30278\,
            I => \N__30259\
        );

    \I__5525\ : Odrv4
    port map (
            O => \N__30275\,
            I => \current_shift_inst.meas_stateZ0Z_0\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__30272\,
            I => \current_shift_inst.meas_stateZ0Z_0\
        );

    \I__5523\ : LocalMux
    port map (
            O => \N__30265\,
            I => \current_shift_inst.meas_stateZ0Z_0\
        );

    \I__5522\ : LocalMux
    port map (
            O => \N__30262\,
            I => \current_shift_inst.meas_stateZ0Z_0\
        );

    \I__5521\ : LocalMux
    port map (
            O => \N__30259\,
            I => \current_shift_inst.meas_stateZ0Z_0\
        );

    \I__5520\ : InMux
    port map (
            O => \N__30248\,
            I => \N__30237\
        );

    \I__5519\ : InMux
    port map (
            O => \N__30247\,
            I => \N__30237\
        );

    \I__5518\ : InMux
    port map (
            O => \N__30246\,
            I => \N__30237\
        );

    \I__5517\ : InMux
    port map (
            O => \N__30245\,
            I => \N__30234\
        );

    \I__5516\ : InMux
    port map (
            O => \N__30244\,
            I => \N__30229\
        );

    \I__5515\ : LocalMux
    port map (
            O => \N__30237\,
            I => \N__30226\
        );

    \I__5514\ : LocalMux
    port map (
            O => \N__30234\,
            I => \N__30223\
        );

    \I__5513\ : InMux
    port map (
            O => \N__30233\,
            I => \N__30220\
        );

    \I__5512\ : InMux
    port map (
            O => \N__30232\,
            I => \N__30217\
        );

    \I__5511\ : LocalMux
    port map (
            O => \N__30229\,
            I => \N__30210\
        );

    \I__5510\ : Span4Mux_v
    port map (
            O => \N__30226\,
            I => \N__30210\
        );

    \I__5509\ : Span4Mux_v
    port map (
            O => \N__30223\,
            I => \N__30210\
        );

    \I__5508\ : LocalMux
    port map (
            O => \N__30220\,
            I => \current_shift_inst.S1_riseZ0\
        );

    \I__5507\ : LocalMux
    port map (
            O => \N__30217\,
            I => \current_shift_inst.S1_riseZ0\
        );

    \I__5506\ : Odrv4
    port map (
            O => \N__30210\,
            I => \current_shift_inst.S1_riseZ0\
        );

    \I__5505\ : InMux
    port map (
            O => \N__30203\,
            I => \N__30199\
        );

    \I__5504\ : InMux
    port map (
            O => \N__30202\,
            I => \N__30195\
        );

    \I__5503\ : LocalMux
    port map (
            O => \N__30199\,
            I => \N__30191\
        );

    \I__5502\ : InMux
    port map (
            O => \N__30198\,
            I => \N__30188\
        );

    \I__5501\ : LocalMux
    port map (
            O => \N__30195\,
            I => \N__30185\
        );

    \I__5500\ : InMux
    port map (
            O => \N__30194\,
            I => \N__30181\
        );

    \I__5499\ : Span12Mux_s8_h
    port map (
            O => \N__30191\,
            I => \N__30178\
        );

    \I__5498\ : LocalMux
    port map (
            O => \N__30188\,
            I => \N__30175\
        );

    \I__5497\ : Span4Mux_h
    port map (
            O => \N__30185\,
            I => \N__30172\
        );

    \I__5496\ : InMux
    port map (
            O => \N__30184\,
            I => \N__30169\
        );

    \I__5495\ : LocalMux
    port map (
            O => \N__30181\,
            I => \N__30164\
        );

    \I__5494\ : Span12Mux_v
    port map (
            O => \N__30178\,
            I => \N__30164\
        );

    \I__5493\ : Span4Mux_h
    port map (
            O => \N__30175\,
            I => \N__30161\
        );

    \I__5492\ : Odrv4
    port map (
            O => \N__30172\,
            I => \current_shift_inst.phase_validZ0\
        );

    \I__5491\ : LocalMux
    port map (
            O => \N__30169\,
            I => \current_shift_inst.phase_validZ0\
        );

    \I__5490\ : Odrv12
    port map (
            O => \N__30164\,
            I => \current_shift_inst.phase_validZ0\
        );

    \I__5489\ : Odrv4
    port map (
            O => \N__30161\,
            I => \current_shift_inst.phase_validZ0\
        );

    \I__5488\ : InMux
    port map (
            O => \N__30152\,
            I => \N__30149\
        );

    \I__5487\ : LocalMux
    port map (
            O => \N__30149\,
            I => \N__30146\
        );

    \I__5486\ : Span4Mux_h
    port map (
            O => \N__30146\,
            I => \N__30143\
        );

    \I__5485\ : Span4Mux_v
    port map (
            O => \N__30143\,
            I => \N__30140\
        );

    \I__5484\ : Odrv4
    port map (
            O => \N__30140\,
            I => il_min_comp1_c
        );

    \I__5483\ : InMux
    port map (
            O => \N__30137\,
            I => \N__30134\
        );

    \I__5482\ : LocalMux
    port map (
            O => \N__30134\,
            I => \il_min_comp1_D1\
        );

    \I__5481\ : InMux
    port map (
            O => \N__30131\,
            I => \N__30128\
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__30128\,
            I => \il_min_comp2_D1\
        );

    \I__5479\ : InMux
    port map (
            O => \N__30125\,
            I => \N__30121\
        );

    \I__5478\ : InMux
    port map (
            O => \N__30124\,
            I => \N__30118\
        );

    \I__5477\ : LocalMux
    port map (
            O => \N__30121\,
            I => \N__30113\
        );

    \I__5476\ : LocalMux
    port map (
            O => \N__30118\,
            I => \N__30110\
        );

    \I__5475\ : InMux
    port map (
            O => \N__30117\,
            I => \N__30105\
        );

    \I__5474\ : InMux
    port map (
            O => \N__30116\,
            I => \N__30105\
        );

    \I__5473\ : Span4Mux_h
    port map (
            O => \N__30113\,
            I => \N__30101\
        );

    \I__5472\ : Span4Mux_v
    port map (
            O => \N__30110\,
            I => \N__30096\
        );

    \I__5471\ : LocalMux
    port map (
            O => \N__30105\,
            I => \N__30096\
        );

    \I__5470\ : InMux
    port map (
            O => \N__30104\,
            I => \N__30093\
        );

    \I__5469\ : Odrv4
    port map (
            O => \N__30101\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_20\
        );

    \I__5468\ : Odrv4
    port map (
            O => \N__30096\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_20\
        );

    \I__5467\ : LocalMux
    port map (
            O => \N__30093\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_20\
        );

    \I__5466\ : CascadeMux
    port map (
            O => \N__30086\,
            I => \N__30083\
        );

    \I__5465\ : InMux
    port map (
            O => \N__30083\,
            I => \N__30079\
        );

    \I__5464\ : InMux
    port map (
            O => \N__30082\,
            I => \N__30076\
        );

    \I__5463\ : LocalMux
    port map (
            O => \N__30079\,
            I => \N__30068\
        );

    \I__5462\ : LocalMux
    port map (
            O => \N__30076\,
            I => \N__30068\
        );

    \I__5461\ : InMux
    port map (
            O => \N__30075\,
            I => \N__30065\
        );

    \I__5460\ : InMux
    port map (
            O => \N__30074\,
            I => \N__30060\
        );

    \I__5459\ : InMux
    port map (
            O => \N__30073\,
            I => \N__30060\
        );

    \I__5458\ : Span4Mux_v
    port map (
            O => \N__30068\,
            I => \N__30057\
        );

    \I__5457\ : LocalMux
    port map (
            O => \N__30065\,
            I => \N__30054\
        );

    \I__5456\ : LocalMux
    port map (
            O => \N__30060\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\
        );

    \I__5455\ : Odrv4
    port map (
            O => \N__30057\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\
        );

    \I__5454\ : Odrv4
    port map (
            O => \N__30054\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\
        );

    \I__5453\ : InMux
    port map (
            O => \N__30047\,
            I => \N__30044\
        );

    \I__5452\ : LocalMux
    port map (
            O => \N__30044\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\
        );

    \I__5451\ : InMux
    port map (
            O => \N__30041\,
            I => \N__30037\
        );

    \I__5450\ : CascadeMux
    port map (
            O => \N__30040\,
            I => \N__30034\
        );

    \I__5449\ : LocalMux
    port map (
            O => \N__30037\,
            I => \N__30031\
        );

    \I__5448\ : InMux
    port map (
            O => \N__30034\,
            I => \N__30028\
        );

    \I__5447\ : Span4Mux_v
    port map (
            O => \N__30031\,
            I => \N__30025\
        );

    \I__5446\ : LocalMux
    port map (
            O => \N__30028\,
            I => \N__30021\
        );

    \I__5445\ : Span4Mux_h
    port map (
            O => \N__30025\,
            I => \N__30018\
        );

    \I__5444\ : InMux
    port map (
            O => \N__30024\,
            I => \N__30015\
        );

    \I__5443\ : Odrv12
    port map (
            O => \N__30021\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__5442\ : Odrv4
    port map (
            O => \N__30018\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__30015\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__5440\ : CascadeMux
    port map (
            O => \N__30008\,
            I => \N__30005\
        );

    \I__5439\ : InMux
    port map (
            O => \N__30005\,
            I => \N__30002\
        );

    \I__5438\ : LocalMux
    port map (
            O => \N__30002\,
            I => \N__29999\
        );

    \I__5437\ : Span4Mux_h
    port map (
            O => \N__29999\,
            I => \N__29996\
        );

    \I__5436\ : Odrv4
    port map (
            O => \N__29996\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\
        );

    \I__5435\ : InMux
    port map (
            O => \N__29993\,
            I => \N__29990\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__29990\,
            I => \current_shift_inst.un4_control_input_axb_17\
        );

    \I__5433\ : InMux
    port map (
            O => \N__29987\,
            I => \N__29984\
        );

    \I__5432\ : LocalMux
    port map (
            O => \N__29984\,
            I => \N__29981\
        );

    \I__5431\ : Odrv4
    port map (
            O => \N__29981\,
            I => \current_shift_inst.un4_control_input_axb_21\
        );

    \I__5430\ : InMux
    port map (
            O => \N__29978\,
            I => \N__29975\
        );

    \I__5429\ : LocalMux
    port map (
            O => \N__29975\,
            I => \current_shift_inst.un4_control_input_axb_26\
        );

    \I__5428\ : InMux
    port map (
            O => \N__29972\,
            I => \N__29969\
        );

    \I__5427\ : LocalMux
    port map (
            O => \N__29969\,
            I => \N__29965\
        );

    \I__5426\ : InMux
    port map (
            O => \N__29968\,
            I => \N__29962\
        );

    \I__5425\ : Span4Mux_v
    port map (
            O => \N__29965\,
            I => \N__29959\
        );

    \I__5424\ : LocalMux
    port map (
            O => \N__29962\,
            I => \N__29956\
        );

    \I__5423\ : Span4Mux_v
    port map (
            O => \N__29959\,
            I => \N__29953\
        );

    \I__5422\ : Odrv4
    port map (
            O => \N__29956\,
            I => \current_shift_inst.z_31\
        );

    \I__5421\ : Odrv4
    port map (
            O => \N__29953\,
            I => \current_shift_inst.z_31\
        );

    \I__5420\ : CascadeMux
    port map (
            O => \N__29948\,
            I => \N__29944\
        );

    \I__5419\ : InMux
    port map (
            O => \N__29947\,
            I => \N__29941\
        );

    \I__5418\ : InMux
    port map (
            O => \N__29944\,
            I => \N__29938\
        );

    \I__5417\ : LocalMux
    port map (
            O => \N__29941\,
            I => \N__29933\
        );

    \I__5416\ : LocalMux
    port map (
            O => \N__29938\,
            I => \N__29933\
        );

    \I__5415\ : Span4Mux_h
    port map (
            O => \N__29933\,
            I => \N__29930\
        );

    \I__5414\ : Span4Mux_v
    port map (
            O => \N__29930\,
            I => \N__29927\
        );

    \I__5413\ : Odrv4
    port map (
            O => \N__29927\,
            I => \current_shift_inst.z_i_31\
        );

    \I__5412\ : InMux
    port map (
            O => \N__29924\,
            I => \N__29921\
        );

    \I__5411\ : LocalMux
    port map (
            O => \N__29921\,
            I => \N__29918\
        );

    \I__5410\ : Odrv4
    port map (
            O => \N__29918\,
            I => \current_shift_inst.un4_control_input_axb_30\
        );

    \I__5409\ : InMux
    port map (
            O => \N__29915\,
            I => \N__29912\
        );

    \I__5408\ : LocalMux
    port map (
            O => \N__29912\,
            I => \N__29909\
        );

    \I__5407\ : Odrv4
    port map (
            O => \N__29909\,
            I => \current_shift_inst.un4_control_input_axb_27\
        );

    \I__5406\ : InMux
    port map (
            O => \N__29906\,
            I => \N__29903\
        );

    \I__5405\ : LocalMux
    port map (
            O => \N__29903\,
            I => \N__29900\
        );

    \I__5404\ : Odrv4
    port map (
            O => \N__29900\,
            I => \current_shift_inst.un4_control_input_axb_29\
        );

    \I__5403\ : InMux
    port map (
            O => \N__29897\,
            I => \N__29894\
        );

    \I__5402\ : LocalMux
    port map (
            O => \N__29894\,
            I => \N__29891\
        );

    \I__5401\ : Odrv4
    port map (
            O => \N__29891\,
            I => \current_shift_inst.un4_control_input_axb_28\
        );

    \I__5400\ : InMux
    port map (
            O => \N__29888\,
            I => \N__29885\
        );

    \I__5399\ : LocalMux
    port map (
            O => \N__29885\,
            I => \current_shift_inst.un4_control_input_axb_12\
        );

    \I__5398\ : InMux
    port map (
            O => \N__29882\,
            I => \N__29879\
        );

    \I__5397\ : LocalMux
    port map (
            O => \N__29879\,
            I => \current_shift_inst.un4_control_input_axb_16\
        );

    \I__5396\ : InMux
    port map (
            O => \N__29876\,
            I => \N__29873\
        );

    \I__5395\ : LocalMux
    port map (
            O => \N__29873\,
            I => \current_shift_inst.un4_control_input_axb_20\
        );

    \I__5394\ : InMux
    port map (
            O => \N__29870\,
            I => \N__29867\
        );

    \I__5393\ : LocalMux
    port map (
            O => \N__29867\,
            I => \current_shift_inst.un4_control_input_axb_18\
        );

    \I__5392\ : InMux
    port map (
            O => \N__29864\,
            I => \N__29861\
        );

    \I__5391\ : LocalMux
    port map (
            O => \N__29861\,
            I => \current_shift_inst.un4_control_input_axb_23\
        );

    \I__5390\ : InMux
    port map (
            O => \N__29858\,
            I => \N__29855\
        );

    \I__5389\ : LocalMux
    port map (
            O => \N__29855\,
            I => \current_shift_inst.un4_control_input_axb_19\
        );

    \I__5388\ : InMux
    port map (
            O => \N__29852\,
            I => \N__29849\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__29849\,
            I => \current_shift_inst.un4_control_input_axb_25\
        );

    \I__5386\ : InMux
    port map (
            O => \N__29846\,
            I => \N__29843\
        );

    \I__5385\ : LocalMux
    port map (
            O => \N__29843\,
            I => \current_shift_inst.un4_control_input_axb_22\
        );

    \I__5384\ : InMux
    port map (
            O => \N__29840\,
            I => \N__29837\
        );

    \I__5383\ : LocalMux
    port map (
            O => \N__29837\,
            I => \current_shift_inst.un4_control_input_axb_24\
        );

    \I__5382\ : InMux
    port map (
            O => \N__29834\,
            I => \N__29831\
        );

    \I__5381\ : LocalMux
    port map (
            O => \N__29831\,
            I => \current_shift_inst.un4_control_input_axb_4\
        );

    \I__5380\ : InMux
    port map (
            O => \N__29828\,
            I => \N__29825\
        );

    \I__5379\ : LocalMux
    port map (
            O => \N__29825\,
            I => \current_shift_inst.un4_control_input_axb_5\
        );

    \I__5378\ : InMux
    port map (
            O => \N__29822\,
            I => \N__29819\
        );

    \I__5377\ : LocalMux
    port map (
            O => \N__29819\,
            I => \current_shift_inst.un4_control_input_axb_6\
        );

    \I__5376\ : CascadeMux
    port map (
            O => \N__29816\,
            I => \N__29813\
        );

    \I__5375\ : InMux
    port map (
            O => \N__29813\,
            I => \N__29810\
        );

    \I__5374\ : LocalMux
    port map (
            O => \N__29810\,
            I => \current_shift_inst.un4_control_input_axb_7\
        );

    \I__5373\ : CascadeMux
    port map (
            O => \N__29807\,
            I => \N__29804\
        );

    \I__5372\ : InMux
    port map (
            O => \N__29804\,
            I => \N__29801\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__29801\,
            I => \current_shift_inst.un4_control_input_axb_8\
        );

    \I__5370\ : InMux
    port map (
            O => \N__29798\,
            I => \N__29795\
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__29795\,
            I => \current_shift_inst.un4_control_input_axb_13\
        );

    \I__5368\ : InMux
    port map (
            O => \N__29792\,
            I => \N__29789\
        );

    \I__5367\ : LocalMux
    port map (
            O => \N__29789\,
            I => \current_shift_inst.un4_control_input_axb_15\
        );

    \I__5366\ : InMux
    port map (
            O => \N__29786\,
            I => \N__29783\
        );

    \I__5365\ : LocalMux
    port map (
            O => \N__29783\,
            I => \current_shift_inst.un4_control_input_axb_9\
        );

    \I__5364\ : InMux
    port map (
            O => \N__29780\,
            I => \N__29777\
        );

    \I__5363\ : LocalMux
    port map (
            O => \N__29777\,
            I => \current_shift_inst.un4_control_input_axb_10\
        );

    \I__5362\ : InMux
    port map (
            O => \N__29774\,
            I => \N__29771\
        );

    \I__5361\ : LocalMux
    port map (
            O => \N__29771\,
            I => \current_shift_inst.un4_control_input_axb_11\
        );

    \I__5360\ : InMux
    port map (
            O => \N__29768\,
            I => \N__29764\
        );

    \I__5359\ : CascadeMux
    port map (
            O => \N__29767\,
            I => \N__29760\
        );

    \I__5358\ : LocalMux
    port map (
            O => \N__29764\,
            I => \N__29757\
        );

    \I__5357\ : InMux
    port map (
            O => \N__29763\,
            I => \N__29754\
        );

    \I__5356\ : InMux
    port map (
            O => \N__29760\,
            I => \N__29751\
        );

    \I__5355\ : Span4Mux_v
    port map (
            O => \N__29757\,
            I => \N__29748\
        );

    \I__5354\ : LocalMux
    port map (
            O => \N__29754\,
            I => \current_shift_inst.elapsed_time_ns_1_fast_31\
        );

    \I__5353\ : LocalMux
    port map (
            O => \N__29751\,
            I => \current_shift_inst.elapsed_time_ns_1_fast_31\
        );

    \I__5352\ : Odrv4
    port map (
            O => \N__29748\,
            I => \current_shift_inst.elapsed_time_ns_1_fast_31\
        );

    \I__5351\ : InMux
    port map (
            O => \N__29741\,
            I => \N__29738\
        );

    \I__5350\ : LocalMux
    port map (
            O => \N__29738\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_1\
        );

    \I__5349\ : InMux
    port map (
            O => \N__29735\,
            I => \N__29732\
        );

    \I__5348\ : LocalMux
    port map (
            O => \N__29732\,
            I => \current_shift_inst.un4_control_input_axb_1\
        );

    \I__5347\ : InMux
    port map (
            O => \N__29729\,
            I => \N__29726\
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__29726\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_2\
        );

    \I__5345\ : InMux
    port map (
            O => \N__29723\,
            I => \N__29720\
        );

    \I__5344\ : LocalMux
    port map (
            O => \N__29720\,
            I => \current_shift_inst.un4_control_input_axb_2\
        );

    \I__5343\ : InMux
    port map (
            O => \N__29717\,
            I => \N__29714\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__29714\,
            I => \current_shift_inst.un4_control_input_axb_14\
        );

    \I__5341\ : InMux
    port map (
            O => \N__29711\,
            I => \N__29708\
        );

    \I__5340\ : LocalMux
    port map (
            O => \N__29708\,
            I => \current_shift_inst.un4_control_input_axb_3\
        );

    \I__5339\ : CascadeMux
    port map (
            O => \N__29705\,
            I => \N__29701\
        );

    \I__5338\ : CascadeMux
    port map (
            O => \N__29704\,
            I => \N__29698\
        );

    \I__5337\ : InMux
    port map (
            O => \N__29701\,
            I => \N__29695\
        );

    \I__5336\ : InMux
    port map (
            O => \N__29698\,
            I => \N__29690\
        );

    \I__5335\ : LocalMux
    port map (
            O => \N__29695\,
            I => \N__29687\
        );

    \I__5334\ : InMux
    port map (
            O => \N__29694\,
            I => \N__29684\
        );

    \I__5333\ : InMux
    port map (
            O => \N__29693\,
            I => \N__29681\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__29690\,
            I => \N__29678\
        );

    \I__5331\ : Span4Mux_v
    port map (
            O => \N__29687\,
            I => \N__29675\
        );

    \I__5330\ : LocalMux
    port map (
            O => \N__29684\,
            I => \N__29672\
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__29681\,
            I => \N__29669\
        );

    \I__5328\ : Span4Mux_v
    port map (
            O => \N__29678\,
            I => \N__29666\
        );

    \I__5327\ : Span4Mux_h
    port map (
            O => \N__29675\,
            I => \N__29659\
        );

    \I__5326\ : Span4Mux_v
    port map (
            O => \N__29672\,
            I => \N__29659\
        );

    \I__5325\ : Span4Mux_v
    port map (
            O => \N__29669\,
            I => \N__29659\
        );

    \I__5324\ : Odrv4
    port map (
            O => \N__29666\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__5323\ : Odrv4
    port map (
            O => \N__29659\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__5322\ : CascadeMux
    port map (
            O => \N__29654\,
            I => \N__29651\
        );

    \I__5321\ : InMux
    port map (
            O => \N__29651\,
            I => \N__29648\
        );

    \I__5320\ : LocalMux
    port map (
            O => \N__29648\,
            I => \N__29645\
        );

    \I__5319\ : Span4Mux_v
    port map (
            O => \N__29645\,
            I => \N__29642\
        );

    \I__5318\ : Odrv4
    port map (
            O => \N__29642\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\
        );

    \I__5317\ : InMux
    port map (
            O => \N__29639\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\
        );

    \I__5316\ : InMux
    port map (
            O => \N__29636\,
            I => \N__29633\
        );

    \I__5315\ : LocalMux
    port map (
            O => \N__29633\,
            I => \N__29628\
        );

    \I__5314\ : InMux
    port map (
            O => \N__29632\,
            I => \N__29625\
        );

    \I__5313\ : CascadeMux
    port map (
            O => \N__29631\,
            I => \N__29622\
        );

    \I__5312\ : Span4Mux_v
    port map (
            O => \N__29628\,
            I => \N__29619\
        );

    \I__5311\ : LocalMux
    port map (
            O => \N__29625\,
            I => \N__29616\
        );

    \I__5310\ : InMux
    port map (
            O => \N__29622\,
            I => \N__29612\
        );

    \I__5309\ : Span4Mux_h
    port map (
            O => \N__29619\,
            I => \N__29607\
        );

    \I__5308\ : Span4Mux_h
    port map (
            O => \N__29616\,
            I => \N__29607\
        );

    \I__5307\ : InMux
    port map (
            O => \N__29615\,
            I => \N__29604\
        );

    \I__5306\ : LocalMux
    port map (
            O => \N__29612\,
            I => \N__29601\
        );

    \I__5305\ : Odrv4
    port map (
            O => \N__29607\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__5304\ : LocalMux
    port map (
            O => \N__29604\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__5303\ : Odrv12
    port map (
            O => \N__29601\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__5302\ : CascadeMux
    port map (
            O => \N__29594\,
            I => \N__29591\
        );

    \I__5301\ : InMux
    port map (
            O => \N__29591\,
            I => \N__29588\
        );

    \I__5300\ : LocalMux
    port map (
            O => \N__29588\,
            I => \N__29585\
        );

    \I__5299\ : Sp12to4
    port map (
            O => \N__29585\,
            I => \N__29582\
        );

    \I__5298\ : Odrv12
    port map (
            O => \N__29582\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\
        );

    \I__5297\ : InMux
    port map (
            O => \N__29579\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\
        );

    \I__5296\ : CascadeMux
    port map (
            O => \N__29576\,
            I => \N__29572\
        );

    \I__5295\ : CascadeMux
    port map (
            O => \N__29575\,
            I => \N__29569\
        );

    \I__5294\ : InMux
    port map (
            O => \N__29572\,
            I => \N__29565\
        );

    \I__5293\ : InMux
    port map (
            O => \N__29569\,
            I => \N__29562\
        );

    \I__5292\ : CascadeMux
    port map (
            O => \N__29568\,
            I => \N__29558\
        );

    \I__5291\ : LocalMux
    port map (
            O => \N__29565\,
            I => \N__29555\
        );

    \I__5290\ : LocalMux
    port map (
            O => \N__29562\,
            I => \N__29552\
        );

    \I__5289\ : InMux
    port map (
            O => \N__29561\,
            I => \N__29549\
        );

    \I__5288\ : InMux
    port map (
            O => \N__29558\,
            I => \N__29546\
        );

    \I__5287\ : Span4Mux_h
    port map (
            O => \N__29555\,
            I => \N__29543\
        );

    \I__5286\ : Span4Mux_h
    port map (
            O => \N__29552\,
            I => \N__29538\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__29549\,
            I => \N__29538\
        );

    \I__5284\ : LocalMux
    port map (
            O => \N__29546\,
            I => \N__29535\
        );

    \I__5283\ : Odrv4
    port map (
            O => \N__29543\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__5282\ : Odrv4
    port map (
            O => \N__29538\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__5281\ : Odrv4
    port map (
            O => \N__29535\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__5280\ : CascadeMux
    port map (
            O => \N__29528\,
            I => \N__29525\
        );

    \I__5279\ : InMux
    port map (
            O => \N__29525\,
            I => \N__29522\
        );

    \I__5278\ : LocalMux
    port map (
            O => \N__29522\,
            I => \N__29519\
        );

    \I__5277\ : Span4Mux_h
    port map (
            O => \N__29519\,
            I => \N__29516\
        );

    \I__5276\ : Odrv4
    port map (
            O => \N__29516\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\
        );

    \I__5275\ : InMux
    port map (
            O => \N__29513\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\
        );

    \I__5274\ : InMux
    port map (
            O => \N__29510\,
            I => \N__29503\
        );

    \I__5273\ : CascadeMux
    port map (
            O => \N__29509\,
            I => \N__29500\
        );

    \I__5272\ : CascadeMux
    port map (
            O => \N__29508\,
            I => \N__29496\
        );

    \I__5271\ : CascadeMux
    port map (
            O => \N__29507\,
            I => \N__29492\
        );

    \I__5270\ : CascadeMux
    port map (
            O => \N__29506\,
            I => \N__29488\
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__29503\,
            I => \N__29485\
        );

    \I__5268\ : InMux
    port map (
            O => \N__29500\,
            I => \N__29470\
        );

    \I__5267\ : InMux
    port map (
            O => \N__29499\,
            I => \N__29470\
        );

    \I__5266\ : InMux
    port map (
            O => \N__29496\,
            I => \N__29470\
        );

    \I__5265\ : InMux
    port map (
            O => \N__29495\,
            I => \N__29470\
        );

    \I__5264\ : InMux
    port map (
            O => \N__29492\,
            I => \N__29470\
        );

    \I__5263\ : InMux
    port map (
            O => \N__29491\,
            I => \N__29470\
        );

    \I__5262\ : InMux
    port map (
            O => \N__29488\,
            I => \N__29470\
        );

    \I__5261\ : Span4Mux_v
    port map (
            O => \N__29485\,
            I => \N__29467\
        );

    \I__5260\ : LocalMux
    port map (
            O => \N__29470\,
            I => \N__29464\
        );

    \I__5259\ : Span4Mux_v
    port map (
            O => \N__29467\,
            I => \N__29461\
        );

    \I__5258\ : Span4Mux_h
    port map (
            O => \N__29464\,
            I => \N__29458\
        );

    \I__5257\ : Odrv4
    port map (
            O => \N__29461\,
            I => \current_shift_inst.control_inputZ0Z_25\
        );

    \I__5256\ : Odrv4
    port map (
            O => \N__29458\,
            I => \current_shift_inst.control_inputZ0Z_25\
        );

    \I__5255\ : InMux
    port map (
            O => \N__29453\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_30\
        );

    \I__5254\ : CascadeMux
    port map (
            O => \N__29450\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto31_cZ0Z_0_cascade_\
        );

    \I__5253\ : InMux
    port map (
            O => \N__29447\,
            I => \N__29443\
        );

    \I__5252\ : InMux
    port map (
            O => \N__29446\,
            I => \N__29440\
        );

    \I__5251\ : LocalMux
    port map (
            O => \N__29443\,
            I => \N__29437\
        );

    \I__5250\ : LocalMux
    port map (
            O => \N__29440\,
            I => \N__29434\
        );

    \I__5249\ : Span4Mux_h
    port map (
            O => \N__29437\,
            I => \N__29431\
        );

    \I__5248\ : Span4Mux_v
    port map (
            O => \N__29434\,
            I => \N__29428\
        );

    \I__5247\ : Odrv4
    port map (
            O => \N__29431\,
            I => \current_shift_inst.control_inputZ0Z_20\
        );

    \I__5246\ : Odrv4
    port map (
            O => \N__29428\,
            I => \current_shift_inst.control_inputZ0Z_20\
        );

    \I__5245\ : InMux
    port map (
            O => \N__29423\,
            I => \N__29419\
        );

    \I__5244\ : CascadeMux
    port map (
            O => \N__29422\,
            I => \N__29414\
        );

    \I__5243\ : LocalMux
    port map (
            O => \N__29419\,
            I => \N__29411\
        );

    \I__5242\ : InMux
    port map (
            O => \N__29418\,
            I => \N__29408\
        );

    \I__5241\ : InMux
    port map (
            O => \N__29417\,
            I => \N__29405\
        );

    \I__5240\ : InMux
    port map (
            O => \N__29414\,
            I => \N__29402\
        );

    \I__5239\ : Span4Mux_h
    port map (
            O => \N__29411\,
            I => \N__29395\
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__29408\,
            I => \N__29395\
        );

    \I__5237\ : LocalMux
    port map (
            O => \N__29405\,
            I => \N__29395\
        );

    \I__5236\ : LocalMux
    port map (
            O => \N__29402\,
            I => \N__29392\
        );

    \I__5235\ : Span4Mux_h
    port map (
            O => \N__29395\,
            I => \N__29389\
        );

    \I__5234\ : Odrv12
    port map (
            O => \N__29392\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__5233\ : Odrv4
    port map (
            O => \N__29389\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__5232\ : CascadeMux
    port map (
            O => \N__29384\,
            I => \N__29381\
        );

    \I__5231\ : InMux
    port map (
            O => \N__29381\,
            I => \N__29378\
        );

    \I__5230\ : LocalMux
    port map (
            O => \N__29378\,
            I => \N__29375\
        );

    \I__5229\ : Span4Mux_h
    port map (
            O => \N__29375\,
            I => \N__29372\
        );

    \I__5228\ : Odrv4
    port map (
            O => \N__29372\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\
        );

    \I__5227\ : InMux
    port map (
            O => \N__29369\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\
        );

    \I__5226\ : CascadeMux
    port map (
            O => \N__29366\,
            I => \N__29363\
        );

    \I__5225\ : InMux
    port map (
            O => \N__29363\,
            I => \N__29360\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__29360\,
            I => \N__29357\
        );

    \I__5223\ : Span4Mux_h
    port map (
            O => \N__29357\,
            I => \N__29351\
        );

    \I__5222\ : InMux
    port map (
            O => \N__29356\,
            I => \N__29348\
        );

    \I__5221\ : InMux
    port map (
            O => \N__29355\,
            I => \N__29343\
        );

    \I__5220\ : InMux
    port map (
            O => \N__29354\,
            I => \N__29343\
        );

    \I__5219\ : Odrv4
    port map (
            O => \N__29351\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__5218\ : LocalMux
    port map (
            O => \N__29348\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__5217\ : LocalMux
    port map (
            O => \N__29343\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__5216\ : CascadeMux
    port map (
            O => \N__29336\,
            I => \N__29332\
        );

    \I__5215\ : InMux
    port map (
            O => \N__29335\,
            I => \N__29329\
        );

    \I__5214\ : InMux
    port map (
            O => \N__29332\,
            I => \N__29326\
        );

    \I__5213\ : LocalMux
    port map (
            O => \N__29329\,
            I => \N__29323\
        );

    \I__5212\ : LocalMux
    port map (
            O => \N__29326\,
            I => \N__29320\
        );

    \I__5211\ : Span4Mux_v
    port map (
            O => \N__29323\,
            I => \N__29317\
        );

    \I__5210\ : Span12Mux_v
    port map (
            O => \N__29320\,
            I => \N__29314\
        );

    \I__5209\ : Odrv4
    port map (
            O => \N__29317\,
            I => \current_shift_inst.control_inputZ0Z_21\
        );

    \I__5208\ : Odrv12
    port map (
            O => \N__29314\,
            I => \current_shift_inst.control_inputZ0Z_21\
        );

    \I__5207\ : CascadeMux
    port map (
            O => \N__29309\,
            I => \N__29306\
        );

    \I__5206\ : InMux
    port map (
            O => \N__29306\,
            I => \N__29303\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__29303\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\
        );

    \I__5204\ : InMux
    port map (
            O => \N__29300\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\
        );

    \I__5203\ : CascadeMux
    port map (
            O => \N__29297\,
            I => \N__29293\
        );

    \I__5202\ : InMux
    port map (
            O => \N__29296\,
            I => \N__29288\
        );

    \I__5201\ : InMux
    port map (
            O => \N__29293\,
            I => \N__29285\
        );

    \I__5200\ : CascadeMux
    port map (
            O => \N__29292\,
            I => \N__29282\
        );

    \I__5199\ : InMux
    port map (
            O => \N__29291\,
            I => \N__29279\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__29288\,
            I => \N__29274\
        );

    \I__5197\ : LocalMux
    port map (
            O => \N__29285\,
            I => \N__29274\
        );

    \I__5196\ : InMux
    port map (
            O => \N__29282\,
            I => \N__29271\
        );

    \I__5195\ : LocalMux
    port map (
            O => \N__29279\,
            I => \N__29268\
        );

    \I__5194\ : Span4Mux_h
    port map (
            O => \N__29274\,
            I => \N__29265\
        );

    \I__5193\ : LocalMux
    port map (
            O => \N__29271\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__5192\ : Odrv4
    port map (
            O => \N__29268\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__5191\ : Odrv4
    port map (
            O => \N__29265\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__5190\ : CascadeMux
    port map (
            O => \N__29258\,
            I => \N__29254\
        );

    \I__5189\ : InMux
    port map (
            O => \N__29257\,
            I => \N__29251\
        );

    \I__5188\ : InMux
    port map (
            O => \N__29254\,
            I => \N__29248\
        );

    \I__5187\ : LocalMux
    port map (
            O => \N__29251\,
            I => \N__29245\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__29248\,
            I => \N__29242\
        );

    \I__5185\ : Span4Mux_h
    port map (
            O => \N__29245\,
            I => \N__29237\
        );

    \I__5184\ : Span4Mux_h
    port map (
            O => \N__29242\,
            I => \N__29237\
        );

    \I__5183\ : Odrv4
    port map (
            O => \N__29237\,
            I => \current_shift_inst.control_inputZ0Z_22\
        );

    \I__5182\ : InMux
    port map (
            O => \N__29234\,
            I => \N__29231\
        );

    \I__5181\ : LocalMux
    port map (
            O => \N__29231\,
            I => \N__29228\
        );

    \I__5180\ : Odrv4
    port map (
            O => \N__29228\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\
        );

    \I__5179\ : InMux
    port map (
            O => \N__29225\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\
        );

    \I__5178\ : InMux
    port map (
            O => \N__29222\,
            I => \N__29219\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__29219\,
            I => \N__29213\
        );

    \I__5176\ : InMux
    port map (
            O => \N__29218\,
            I => \N__29210\
        );

    \I__5175\ : InMux
    port map (
            O => \N__29217\,
            I => \N__29207\
        );

    \I__5174\ : InMux
    port map (
            O => \N__29216\,
            I => \N__29204\
        );

    \I__5173\ : Span4Mux_h
    port map (
            O => \N__29213\,
            I => \N__29201\
        );

    \I__5172\ : LocalMux
    port map (
            O => \N__29210\,
            I => \N__29198\
        );

    \I__5171\ : LocalMux
    port map (
            O => \N__29207\,
            I => \N__29193\
        );

    \I__5170\ : LocalMux
    port map (
            O => \N__29204\,
            I => \N__29193\
        );

    \I__5169\ : Odrv4
    port map (
            O => \N__29201\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__5168\ : Odrv4
    port map (
            O => \N__29198\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__5167\ : Odrv4
    port map (
            O => \N__29193\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__5166\ : CascadeMux
    port map (
            O => \N__29186\,
            I => \N__29182\
        );

    \I__5165\ : InMux
    port map (
            O => \N__29185\,
            I => \N__29179\
        );

    \I__5164\ : InMux
    port map (
            O => \N__29182\,
            I => \N__29176\
        );

    \I__5163\ : LocalMux
    port map (
            O => \N__29179\,
            I => \N__29173\
        );

    \I__5162\ : LocalMux
    port map (
            O => \N__29176\,
            I => \N__29170\
        );

    \I__5161\ : Span4Mux_v
    port map (
            O => \N__29173\,
            I => \N__29165\
        );

    \I__5160\ : Span4Mux_v
    port map (
            O => \N__29170\,
            I => \N__29165\
        );

    \I__5159\ : Odrv4
    port map (
            O => \N__29165\,
            I => \current_shift_inst.control_inputZ0Z_23\
        );

    \I__5158\ : CascadeMux
    port map (
            O => \N__29162\,
            I => \N__29159\
        );

    \I__5157\ : InMux
    port map (
            O => \N__29159\,
            I => \N__29156\
        );

    \I__5156\ : LocalMux
    port map (
            O => \N__29156\,
            I => \N__29153\
        );

    \I__5155\ : Odrv4
    port map (
            O => \N__29153\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\
        );

    \I__5154\ : InMux
    port map (
            O => \N__29150\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\
        );

    \I__5153\ : CascadeMux
    port map (
            O => \N__29147\,
            I => \N__29143\
        );

    \I__5152\ : InMux
    port map (
            O => \N__29146\,
            I => \N__29140\
        );

    \I__5151\ : InMux
    port map (
            O => \N__29143\,
            I => \N__29137\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__29140\,
            I => \N__29134\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__29137\,
            I => \N__29131\
        );

    \I__5148\ : Span12Mux_v
    port map (
            O => \N__29134\,
            I => \N__29128\
        );

    \I__5147\ : Span4Mux_h
    port map (
            O => \N__29131\,
            I => \N__29125\
        );

    \I__5146\ : Odrv12
    port map (
            O => \N__29128\,
            I => \current_shift_inst.control_inputZ0Z_24\
        );

    \I__5145\ : Odrv4
    port map (
            O => \N__29125\,
            I => \current_shift_inst.control_inputZ0Z_24\
        );

    \I__5144\ : InMux
    port map (
            O => \N__29120\,
            I => \bfn_11_13_0_\
        );

    \I__5143\ : InMux
    port map (
            O => \N__29117\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\
        );

    \I__5142\ : CascadeMux
    port map (
            O => \N__29114\,
            I => \N__29111\
        );

    \I__5141\ : InMux
    port map (
            O => \N__29111\,
            I => \N__29108\
        );

    \I__5140\ : LocalMux
    port map (
            O => \N__29108\,
            I => \N__29104\
        );

    \I__5139\ : CascadeMux
    port map (
            O => \N__29107\,
            I => \N__29101\
        );

    \I__5138\ : Span4Mux_v
    port map (
            O => \N__29104\,
            I => \N__29097\
        );

    \I__5137\ : InMux
    port map (
            O => \N__29101\,
            I => \N__29094\
        );

    \I__5136\ : CascadeMux
    port map (
            O => \N__29100\,
            I => \N__29090\
        );

    \I__5135\ : Span4Mux_h
    port map (
            O => \N__29097\,
            I => \N__29087\
        );

    \I__5134\ : LocalMux
    port map (
            O => \N__29094\,
            I => \N__29084\
        );

    \I__5133\ : InMux
    port map (
            O => \N__29093\,
            I => \N__29079\
        );

    \I__5132\ : InMux
    port map (
            O => \N__29090\,
            I => \N__29079\
        );

    \I__5131\ : Odrv4
    port map (
            O => \N__29087\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__5130\ : Odrv4
    port map (
            O => \N__29084\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__5129\ : LocalMux
    port map (
            O => \N__29079\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__5128\ : InMux
    port map (
            O => \N__29072\,
            I => \N__29069\
        );

    \I__5127\ : LocalMux
    port map (
            O => \N__29069\,
            I => \N__29066\
        );

    \I__5126\ : Odrv4
    port map (
            O => \N__29066\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\
        );

    \I__5125\ : InMux
    port map (
            O => \N__29063\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\
        );

    \I__5124\ : InMux
    port map (
            O => \N__29060\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\
        );

    \I__5123\ : CascadeMux
    port map (
            O => \N__29057\,
            I => \N__29053\
        );

    \I__5122\ : InMux
    port map (
            O => \N__29056\,
            I => \N__29050\
        );

    \I__5121\ : InMux
    port map (
            O => \N__29053\,
            I => \N__29047\
        );

    \I__5120\ : LocalMux
    port map (
            O => \N__29050\,
            I => \N__29042\
        );

    \I__5119\ : LocalMux
    port map (
            O => \N__29047\,
            I => \N__29039\
        );

    \I__5118\ : InMux
    port map (
            O => \N__29046\,
            I => \N__29036\
        );

    \I__5117\ : InMux
    port map (
            O => \N__29045\,
            I => \N__29033\
        );

    \I__5116\ : Odrv12
    port map (
            O => \N__29042\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__5115\ : Odrv4
    port map (
            O => \N__29039\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__5114\ : LocalMux
    port map (
            O => \N__29036\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__5113\ : LocalMux
    port map (
            O => \N__29033\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__5112\ : CascadeMux
    port map (
            O => \N__29024\,
            I => \N__29020\
        );

    \I__5111\ : InMux
    port map (
            O => \N__29023\,
            I => \N__29017\
        );

    \I__5110\ : InMux
    port map (
            O => \N__29020\,
            I => \N__29014\
        );

    \I__5109\ : LocalMux
    port map (
            O => \N__29017\,
            I => \N__29011\
        );

    \I__5108\ : LocalMux
    port map (
            O => \N__29014\,
            I => \N__29008\
        );

    \I__5107\ : Span4Mux_h
    port map (
            O => \N__29011\,
            I => \N__29005\
        );

    \I__5106\ : Span12Mux_v
    port map (
            O => \N__29008\,
            I => \N__29002\
        );

    \I__5105\ : Odrv4
    port map (
            O => \N__29005\,
            I => \current_shift_inst.control_inputZ0Z_13\
        );

    \I__5104\ : Odrv12
    port map (
            O => \N__29002\,
            I => \current_shift_inst.control_inputZ0Z_13\
        );

    \I__5103\ : CascadeMux
    port map (
            O => \N__28997\,
            I => \N__28994\
        );

    \I__5102\ : InMux
    port map (
            O => \N__28994\,
            I => \N__28991\
        );

    \I__5101\ : LocalMux
    port map (
            O => \N__28991\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\
        );

    \I__5100\ : InMux
    port map (
            O => \N__28988\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\
        );

    \I__5099\ : InMux
    port map (
            O => \N__28985\,
            I => \N__28981\
        );

    \I__5098\ : InMux
    port map (
            O => \N__28984\,
            I => \N__28976\
        );

    \I__5097\ : LocalMux
    port map (
            O => \N__28981\,
            I => \N__28973\
        );

    \I__5096\ : InMux
    port map (
            O => \N__28980\,
            I => \N__28970\
        );

    \I__5095\ : InMux
    port map (
            O => \N__28979\,
            I => \N__28967\
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__28976\,
            I => \N__28964\
        );

    \I__5093\ : Odrv12
    port map (
            O => \N__28973\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__5092\ : LocalMux
    port map (
            O => \N__28970\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__5091\ : LocalMux
    port map (
            O => \N__28967\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__5090\ : Odrv4
    port map (
            O => \N__28964\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__5089\ : CascadeMux
    port map (
            O => \N__28955\,
            I => \N__28952\
        );

    \I__5088\ : InMux
    port map (
            O => \N__28952\,
            I => \N__28948\
        );

    \I__5087\ : InMux
    port map (
            O => \N__28951\,
            I => \N__28945\
        );

    \I__5086\ : LocalMux
    port map (
            O => \N__28948\,
            I => \N__28942\
        );

    \I__5085\ : LocalMux
    port map (
            O => \N__28945\,
            I => \N__28939\
        );

    \I__5084\ : Span4Mux_h
    port map (
            O => \N__28942\,
            I => \N__28936\
        );

    \I__5083\ : Span4Mux_v
    port map (
            O => \N__28939\,
            I => \N__28933\
        );

    \I__5082\ : Span4Mux_h
    port map (
            O => \N__28936\,
            I => \N__28930\
        );

    \I__5081\ : Odrv4
    port map (
            O => \N__28933\,
            I => \current_shift_inst.control_inputZ0Z_14\
        );

    \I__5080\ : Odrv4
    port map (
            O => \N__28930\,
            I => \current_shift_inst.control_inputZ0Z_14\
        );

    \I__5079\ : CascadeMux
    port map (
            O => \N__28925\,
            I => \N__28922\
        );

    \I__5078\ : InMux
    port map (
            O => \N__28922\,
            I => \N__28919\
        );

    \I__5077\ : LocalMux
    port map (
            O => \N__28919\,
            I => \N__28916\
        );

    \I__5076\ : Odrv4
    port map (
            O => \N__28916\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\
        );

    \I__5075\ : InMux
    port map (
            O => \N__28913\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\
        );

    \I__5074\ : CascadeMux
    port map (
            O => \N__28910\,
            I => \N__28907\
        );

    \I__5073\ : InMux
    port map (
            O => \N__28907\,
            I => \N__28903\
        );

    \I__5072\ : InMux
    port map (
            O => \N__28906\,
            I => \N__28898\
        );

    \I__5071\ : LocalMux
    port map (
            O => \N__28903\,
            I => \N__28895\
        );

    \I__5070\ : InMux
    port map (
            O => \N__28902\,
            I => \N__28892\
        );

    \I__5069\ : InMux
    port map (
            O => \N__28901\,
            I => \N__28889\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__28898\,
            I => \N__28886\
        );

    \I__5067\ : Odrv12
    port map (
            O => \N__28895\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__28892\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__5065\ : LocalMux
    port map (
            O => \N__28889\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__5064\ : Odrv4
    port map (
            O => \N__28886\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__5063\ : CascadeMux
    port map (
            O => \N__28877\,
            I => \N__28873\
        );

    \I__5062\ : InMux
    port map (
            O => \N__28876\,
            I => \N__28870\
        );

    \I__5061\ : InMux
    port map (
            O => \N__28873\,
            I => \N__28867\
        );

    \I__5060\ : LocalMux
    port map (
            O => \N__28870\,
            I => \N__28864\
        );

    \I__5059\ : LocalMux
    port map (
            O => \N__28867\,
            I => \N__28861\
        );

    \I__5058\ : Span4Mux_h
    port map (
            O => \N__28864\,
            I => \N__28856\
        );

    \I__5057\ : Span4Mux_h
    port map (
            O => \N__28861\,
            I => \N__28856\
        );

    \I__5056\ : Span4Mux_h
    port map (
            O => \N__28856\,
            I => \N__28853\
        );

    \I__5055\ : Odrv4
    port map (
            O => \N__28853\,
            I => \current_shift_inst.control_inputZ0Z_15\
        );

    \I__5054\ : InMux
    port map (
            O => \N__28850\,
            I => \N__28847\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__28847\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\
        );

    \I__5052\ : InMux
    port map (
            O => \N__28844\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\
        );

    \I__5051\ : CascadeMux
    port map (
            O => \N__28841\,
            I => \N__28838\
        );

    \I__5050\ : InMux
    port map (
            O => \N__28838\,
            I => \N__28834\
        );

    \I__5049\ : CascadeMux
    port map (
            O => \N__28837\,
            I => \N__28830\
        );

    \I__5048\ : LocalMux
    port map (
            O => \N__28834\,
            I => \N__28827\
        );

    \I__5047\ : InMux
    port map (
            O => \N__28833\,
            I => \N__28823\
        );

    \I__5046\ : InMux
    port map (
            O => \N__28830\,
            I => \N__28820\
        );

    \I__5045\ : Span4Mux_h
    port map (
            O => \N__28827\,
            I => \N__28817\
        );

    \I__5044\ : InMux
    port map (
            O => \N__28826\,
            I => \N__28814\
        );

    \I__5043\ : LocalMux
    port map (
            O => \N__28823\,
            I => \N__28809\
        );

    \I__5042\ : LocalMux
    port map (
            O => \N__28820\,
            I => \N__28809\
        );

    \I__5041\ : Span4Mux_h
    port map (
            O => \N__28817\,
            I => \N__28806\
        );

    \I__5040\ : LocalMux
    port map (
            O => \N__28814\,
            I => \N__28803\
        );

    \I__5039\ : Span4Mux_h
    port map (
            O => \N__28809\,
            I => \N__28800\
        );

    \I__5038\ : Odrv4
    port map (
            O => \N__28806\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__5037\ : Odrv12
    port map (
            O => \N__28803\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__5036\ : Odrv4
    port map (
            O => \N__28800\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__5035\ : CascadeMux
    port map (
            O => \N__28793\,
            I => \N__28789\
        );

    \I__5034\ : InMux
    port map (
            O => \N__28792\,
            I => \N__28786\
        );

    \I__5033\ : InMux
    port map (
            O => \N__28789\,
            I => \N__28783\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__28786\,
            I => \N__28780\
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__28783\,
            I => \N__28777\
        );

    \I__5030\ : Span4Mux_h
    port map (
            O => \N__28780\,
            I => \N__28774\
        );

    \I__5029\ : Span4Mux_h
    port map (
            O => \N__28777\,
            I => \N__28771\
        );

    \I__5028\ : Odrv4
    port map (
            O => \N__28774\,
            I => \current_shift_inst.control_inputZ0Z_16\
        );

    \I__5027\ : Odrv4
    port map (
            O => \N__28771\,
            I => \current_shift_inst.control_inputZ0Z_16\
        );

    \I__5026\ : CascadeMux
    port map (
            O => \N__28766\,
            I => \N__28763\
        );

    \I__5025\ : InMux
    port map (
            O => \N__28763\,
            I => \N__28760\
        );

    \I__5024\ : LocalMux
    port map (
            O => \N__28760\,
            I => \N__28757\
        );

    \I__5023\ : Odrv4
    port map (
            O => \N__28757\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\
        );

    \I__5022\ : InMux
    port map (
            O => \N__28754\,
            I => \bfn_11_12_0_\
        );

    \I__5021\ : InMux
    port map (
            O => \N__28751\,
            I => \N__28748\
        );

    \I__5020\ : LocalMux
    port map (
            O => \N__28748\,
            I => \N__28744\
        );

    \I__5019\ : InMux
    port map (
            O => \N__28747\,
            I => \N__28740\
        );

    \I__5018\ : Span4Mux_v
    port map (
            O => \N__28744\,
            I => \N__28737\
        );

    \I__5017\ : InMux
    port map (
            O => \N__28743\,
            I => \N__28733\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__28740\,
            I => \N__28730\
        );

    \I__5015\ : Span4Mux_h
    port map (
            O => \N__28737\,
            I => \N__28727\
        );

    \I__5014\ : InMux
    port map (
            O => \N__28736\,
            I => \N__28724\
        );

    \I__5013\ : LocalMux
    port map (
            O => \N__28733\,
            I => \N__28719\
        );

    \I__5012\ : Span4Mux_v
    port map (
            O => \N__28730\,
            I => \N__28719\
        );

    \I__5011\ : Odrv4
    port map (
            O => \N__28727\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__5010\ : LocalMux
    port map (
            O => \N__28724\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__5009\ : Odrv4
    port map (
            O => \N__28719\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__5008\ : CascadeMux
    port map (
            O => \N__28712\,
            I => \N__28709\
        );

    \I__5007\ : InMux
    port map (
            O => \N__28709\,
            I => \N__28705\
        );

    \I__5006\ : InMux
    port map (
            O => \N__28708\,
            I => \N__28702\
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__28705\,
            I => \N__28699\
        );

    \I__5004\ : LocalMux
    port map (
            O => \N__28702\,
            I => \N__28696\
        );

    \I__5003\ : Span4Mux_h
    port map (
            O => \N__28699\,
            I => \N__28693\
        );

    \I__5002\ : Odrv4
    port map (
            O => \N__28696\,
            I => \current_shift_inst.control_inputZ0Z_17\
        );

    \I__5001\ : Odrv4
    port map (
            O => \N__28693\,
            I => \current_shift_inst.control_inputZ0Z_17\
        );

    \I__5000\ : CascadeMux
    port map (
            O => \N__28688\,
            I => \N__28685\
        );

    \I__4999\ : InMux
    port map (
            O => \N__28685\,
            I => \N__28682\
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__28682\,
            I => \N__28679\
        );

    \I__4997\ : Span4Mux_h
    port map (
            O => \N__28679\,
            I => \N__28676\
        );

    \I__4996\ : Odrv4
    port map (
            O => \N__28676\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\
        );

    \I__4995\ : InMux
    port map (
            O => \N__28673\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\
        );

    \I__4994\ : InMux
    port map (
            O => \N__28670\,
            I => \N__28667\
        );

    \I__4993\ : LocalMux
    port map (
            O => \N__28667\,
            I => \N__28664\
        );

    \I__4992\ : Span4Mux_h
    port map (
            O => \N__28664\,
            I => \N__28660\
        );

    \I__4991\ : InMux
    port map (
            O => \N__28663\,
            I => \N__28656\
        );

    \I__4990\ : Span4Mux_h
    port map (
            O => \N__28660\,
            I => \N__28652\
        );

    \I__4989\ : InMux
    port map (
            O => \N__28659\,
            I => \N__28649\
        );

    \I__4988\ : LocalMux
    port map (
            O => \N__28656\,
            I => \N__28646\
        );

    \I__4987\ : InMux
    port map (
            O => \N__28655\,
            I => \N__28643\
        );

    \I__4986\ : Odrv4
    port map (
            O => \N__28652\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__4985\ : LocalMux
    port map (
            O => \N__28649\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__4984\ : Odrv4
    port map (
            O => \N__28646\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__28643\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__4982\ : CascadeMux
    port map (
            O => \N__28634\,
            I => \N__28630\
        );

    \I__4981\ : InMux
    port map (
            O => \N__28633\,
            I => \N__28627\
        );

    \I__4980\ : InMux
    port map (
            O => \N__28630\,
            I => \N__28624\
        );

    \I__4979\ : LocalMux
    port map (
            O => \N__28627\,
            I => \N__28621\
        );

    \I__4978\ : LocalMux
    port map (
            O => \N__28624\,
            I => \N__28618\
        );

    \I__4977\ : Span4Mux_h
    port map (
            O => \N__28621\,
            I => \N__28615\
        );

    \I__4976\ : Span4Mux_h
    port map (
            O => \N__28618\,
            I => \N__28612\
        );

    \I__4975\ : Odrv4
    port map (
            O => \N__28615\,
            I => \current_shift_inst.control_inputZ0Z_18\
        );

    \I__4974\ : Odrv4
    port map (
            O => \N__28612\,
            I => \current_shift_inst.control_inputZ0Z_18\
        );

    \I__4973\ : CascadeMux
    port map (
            O => \N__28607\,
            I => \N__28604\
        );

    \I__4972\ : InMux
    port map (
            O => \N__28604\,
            I => \N__28601\
        );

    \I__4971\ : LocalMux
    port map (
            O => \N__28601\,
            I => \N__28598\
        );

    \I__4970\ : Odrv4
    port map (
            O => \N__28598\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\
        );

    \I__4969\ : InMux
    port map (
            O => \N__28595\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\
        );

    \I__4968\ : InMux
    port map (
            O => \N__28592\,
            I => \N__28587\
        );

    \I__4967\ : InMux
    port map (
            O => \N__28591\,
            I => \N__28584\
        );

    \I__4966\ : InMux
    port map (
            O => \N__28590\,
            I => \N__28580\
        );

    \I__4965\ : LocalMux
    port map (
            O => \N__28587\,
            I => \N__28577\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__28584\,
            I => \N__28574\
        );

    \I__4963\ : InMux
    port map (
            O => \N__28583\,
            I => \N__28571\
        );

    \I__4962\ : LocalMux
    port map (
            O => \N__28580\,
            I => \N__28568\
        );

    \I__4961\ : Span4Mux_h
    port map (
            O => \N__28577\,
            I => \N__28563\
        );

    \I__4960\ : Span4Mux_h
    port map (
            O => \N__28574\,
            I => \N__28563\
        );

    \I__4959\ : LocalMux
    port map (
            O => \N__28571\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__4958\ : Odrv4
    port map (
            O => \N__28568\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__4957\ : Odrv4
    port map (
            O => \N__28563\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__4956\ : CascadeMux
    port map (
            O => \N__28556\,
            I => \N__28552\
        );

    \I__4955\ : InMux
    port map (
            O => \N__28555\,
            I => \N__28549\
        );

    \I__4954\ : InMux
    port map (
            O => \N__28552\,
            I => \N__28546\
        );

    \I__4953\ : LocalMux
    port map (
            O => \N__28549\,
            I => \N__28543\
        );

    \I__4952\ : LocalMux
    port map (
            O => \N__28546\,
            I => \N__28540\
        );

    \I__4951\ : Span4Mux_v
    port map (
            O => \N__28543\,
            I => \N__28537\
        );

    \I__4950\ : Span4Mux_h
    port map (
            O => \N__28540\,
            I => \N__28534\
        );

    \I__4949\ : Odrv4
    port map (
            O => \N__28537\,
            I => \current_shift_inst.control_inputZ0Z_19\
        );

    \I__4948\ : Odrv4
    port map (
            O => \N__28534\,
            I => \current_shift_inst.control_inputZ0Z_19\
        );

    \I__4947\ : InMux
    port map (
            O => \N__28529\,
            I => \N__28526\
        );

    \I__4946\ : LocalMux
    port map (
            O => \N__28526\,
            I => \N__28523\
        );

    \I__4945\ : Odrv12
    port map (
            O => \N__28523\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\
        );

    \I__4944\ : InMux
    port map (
            O => \N__28520\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\
        );

    \I__4943\ : InMux
    port map (
            O => \N__28517\,
            I => \N__28514\
        );

    \I__4942\ : LocalMux
    port map (
            O => \N__28514\,
            I => \N__28511\
        );

    \I__4941\ : Span4Mux_h
    port map (
            O => \N__28511\,
            I => \N__28506\
        );

    \I__4940\ : InMux
    port map (
            O => \N__28510\,
            I => \N__28500\
        );

    \I__4939\ : InMux
    port map (
            O => \N__28509\,
            I => \N__28500\
        );

    \I__4938\ : Span4Mux_h
    port map (
            O => \N__28506\,
            I => \N__28497\
        );

    \I__4937\ : InMux
    port map (
            O => \N__28505\,
            I => \N__28494\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__28500\,
            I => \N__28491\
        );

    \I__4935\ : Odrv4
    port map (
            O => \N__28497\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__4934\ : LocalMux
    port map (
            O => \N__28494\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__4933\ : Odrv4
    port map (
            O => \N__28491\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__4932\ : CascadeMux
    port map (
            O => \N__28484\,
            I => \N__28480\
        );

    \I__4931\ : InMux
    port map (
            O => \N__28483\,
            I => \N__28477\
        );

    \I__4930\ : InMux
    port map (
            O => \N__28480\,
            I => \N__28474\
        );

    \I__4929\ : LocalMux
    port map (
            O => \N__28477\,
            I => \N__28471\
        );

    \I__4928\ : LocalMux
    port map (
            O => \N__28474\,
            I => \N__28468\
        );

    \I__4927\ : Span12Mux_v
    port map (
            O => \N__28471\,
            I => \N__28465\
        );

    \I__4926\ : Span4Mux_h
    port map (
            O => \N__28468\,
            I => \N__28462\
        );

    \I__4925\ : Odrv12
    port map (
            O => \N__28465\,
            I => \current_shift_inst.control_inputZ0Z_6\
        );

    \I__4924\ : Odrv4
    port map (
            O => \N__28462\,
            I => \current_shift_inst.control_inputZ0Z_6\
        );

    \I__4923\ : InMux
    port map (
            O => \N__28457\,
            I => \N__28454\
        );

    \I__4922\ : LocalMux
    port map (
            O => \N__28454\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\
        );

    \I__4921\ : InMux
    port map (
            O => \N__28451\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\
        );

    \I__4920\ : CascadeMux
    port map (
            O => \N__28448\,
            I => \N__28445\
        );

    \I__4919\ : InMux
    port map (
            O => \N__28445\,
            I => \N__28442\
        );

    \I__4918\ : LocalMux
    port map (
            O => \N__28442\,
            I => \N__28437\
        );

    \I__4917\ : InMux
    port map (
            O => \N__28441\,
            I => \N__28434\
        );

    \I__4916\ : InMux
    port map (
            O => \N__28440\,
            I => \N__28431\
        );

    \I__4915\ : Span4Mux_v
    port map (
            O => \N__28437\,
            I => \N__28424\
        );

    \I__4914\ : LocalMux
    port map (
            O => \N__28434\,
            I => \N__28424\
        );

    \I__4913\ : LocalMux
    port map (
            O => \N__28431\,
            I => \N__28424\
        );

    \I__4912\ : Span4Mux_h
    port map (
            O => \N__28424\,
            I => \N__28420\
        );

    \I__4911\ : InMux
    port map (
            O => \N__28423\,
            I => \N__28417\
        );

    \I__4910\ : Odrv4
    port map (
            O => \N__28420\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__4909\ : LocalMux
    port map (
            O => \N__28417\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__4908\ : InMux
    port map (
            O => \N__28412\,
            I => \N__28408\
        );

    \I__4907\ : CascadeMux
    port map (
            O => \N__28411\,
            I => \N__28405\
        );

    \I__4906\ : LocalMux
    port map (
            O => \N__28408\,
            I => \N__28402\
        );

    \I__4905\ : InMux
    port map (
            O => \N__28405\,
            I => \N__28399\
        );

    \I__4904\ : Span4Mux_h
    port map (
            O => \N__28402\,
            I => \N__28396\
        );

    \I__4903\ : LocalMux
    port map (
            O => \N__28399\,
            I => \N__28393\
        );

    \I__4902\ : Span4Mux_v
    port map (
            O => \N__28396\,
            I => \N__28388\
        );

    \I__4901\ : Span4Mux_v
    port map (
            O => \N__28393\,
            I => \N__28388\
        );

    \I__4900\ : Odrv4
    port map (
            O => \N__28388\,
            I => \current_shift_inst.control_inputZ0Z_7\
        );

    \I__4899\ : CascadeMux
    port map (
            O => \N__28385\,
            I => \N__28382\
        );

    \I__4898\ : InMux
    port map (
            O => \N__28382\,
            I => \N__28379\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__28379\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\
        );

    \I__4896\ : InMux
    port map (
            O => \N__28376\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\
        );

    \I__4895\ : InMux
    port map (
            O => \N__28373\,
            I => \N__28370\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__28370\,
            I => \N__28367\
        );

    \I__4893\ : Span4Mux_h
    port map (
            O => \N__28367\,
            I => \N__28362\
        );

    \I__4892\ : InMux
    port map (
            O => \N__28366\,
            I => \N__28356\
        );

    \I__4891\ : InMux
    port map (
            O => \N__28365\,
            I => \N__28356\
        );

    \I__4890\ : Span4Mux_h
    port map (
            O => \N__28362\,
            I => \N__28353\
        );

    \I__4889\ : InMux
    port map (
            O => \N__28361\,
            I => \N__28350\
        );

    \I__4888\ : LocalMux
    port map (
            O => \N__28356\,
            I => \N__28347\
        );

    \I__4887\ : Odrv4
    port map (
            O => \N__28353\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__4886\ : LocalMux
    port map (
            O => \N__28350\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__4885\ : Odrv4
    port map (
            O => \N__28347\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__4884\ : CascadeMux
    port map (
            O => \N__28340\,
            I => \N__28336\
        );

    \I__4883\ : InMux
    port map (
            O => \N__28339\,
            I => \N__28333\
        );

    \I__4882\ : InMux
    port map (
            O => \N__28336\,
            I => \N__28330\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__28333\,
            I => \N__28327\
        );

    \I__4880\ : LocalMux
    port map (
            O => \N__28330\,
            I => \N__28324\
        );

    \I__4879\ : Span4Mux_h
    port map (
            O => \N__28327\,
            I => \N__28319\
        );

    \I__4878\ : Span4Mux_h
    port map (
            O => \N__28324\,
            I => \N__28319\
        );

    \I__4877\ : Odrv4
    port map (
            O => \N__28319\,
            I => \current_shift_inst.control_inputZ0Z_8\
        );

    \I__4876\ : InMux
    port map (
            O => \N__28316\,
            I => \N__28313\
        );

    \I__4875\ : LocalMux
    port map (
            O => \N__28313\,
            I => \N__28310\
        );

    \I__4874\ : Odrv4
    port map (
            O => \N__28310\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\
        );

    \I__4873\ : InMux
    port map (
            O => \N__28307\,
            I => \bfn_11_11_0_\
        );

    \I__4872\ : CascadeMux
    port map (
            O => \N__28304\,
            I => \N__28300\
        );

    \I__4871\ : InMux
    port map (
            O => \N__28303\,
            I => \N__28297\
        );

    \I__4870\ : InMux
    port map (
            O => \N__28300\,
            I => \N__28293\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__28297\,
            I => \N__28290\
        );

    \I__4868\ : CascadeMux
    port map (
            O => \N__28296\,
            I => \N__28287\
        );

    \I__4867\ : LocalMux
    port map (
            O => \N__28293\,
            I => \N__28281\
        );

    \I__4866\ : Span4Mux_v
    port map (
            O => \N__28290\,
            I => \N__28281\
        );

    \I__4865\ : InMux
    port map (
            O => \N__28287\,
            I => \N__28278\
        );

    \I__4864\ : InMux
    port map (
            O => \N__28286\,
            I => \N__28275\
        );

    \I__4863\ : Sp12to4
    port map (
            O => \N__28281\,
            I => \N__28270\
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__28278\,
            I => \N__28270\
        );

    \I__4861\ : LocalMux
    port map (
            O => \N__28275\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__4860\ : Odrv12
    port map (
            O => \N__28270\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__4859\ : InMux
    port map (
            O => \N__28265\,
            I => \N__28262\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__28262\,
            I => \N__28258\
        );

    \I__4857\ : CascadeMux
    port map (
            O => \N__28261\,
            I => \N__28255\
        );

    \I__4856\ : Span4Mux_v
    port map (
            O => \N__28258\,
            I => \N__28252\
        );

    \I__4855\ : InMux
    port map (
            O => \N__28255\,
            I => \N__28249\
        );

    \I__4854\ : Span4Mux_v
    port map (
            O => \N__28252\,
            I => \N__28246\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__28249\,
            I => \N__28243\
        );

    \I__4852\ : Span4Mux_h
    port map (
            O => \N__28246\,
            I => \N__28240\
        );

    \I__4851\ : Span4Mux_h
    port map (
            O => \N__28243\,
            I => \N__28237\
        );

    \I__4850\ : Odrv4
    port map (
            O => \N__28240\,
            I => \current_shift_inst.control_inputZ0Z_9\
        );

    \I__4849\ : Odrv4
    port map (
            O => \N__28237\,
            I => \current_shift_inst.control_inputZ0Z_9\
        );

    \I__4848\ : CascadeMux
    port map (
            O => \N__28232\,
            I => \N__28229\
        );

    \I__4847\ : InMux
    port map (
            O => \N__28229\,
            I => \N__28226\
        );

    \I__4846\ : LocalMux
    port map (
            O => \N__28226\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\
        );

    \I__4845\ : InMux
    port map (
            O => \N__28223\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\
        );

    \I__4844\ : InMux
    port map (
            O => \N__28220\,
            I => \N__28216\
        );

    \I__4843\ : CascadeMux
    port map (
            O => \N__28219\,
            I => \N__28213\
        );

    \I__4842\ : LocalMux
    port map (
            O => \N__28216\,
            I => \N__28209\
        );

    \I__4841\ : InMux
    port map (
            O => \N__28213\,
            I => \N__28206\
        );

    \I__4840\ : InMux
    port map (
            O => \N__28212\,
            I => \N__28203\
        );

    \I__4839\ : Span4Mux_h
    port map (
            O => \N__28209\,
            I => \N__28196\
        );

    \I__4838\ : LocalMux
    port map (
            O => \N__28206\,
            I => \N__28196\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__28203\,
            I => \N__28196\
        );

    \I__4836\ : Span4Mux_h
    port map (
            O => \N__28196\,
            I => \N__28192\
        );

    \I__4835\ : InMux
    port map (
            O => \N__28195\,
            I => \N__28189\
        );

    \I__4834\ : Odrv4
    port map (
            O => \N__28192\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__4833\ : LocalMux
    port map (
            O => \N__28189\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__4832\ : InMux
    port map (
            O => \N__28184\,
            I => \N__28180\
        );

    \I__4831\ : CascadeMux
    port map (
            O => \N__28183\,
            I => \N__28177\
        );

    \I__4830\ : LocalMux
    port map (
            O => \N__28180\,
            I => \N__28174\
        );

    \I__4829\ : InMux
    port map (
            O => \N__28177\,
            I => \N__28171\
        );

    \I__4828\ : Span4Mux_v
    port map (
            O => \N__28174\,
            I => \N__28168\
        );

    \I__4827\ : LocalMux
    port map (
            O => \N__28171\,
            I => \N__28165\
        );

    \I__4826\ : Span4Mux_h
    port map (
            O => \N__28168\,
            I => \N__28160\
        );

    \I__4825\ : Span4Mux_h
    port map (
            O => \N__28165\,
            I => \N__28160\
        );

    \I__4824\ : Odrv4
    port map (
            O => \N__28160\,
            I => \current_shift_inst.control_inputZ0Z_10\
        );

    \I__4823\ : CascadeMux
    port map (
            O => \N__28157\,
            I => \N__28154\
        );

    \I__4822\ : InMux
    port map (
            O => \N__28154\,
            I => \N__28151\
        );

    \I__4821\ : LocalMux
    port map (
            O => \N__28151\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\
        );

    \I__4820\ : InMux
    port map (
            O => \N__28148\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\
        );

    \I__4819\ : InMux
    port map (
            O => \N__28145\,
            I => \N__28141\
        );

    \I__4818\ : InMux
    port map (
            O => \N__28144\,
            I => \N__28138\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__28141\,
            I => \N__28135\
        );

    \I__4816\ : LocalMux
    port map (
            O => \N__28138\,
            I => \N__28130\
        );

    \I__4815\ : Span12Mux_s10_v
    port map (
            O => \N__28135\,
            I => \N__28127\
        );

    \I__4814\ : InMux
    port map (
            O => \N__28134\,
            I => \N__28124\
        );

    \I__4813\ : InMux
    port map (
            O => \N__28133\,
            I => \N__28121\
        );

    \I__4812\ : Span4Mux_v
    port map (
            O => \N__28130\,
            I => \N__28118\
        );

    \I__4811\ : Odrv12
    port map (
            O => \N__28127\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__4810\ : LocalMux
    port map (
            O => \N__28124\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__4809\ : LocalMux
    port map (
            O => \N__28121\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__4808\ : Odrv4
    port map (
            O => \N__28118\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__4807\ : CascadeMux
    port map (
            O => \N__28109\,
            I => \N__28105\
        );

    \I__4806\ : InMux
    port map (
            O => \N__28108\,
            I => \N__28102\
        );

    \I__4805\ : InMux
    port map (
            O => \N__28105\,
            I => \N__28099\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__28102\,
            I => \N__28096\
        );

    \I__4803\ : LocalMux
    port map (
            O => \N__28099\,
            I => \N__28093\
        );

    \I__4802\ : Span4Mux_v
    port map (
            O => \N__28096\,
            I => \N__28090\
        );

    \I__4801\ : Span4Mux_h
    port map (
            O => \N__28093\,
            I => \N__28087\
        );

    \I__4800\ : Odrv4
    port map (
            O => \N__28090\,
            I => \current_shift_inst.control_inputZ0Z_11\
        );

    \I__4799\ : Odrv4
    port map (
            O => \N__28087\,
            I => \current_shift_inst.control_inputZ0Z_11\
        );

    \I__4798\ : CascadeMux
    port map (
            O => \N__28082\,
            I => \N__28079\
        );

    \I__4797\ : InMux
    port map (
            O => \N__28079\,
            I => \N__28076\
        );

    \I__4796\ : LocalMux
    port map (
            O => \N__28076\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\
        );

    \I__4795\ : InMux
    port map (
            O => \N__28073\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\
        );

    \I__4794\ : InMux
    port map (
            O => \N__28070\,
            I => \N__28066\
        );

    \I__4793\ : CascadeMux
    port map (
            O => \N__28069\,
            I => \N__28063\
        );

    \I__4792\ : LocalMux
    port map (
            O => \N__28066\,
            I => \N__28060\
        );

    \I__4791\ : InMux
    port map (
            O => \N__28063\,
            I => \N__28057\
        );

    \I__4790\ : Span4Mux_h
    port map (
            O => \N__28060\,
            I => \N__28051\
        );

    \I__4789\ : LocalMux
    port map (
            O => \N__28057\,
            I => \N__28051\
        );

    \I__4788\ : InMux
    port map (
            O => \N__28056\,
            I => \N__28047\
        );

    \I__4787\ : Span4Mux_h
    port map (
            O => \N__28051\,
            I => \N__28044\
        );

    \I__4786\ : InMux
    port map (
            O => \N__28050\,
            I => \N__28041\
        );

    \I__4785\ : LocalMux
    port map (
            O => \N__28047\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__4784\ : Odrv4
    port map (
            O => \N__28044\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__28041\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__4782\ : CascadeMux
    port map (
            O => \N__28034\,
            I => \N__28031\
        );

    \I__4781\ : InMux
    port map (
            O => \N__28031\,
            I => \N__28027\
        );

    \I__4780\ : InMux
    port map (
            O => \N__28030\,
            I => \N__28024\
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__28027\,
            I => \N__28021\
        );

    \I__4778\ : LocalMux
    port map (
            O => \N__28024\,
            I => \N__28018\
        );

    \I__4777\ : Span4Mux_v
    port map (
            O => \N__28021\,
            I => \N__28015\
        );

    \I__4776\ : Span4Mux_h
    port map (
            O => \N__28018\,
            I => \N__28012\
        );

    \I__4775\ : Span4Mux_h
    port map (
            O => \N__28015\,
            I => \N__28009\
        );

    \I__4774\ : Odrv4
    port map (
            O => \N__28012\,
            I => \current_shift_inst.control_inputZ0Z_12\
        );

    \I__4773\ : Odrv4
    port map (
            O => \N__28009\,
            I => \current_shift_inst.control_inputZ0Z_12\
        );

    \I__4772\ : InMux
    port map (
            O => \N__28004\,
            I => \N__28001\
        );

    \I__4771\ : LocalMux
    port map (
            O => \N__28001\,
            I => \N__27998\
        );

    \I__4770\ : Odrv4
    port map (
            O => \N__27998\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\
        );

    \I__4769\ : InMux
    port map (
            O => \N__27995\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\
        );

    \I__4768\ : InMux
    port map (
            O => \N__27992\,
            I => \N__27988\
        );

    \I__4767\ : InMux
    port map (
            O => \N__27991\,
            I => \N__27985\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__27988\,
            I => \N__27981\
        );

    \I__4765\ : LocalMux
    port map (
            O => \N__27985\,
            I => \N__27978\
        );

    \I__4764\ : InMux
    port map (
            O => \N__27984\,
            I => \N__27975\
        );

    \I__4763\ : Span4Mux_v
    port map (
            O => \N__27981\,
            I => \N__27972\
        );

    \I__4762\ : Odrv12
    port map (
            O => \N__27978\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_0\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__27975\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_0\
        );

    \I__4760\ : Odrv4
    port map (
            O => \N__27972\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_0\
        );

    \I__4759\ : InMux
    port map (
            O => \N__27965\,
            I => \N__27961\
        );

    \I__4758\ : CascadeMux
    port map (
            O => \N__27964\,
            I => \N__27958\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__27961\,
            I => \N__27955\
        );

    \I__4756\ : InMux
    port map (
            O => \N__27958\,
            I => \N__27952\
        );

    \I__4755\ : Span4Mux_v
    port map (
            O => \N__27955\,
            I => \N__27949\
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__27952\,
            I => \N__27946\
        );

    \I__4753\ : Span4Mux_h
    port map (
            O => \N__27949\,
            I => \N__27941\
        );

    \I__4752\ : Span4Mux_h
    port map (
            O => \N__27946\,
            I => \N__27941\
        );

    \I__4751\ : Odrv4
    port map (
            O => \N__27941\,
            I => \current_shift_inst.control_inputZ0Z_0\
        );

    \I__4750\ : CascadeMux
    port map (
            O => \N__27938\,
            I => \N__27935\
        );

    \I__4749\ : InMux
    port map (
            O => \N__27935\,
            I => \N__27932\
        );

    \I__4748\ : LocalMux
    port map (
            O => \N__27932\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_axb_0\
        );

    \I__4747\ : InMux
    port map (
            O => \N__27929\,
            I => \N__27926\
        );

    \I__4746\ : LocalMux
    port map (
            O => \N__27926\,
            I => \N__27923\
        );

    \I__4745\ : Span4Mux_h
    port map (
            O => \N__27923\,
            I => \N__27919\
        );

    \I__4744\ : InMux
    port map (
            O => \N__27922\,
            I => \N__27915\
        );

    \I__4743\ : Span4Mux_h
    port map (
            O => \N__27919\,
            I => \N__27912\
        );

    \I__4742\ : InMux
    port map (
            O => \N__27918\,
            I => \N__27909\
        );

    \I__4741\ : LocalMux
    port map (
            O => \N__27915\,
            I => \N__27906\
        );

    \I__4740\ : Odrv4
    port map (
            O => \N__27912\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__4739\ : LocalMux
    port map (
            O => \N__27909\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__4738\ : Odrv4
    port map (
            O => \N__27906\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__4737\ : CascadeMux
    port map (
            O => \N__27899\,
            I => \N__27896\
        );

    \I__4736\ : InMux
    port map (
            O => \N__27896\,
            I => \N__27892\
        );

    \I__4735\ : InMux
    port map (
            O => \N__27895\,
            I => \N__27889\
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__27892\,
            I => \N__27886\
        );

    \I__4733\ : LocalMux
    port map (
            O => \N__27889\,
            I => \N__27883\
        );

    \I__4732\ : Span4Mux_h
    port map (
            O => \N__27886\,
            I => \N__27880\
        );

    \I__4731\ : Odrv4
    port map (
            O => \N__27883\,
            I => \current_shift_inst.control_inputZ0Z_1\
        );

    \I__4730\ : Odrv4
    port map (
            O => \N__27880\,
            I => \current_shift_inst.control_inputZ0Z_1\
        );

    \I__4729\ : CascadeMux
    port map (
            O => \N__27875\,
            I => \N__27872\
        );

    \I__4728\ : InMux
    port map (
            O => \N__27872\,
            I => \N__27869\
        );

    \I__4727\ : LocalMux
    port map (
            O => \N__27869\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1\
        );

    \I__4726\ : InMux
    port map (
            O => \N__27866\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_0\
        );

    \I__4725\ : CascadeMux
    port map (
            O => \N__27863\,
            I => \N__27860\
        );

    \I__4724\ : InMux
    port map (
            O => \N__27860\,
            I => \N__27856\
        );

    \I__4723\ : InMux
    port map (
            O => \N__27859\,
            I => \N__27853\
        );

    \I__4722\ : LocalMux
    port map (
            O => \N__27856\,
            I => \N__27850\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__27853\,
            I => \N__27847\
        );

    \I__4720\ : Span4Mux_h
    port map (
            O => \N__27850\,
            I => \N__27844\
        );

    \I__4719\ : Odrv4
    port map (
            O => \N__27847\,
            I => \current_shift_inst.control_inputZ0Z_2\
        );

    \I__4718\ : Odrv4
    port map (
            O => \N__27844\,
            I => \current_shift_inst.control_inputZ0Z_2\
        );

    \I__4717\ : InMux
    port map (
            O => \N__27839\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\
        );

    \I__4716\ : InMux
    port map (
            O => \N__27836\,
            I => \N__27833\
        );

    \I__4715\ : LocalMux
    port map (
            O => \N__27833\,
            I => \N__27829\
        );

    \I__4714\ : InMux
    port map (
            O => \N__27832\,
            I => \N__27826\
        );

    \I__4713\ : Span4Mux_v
    port map (
            O => \N__27829\,
            I => \N__27823\
        );

    \I__4712\ : LocalMux
    port map (
            O => \N__27826\,
            I => \N__27820\
        );

    \I__4711\ : Span4Mux_h
    port map (
            O => \N__27823\,
            I => \N__27817\
        );

    \I__4710\ : Span4Mux_h
    port map (
            O => \N__27820\,
            I => \N__27814\
        );

    \I__4709\ : Odrv4
    port map (
            O => \N__27817\,
            I => \current_shift_inst.control_inputZ0Z_3\
        );

    \I__4708\ : Odrv4
    port map (
            O => \N__27814\,
            I => \current_shift_inst.control_inputZ0Z_3\
        );

    \I__4707\ : InMux
    port map (
            O => \N__27809\,
            I => \N__27806\
        );

    \I__4706\ : LocalMux
    port map (
            O => \N__27806\,
            I => \N__27800\
        );

    \I__4705\ : InMux
    port map (
            O => \N__27805\,
            I => \N__27797\
        );

    \I__4704\ : InMux
    port map (
            O => \N__27804\,
            I => \N__27794\
        );

    \I__4703\ : CascadeMux
    port map (
            O => \N__27803\,
            I => \N__27791\
        );

    \I__4702\ : Span4Mux_v
    port map (
            O => \N__27800\,
            I => \N__27784\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__27797\,
            I => \N__27784\
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__27794\,
            I => \N__27784\
        );

    \I__4699\ : InMux
    port map (
            O => \N__27791\,
            I => \N__27781\
        );

    \I__4698\ : Span4Mux_h
    port map (
            O => \N__27784\,
            I => \N__27778\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__27781\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__4696\ : Odrv4
    port map (
            O => \N__27778\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__4695\ : CascadeMux
    port map (
            O => \N__27773\,
            I => \N__27770\
        );

    \I__4694\ : InMux
    port map (
            O => \N__27770\,
            I => \N__27767\
        );

    \I__4693\ : LocalMux
    port map (
            O => \N__27767\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\
        );

    \I__4692\ : InMux
    port map (
            O => \N__27764\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\
        );

    \I__4691\ : InMux
    port map (
            O => \N__27761\,
            I => \N__27755\
        );

    \I__4690\ : InMux
    port map (
            O => \N__27760\,
            I => \N__27755\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__27755\,
            I => \N__27751\
        );

    \I__4688\ : InMux
    port map (
            O => \N__27754\,
            I => \N__27748\
        );

    \I__4687\ : Span4Mux_v
    port map (
            O => \N__27751\,
            I => \N__27745\
        );

    \I__4686\ : LocalMux
    port map (
            O => \N__27748\,
            I => \N__27741\
        );

    \I__4685\ : Span4Mux_h
    port map (
            O => \N__27745\,
            I => \N__27738\
        );

    \I__4684\ : InMux
    port map (
            O => \N__27744\,
            I => \N__27735\
        );

    \I__4683\ : Odrv12
    port map (
            O => \N__27741\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__4682\ : Odrv4
    port map (
            O => \N__27738\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__27735\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__4680\ : CascadeMux
    port map (
            O => \N__27728\,
            I => \N__27725\
        );

    \I__4679\ : InMux
    port map (
            O => \N__27725\,
            I => \N__27722\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__27722\,
            I => \N__27718\
        );

    \I__4677\ : InMux
    port map (
            O => \N__27721\,
            I => \N__27715\
        );

    \I__4676\ : Span4Mux_v
    port map (
            O => \N__27718\,
            I => \N__27712\
        );

    \I__4675\ : LocalMux
    port map (
            O => \N__27715\,
            I => \N__27707\
        );

    \I__4674\ : Span4Mux_h
    port map (
            O => \N__27712\,
            I => \N__27707\
        );

    \I__4673\ : Odrv4
    port map (
            O => \N__27707\,
            I => \current_shift_inst.control_inputZ0Z_4\
        );

    \I__4672\ : CascadeMux
    port map (
            O => \N__27704\,
            I => \N__27701\
        );

    \I__4671\ : InMux
    port map (
            O => \N__27701\,
            I => \N__27698\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__27698\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\
        );

    \I__4669\ : InMux
    port map (
            O => \N__27695\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\
        );

    \I__4668\ : InMux
    port map (
            O => \N__27692\,
            I => \N__27687\
        );

    \I__4667\ : InMux
    port map (
            O => \N__27691\,
            I => \N__27684\
        );

    \I__4666\ : InMux
    port map (
            O => \N__27690\,
            I => \N__27681\
        );

    \I__4665\ : LocalMux
    port map (
            O => \N__27687\,
            I => \N__27678\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__27684\,
            I => \N__27672\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__27681\,
            I => \N__27672\
        );

    \I__4662\ : Span4Mux_h
    port map (
            O => \N__27678\,
            I => \N__27669\
        );

    \I__4661\ : InMux
    port map (
            O => \N__27677\,
            I => \N__27666\
        );

    \I__4660\ : Span4Mux_h
    port map (
            O => \N__27672\,
            I => \N__27663\
        );

    \I__4659\ : Odrv4
    port map (
            O => \N__27669\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__27666\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__4657\ : Odrv4
    port map (
            O => \N__27663\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__4656\ : InMux
    port map (
            O => \N__27656\,
            I => \N__27652\
        );

    \I__4655\ : CascadeMux
    port map (
            O => \N__27655\,
            I => \N__27649\
        );

    \I__4654\ : LocalMux
    port map (
            O => \N__27652\,
            I => \N__27646\
        );

    \I__4653\ : InMux
    port map (
            O => \N__27649\,
            I => \N__27643\
        );

    \I__4652\ : Span4Mux_h
    port map (
            O => \N__27646\,
            I => \N__27640\
        );

    \I__4651\ : LocalMux
    port map (
            O => \N__27643\,
            I => \N__27637\
        );

    \I__4650\ : Span4Mux_h
    port map (
            O => \N__27640\,
            I => \N__27634\
        );

    \I__4649\ : Span12Mux_v
    port map (
            O => \N__27637\,
            I => \N__27631\
        );

    \I__4648\ : Odrv4
    port map (
            O => \N__27634\,
            I => \current_shift_inst.control_inputZ0Z_5\
        );

    \I__4647\ : Odrv12
    port map (
            O => \N__27631\,
            I => \current_shift_inst.control_inputZ0Z_5\
        );

    \I__4646\ : CascadeMux
    port map (
            O => \N__27626\,
            I => \N__27623\
        );

    \I__4645\ : InMux
    port map (
            O => \N__27623\,
            I => \N__27620\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__27620\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\
        );

    \I__4643\ : InMux
    port map (
            O => \N__27617\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\
        );

    \I__4642\ : CascadeMux
    port map (
            O => \N__27614\,
            I => \N__27609\
        );

    \I__4641\ : CascadeMux
    port map (
            O => \N__27613\,
            I => \N__27606\
        );

    \I__4640\ : CascadeMux
    port map (
            O => \N__27612\,
            I => \N__27603\
        );

    \I__4639\ : InMux
    port map (
            O => \N__27609\,
            I => \N__27598\
        );

    \I__4638\ : InMux
    port map (
            O => \N__27606\,
            I => \N__27595\
        );

    \I__4637\ : InMux
    port map (
            O => \N__27603\,
            I => \N__27590\
        );

    \I__4636\ : InMux
    port map (
            O => \N__27602\,
            I => \N__27590\
        );

    \I__4635\ : InMux
    port map (
            O => \N__27601\,
            I => \N__27587\
        );

    \I__4634\ : LocalMux
    port map (
            O => \N__27598\,
            I => \N__27584\
        );

    \I__4633\ : LocalMux
    port map (
            O => \N__27595\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__4632\ : LocalMux
    port map (
            O => \N__27590\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__27587\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__4630\ : Odrv12
    port map (
            O => \N__27584\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__4629\ : InMux
    port map (
            O => \N__27575\,
            I => \N__27572\
        );

    \I__4628\ : LocalMux
    port map (
            O => \N__27572\,
            I => \N__27569\
        );

    \I__4627\ : Span4Mux_h
    port map (
            O => \N__27569\,
            I => \N__27564\
        );

    \I__4626\ : InMux
    port map (
            O => \N__27568\,
            I => \N__27560\
        );

    \I__4625\ : InMux
    port map (
            O => \N__27567\,
            I => \N__27557\
        );

    \I__4624\ : Sp12to4
    port map (
            O => \N__27564\,
            I => \N__27554\
        );

    \I__4623\ : InMux
    port map (
            O => \N__27563\,
            I => \N__27551\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__27560\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__27557\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__4620\ : Odrv12
    port map (
            O => \N__27554\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__4619\ : LocalMux
    port map (
            O => \N__27551\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__4618\ : InMux
    port map (
            O => \N__27542\,
            I => \N__27536\
        );

    \I__4617\ : InMux
    port map (
            O => \N__27541\,
            I => \N__27533\
        );

    \I__4616\ : InMux
    port map (
            O => \N__27540\,
            I => \N__27530\
        );

    \I__4615\ : InMux
    port map (
            O => \N__27539\,
            I => \N__27527\
        );

    \I__4614\ : LocalMux
    port map (
            O => \N__27536\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__4613\ : LocalMux
    port map (
            O => \N__27533\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__4612\ : LocalMux
    port map (
            O => \N__27530\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__27527\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__4610\ : CEMux
    port map (
            O => \N__27518\,
            I => \N__27514\
        );

    \I__4609\ : CEMux
    port map (
            O => \N__27517\,
            I => \N__27511\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__27514\,
            I => \N__27508\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__27511\,
            I => \N__27503\
        );

    \I__4606\ : Span4Mux_v
    port map (
            O => \N__27508\,
            I => \N__27500\
        );

    \I__4605\ : CEMux
    port map (
            O => \N__27507\,
            I => \N__27497\
        );

    \I__4604\ : CEMux
    port map (
            O => \N__27506\,
            I => \N__27494\
        );

    \I__4603\ : Span4Mux_v
    port map (
            O => \N__27503\,
            I => \N__27491\
        );

    \I__4602\ : Span4Mux_h
    port map (
            O => \N__27500\,
            I => \N__27488\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__27497\,
            I => \N__27485\
        );

    \I__4600\ : LocalMux
    port map (
            O => \N__27494\,
            I => \N__27482\
        );

    \I__4599\ : Odrv4
    port map (
            O => \N__27491\,
            I => \current_shift_inst.timer_s1.N_192_i\
        );

    \I__4598\ : Odrv4
    port map (
            O => \N__27488\,
            I => \current_shift_inst.timer_s1.N_192_i\
        );

    \I__4597\ : Odrv4
    port map (
            O => \N__27485\,
            I => \current_shift_inst.timer_s1.N_192_i\
        );

    \I__4596\ : Odrv12
    port map (
            O => \N__27482\,
            I => \current_shift_inst.timer_s1.N_192_i\
        );

    \I__4595\ : InMux
    port map (
            O => \N__27473\,
            I => \N__27467\
        );

    \I__4594\ : InMux
    port map (
            O => \N__27472\,
            I => \N__27462\
        );

    \I__4593\ : InMux
    port map (
            O => \N__27471\,
            I => \N__27462\
        );

    \I__4592\ : InMux
    port map (
            O => \N__27470\,
            I => \N__27459\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__27467\,
            I => \current_shift_inst.timer_phase.runningZ0\
        );

    \I__4590\ : LocalMux
    port map (
            O => \N__27462\,
            I => \current_shift_inst.timer_phase.runningZ0\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__27459\,
            I => \current_shift_inst.timer_phase.runningZ0\
        );

    \I__4588\ : InMux
    port map (
            O => \N__27452\,
            I => \N__27447\
        );

    \I__4587\ : InMux
    port map (
            O => \N__27451\,
            I => \N__27443\
        );

    \I__4586\ : InMux
    port map (
            O => \N__27450\,
            I => \N__27440\
        );

    \I__4585\ : LocalMux
    port map (
            O => \N__27447\,
            I => \N__27437\
        );

    \I__4584\ : InMux
    port map (
            O => \N__27446\,
            I => \N__27434\
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__27443\,
            I => \current_shift_inst.stop_timer_phaseZ0\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__27440\,
            I => \current_shift_inst.stop_timer_phaseZ0\
        );

    \I__4581\ : Odrv4
    port map (
            O => \N__27437\,
            I => \current_shift_inst.stop_timer_phaseZ0\
        );

    \I__4580\ : LocalMux
    port map (
            O => \N__27434\,
            I => \current_shift_inst.stop_timer_phaseZ0\
        );

    \I__4579\ : IoInMux
    port map (
            O => \N__27425\,
            I => \N__27422\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__27422\,
            I => \N__27419\
        );

    \I__4577\ : IoSpan4Mux
    port map (
            O => \N__27419\,
            I => \N__27416\
        );

    \I__4576\ : Span4Mux_s1_v
    port map (
            O => \N__27416\,
            I => \N__27413\
        );

    \I__4575\ : Odrv4
    port map (
            O => \N__27413\,
            I => \current_shift_inst.timer_phase.N_188_i\
        );

    \I__4574\ : InMux
    port map (
            O => \N__27410\,
            I => \N__27407\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__27407\,
            I => \N__27404\
        );

    \I__4572\ : Span12Mux_h
    port map (
            O => \N__27404\,
            I => \N__27401\
        );

    \I__4571\ : Odrv12
    port map (
            O => \N__27401\,
            I => il_max_comp2_c
        );

    \I__4570\ : InMux
    port map (
            O => \N__27398\,
            I => \N__27395\
        );

    \I__4569\ : LocalMux
    port map (
            O => \N__27395\,
            I => \N__27392\
        );

    \I__4568\ : Span4Mux_v
    port map (
            O => \N__27392\,
            I => \N__27389\
        );

    \I__4567\ : Span4Mux_h
    port map (
            O => \N__27389\,
            I => \N__27386\
        );

    \I__4566\ : Odrv4
    port map (
            O => \N__27386\,
            I => il_min_comp2_c
        );

    \I__4565\ : InMux
    port map (
            O => \N__27383\,
            I => \current_shift_inst.timer_s1.counter_cry_20\
        );

    \I__4564\ : InMux
    port map (
            O => \N__27380\,
            I => \current_shift_inst.timer_s1.counter_cry_21\
        );

    \I__4563\ : InMux
    port map (
            O => \N__27377\,
            I => \current_shift_inst.timer_s1.counter_cry_22\
        );

    \I__4562\ : InMux
    port map (
            O => \N__27374\,
            I => \bfn_10_24_0_\
        );

    \I__4561\ : InMux
    port map (
            O => \N__27371\,
            I => \current_shift_inst.timer_s1.counter_cry_24\
        );

    \I__4560\ : InMux
    port map (
            O => \N__27368\,
            I => \current_shift_inst.timer_s1.counter_cry_25\
        );

    \I__4559\ : InMux
    port map (
            O => \N__27365\,
            I => \current_shift_inst.timer_s1.counter_cry_26\
        );

    \I__4558\ : InMux
    port map (
            O => \N__27362\,
            I => \current_shift_inst.timer_s1.counter_cry_27\
        );

    \I__4557\ : InMux
    port map (
            O => \N__27359\,
            I => \N__27325\
        );

    \I__4556\ : InMux
    port map (
            O => \N__27358\,
            I => \N__27325\
        );

    \I__4555\ : InMux
    port map (
            O => \N__27357\,
            I => \N__27316\
        );

    \I__4554\ : InMux
    port map (
            O => \N__27356\,
            I => \N__27316\
        );

    \I__4553\ : InMux
    port map (
            O => \N__27355\,
            I => \N__27316\
        );

    \I__4552\ : InMux
    port map (
            O => \N__27354\,
            I => \N__27316\
        );

    \I__4551\ : InMux
    port map (
            O => \N__27353\,
            I => \N__27307\
        );

    \I__4550\ : InMux
    port map (
            O => \N__27352\,
            I => \N__27307\
        );

    \I__4549\ : InMux
    port map (
            O => \N__27351\,
            I => \N__27307\
        );

    \I__4548\ : InMux
    port map (
            O => \N__27350\,
            I => \N__27307\
        );

    \I__4547\ : InMux
    port map (
            O => \N__27349\,
            I => \N__27298\
        );

    \I__4546\ : InMux
    port map (
            O => \N__27348\,
            I => \N__27298\
        );

    \I__4545\ : InMux
    port map (
            O => \N__27347\,
            I => \N__27298\
        );

    \I__4544\ : InMux
    port map (
            O => \N__27346\,
            I => \N__27298\
        );

    \I__4543\ : InMux
    port map (
            O => \N__27345\,
            I => \N__27289\
        );

    \I__4542\ : InMux
    port map (
            O => \N__27344\,
            I => \N__27289\
        );

    \I__4541\ : InMux
    port map (
            O => \N__27343\,
            I => \N__27289\
        );

    \I__4540\ : InMux
    port map (
            O => \N__27342\,
            I => \N__27289\
        );

    \I__4539\ : InMux
    port map (
            O => \N__27341\,
            I => \N__27280\
        );

    \I__4538\ : InMux
    port map (
            O => \N__27340\,
            I => \N__27280\
        );

    \I__4537\ : InMux
    port map (
            O => \N__27339\,
            I => \N__27280\
        );

    \I__4536\ : InMux
    port map (
            O => \N__27338\,
            I => \N__27280\
        );

    \I__4535\ : InMux
    port map (
            O => \N__27337\,
            I => \N__27271\
        );

    \I__4534\ : InMux
    port map (
            O => \N__27336\,
            I => \N__27271\
        );

    \I__4533\ : InMux
    port map (
            O => \N__27335\,
            I => \N__27271\
        );

    \I__4532\ : InMux
    port map (
            O => \N__27334\,
            I => \N__27271\
        );

    \I__4531\ : InMux
    port map (
            O => \N__27333\,
            I => \N__27262\
        );

    \I__4530\ : InMux
    port map (
            O => \N__27332\,
            I => \N__27262\
        );

    \I__4529\ : InMux
    port map (
            O => \N__27331\,
            I => \N__27262\
        );

    \I__4528\ : InMux
    port map (
            O => \N__27330\,
            I => \N__27262\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__27325\,
            I => \N__27255\
        );

    \I__4526\ : LocalMux
    port map (
            O => \N__27316\,
            I => \N__27255\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__27307\,
            I => \N__27255\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__27298\,
            I => \N__27242\
        );

    \I__4523\ : LocalMux
    port map (
            O => \N__27289\,
            I => \N__27242\
        );

    \I__4522\ : LocalMux
    port map (
            O => \N__27280\,
            I => \N__27242\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__27271\,
            I => \N__27242\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__27262\,
            I => \N__27242\
        );

    \I__4519\ : Sp12to4
    port map (
            O => \N__27255\,
            I => \N__27242\
        );

    \I__4518\ : Odrv12
    port map (
            O => \N__27242\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__4517\ : InMux
    port map (
            O => \N__27239\,
            I => \current_shift_inst.timer_s1.counter_cry_28\
        );

    \I__4516\ : InMux
    port map (
            O => \N__27236\,
            I => \current_shift_inst.timer_s1.counter_cry_10\
        );

    \I__4515\ : InMux
    port map (
            O => \N__27233\,
            I => \current_shift_inst.timer_s1.counter_cry_11\
        );

    \I__4514\ : InMux
    port map (
            O => \N__27230\,
            I => \current_shift_inst.timer_s1.counter_cry_12\
        );

    \I__4513\ : InMux
    port map (
            O => \N__27227\,
            I => \current_shift_inst.timer_s1.counter_cry_13\
        );

    \I__4512\ : InMux
    port map (
            O => \N__27224\,
            I => \current_shift_inst.timer_s1.counter_cry_14\
        );

    \I__4511\ : InMux
    port map (
            O => \N__27221\,
            I => \bfn_10_23_0_\
        );

    \I__4510\ : InMux
    port map (
            O => \N__27218\,
            I => \current_shift_inst.timer_s1.counter_cry_16\
        );

    \I__4509\ : InMux
    port map (
            O => \N__27215\,
            I => \current_shift_inst.timer_s1.counter_cry_17\
        );

    \I__4508\ : InMux
    port map (
            O => \N__27212\,
            I => \current_shift_inst.timer_s1.counter_cry_18\
        );

    \I__4507\ : InMux
    port map (
            O => \N__27209\,
            I => \current_shift_inst.timer_s1.counter_cry_19\
        );

    \I__4506\ : InMux
    port map (
            O => \N__27206\,
            I => \current_shift_inst.timer_s1.counter_cry_1\
        );

    \I__4505\ : InMux
    port map (
            O => \N__27203\,
            I => \current_shift_inst.timer_s1.counter_cry_2\
        );

    \I__4504\ : InMux
    port map (
            O => \N__27200\,
            I => \current_shift_inst.timer_s1.counter_cry_3\
        );

    \I__4503\ : InMux
    port map (
            O => \N__27197\,
            I => \current_shift_inst.timer_s1.counter_cry_4\
        );

    \I__4502\ : InMux
    port map (
            O => \N__27194\,
            I => \current_shift_inst.timer_s1.counter_cry_5\
        );

    \I__4501\ : InMux
    port map (
            O => \N__27191\,
            I => \current_shift_inst.timer_s1.counter_cry_6\
        );

    \I__4500\ : InMux
    port map (
            O => \N__27188\,
            I => \bfn_10_22_0_\
        );

    \I__4499\ : InMux
    port map (
            O => \N__27185\,
            I => \current_shift_inst.timer_s1.counter_cry_8\
        );

    \I__4498\ : InMux
    port map (
            O => \N__27182\,
            I => \current_shift_inst.timer_s1.counter_cry_9\
        );

    \I__4497\ : InMux
    port map (
            O => \N__27179\,
            I => \current_shift_inst.un4_control_input_cry_26\
        );

    \I__4496\ : InMux
    port map (
            O => \N__27176\,
            I => \current_shift_inst.un4_control_input_cry_27\
        );

    \I__4495\ : InMux
    port map (
            O => \N__27173\,
            I => \current_shift_inst.un4_control_input_cry_28\
        );

    \I__4494\ : InMux
    port map (
            O => \N__27170\,
            I => \N__27164\
        );

    \I__4493\ : InMux
    port map (
            O => \N__27169\,
            I => \N__27164\
        );

    \I__4492\ : LocalMux
    port map (
            O => \N__27164\,
            I => \N__27161\
        );

    \I__4491\ : Span4Mux_h
    port map (
            O => \N__27161\,
            I => \N__27157\
        );

    \I__4490\ : InMux
    port map (
            O => \N__27160\,
            I => \N__27154\
        );

    \I__4489\ : Odrv4
    port map (
            O => \N__27157\,
            I => \current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__27154\,
            I => \current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0\
        );

    \I__4487\ : InMux
    port map (
            O => \N__27149\,
            I => \current_shift_inst.un4_control_input_cry_29\
        );

    \I__4486\ : CascadeMux
    port map (
            O => \N__27146\,
            I => \N__27143\
        );

    \I__4485\ : InMux
    port map (
            O => \N__27143\,
            I => \N__27139\
        );

    \I__4484\ : InMux
    port map (
            O => \N__27142\,
            I => \N__27136\
        );

    \I__4483\ : LocalMux
    port map (
            O => \N__27139\,
            I => \N__27126\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__27136\,
            I => \N__27126\
        );

    \I__4481\ : InMux
    port map (
            O => \N__27135\,
            I => \N__27123\
        );

    \I__4480\ : InMux
    port map (
            O => \N__27134\,
            I => \N__27120\
        );

    \I__4479\ : InMux
    port map (
            O => \N__27133\,
            I => \N__27116\
        );

    \I__4478\ : CascadeMux
    port map (
            O => \N__27132\,
            I => \N__27113\
        );

    \I__4477\ : CascadeMux
    port map (
            O => \N__27131\,
            I => \N__27109\
        );

    \I__4476\ : Span4Mux_v
    port map (
            O => \N__27126\,
            I => \N__27106\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__27123\,
            I => \N__27103\
        );

    \I__4474\ : LocalMux
    port map (
            O => \N__27120\,
            I => \N__27100\
        );

    \I__4473\ : InMux
    port map (
            O => \N__27119\,
            I => \N__27097\
        );

    \I__4472\ : LocalMux
    port map (
            O => \N__27116\,
            I => \N__27094\
        );

    \I__4471\ : InMux
    port map (
            O => \N__27113\,
            I => \N__27087\
        );

    \I__4470\ : InMux
    port map (
            O => \N__27112\,
            I => \N__27087\
        );

    \I__4469\ : InMux
    port map (
            O => \N__27109\,
            I => \N__27087\
        );

    \I__4468\ : Span4Mux_v
    port map (
            O => \N__27106\,
            I => \N__27082\
        );

    \I__4467\ : Span4Mux_v
    port map (
            O => \N__27103\,
            I => \N__27082\
        );

    \I__4466\ : Span4Mux_h
    port map (
            O => \N__27100\,
            I => \N__27079\
        );

    \I__4465\ : LocalMux
    port map (
            O => \N__27097\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__4464\ : Odrv12
    port map (
            O => \N__27094\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__4463\ : LocalMux
    port map (
            O => \N__27087\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__4462\ : Odrv4
    port map (
            O => \N__27082\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__4461\ : Odrv4
    port map (
            O => \N__27079\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__4460\ : InMux
    port map (
            O => \N__27068\,
            I => \current_shift_inst.un4_control_input_cry_30\
        );

    \I__4459\ : InMux
    port map (
            O => \N__27065\,
            I => \N__27059\
        );

    \I__4458\ : InMux
    port map (
            O => \N__27064\,
            I => \N__27059\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__27059\,
            I => \N__27056\
        );

    \I__4456\ : Span4Mux_h
    port map (
            O => \N__27056\,
            I => \N__27052\
        );

    \I__4455\ : InMux
    port map (
            O => \N__27055\,
            I => \N__27049\
        );

    \I__4454\ : Odrv4
    port map (
            O => \N__27052\,
            I => \current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0\
        );

    \I__4453\ : LocalMux
    port map (
            O => \N__27049\,
            I => \current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0\
        );

    \I__4452\ : InMux
    port map (
            O => \N__27044\,
            I => \N__27039\
        );

    \I__4451\ : InMux
    port map (
            O => \N__27043\,
            I => \N__27033\
        );

    \I__4450\ : InMux
    port map (
            O => \N__27042\,
            I => \N__27033\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__27039\,
            I => \N__27030\
        );

    \I__4448\ : InMux
    port map (
            O => \N__27038\,
            I => \N__27027\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__27033\,
            I => \N__27024\
        );

    \I__4446\ : Span4Mux_h
    port map (
            O => \N__27030\,
            I => \N__27021\
        );

    \I__4445\ : LocalMux
    port map (
            O => \N__27027\,
            I => \N__27018\
        );

    \I__4444\ : Odrv12
    port map (
            O => \N__27024\,
            I => \current_shift_inst.elapsed_time_ns_phase_28\
        );

    \I__4443\ : Odrv4
    port map (
            O => \N__27021\,
            I => \current_shift_inst.elapsed_time_ns_phase_28\
        );

    \I__4442\ : Odrv4
    port map (
            O => \N__27018\,
            I => \current_shift_inst.elapsed_time_ns_phase_28\
        );

    \I__4441\ : CascadeMux
    port map (
            O => \N__27011\,
            I => \N__27008\
        );

    \I__4440\ : InMux
    port map (
            O => \N__27008\,
            I => \N__27002\
        );

    \I__4439\ : InMux
    port map (
            O => \N__27007\,
            I => \N__27002\
        );

    \I__4438\ : LocalMux
    port map (
            O => \N__27002\,
            I => \N__26997\
        );

    \I__4437\ : CascadeMux
    port map (
            O => \N__27001\,
            I => \N__26994\
        );

    \I__4436\ : InMux
    port map (
            O => \N__27000\,
            I => \N__26991\
        );

    \I__4435\ : Span4Mux_h
    port map (
            O => \N__26997\,
            I => \N__26988\
        );

    \I__4434\ : InMux
    port map (
            O => \N__26994\,
            I => \N__26985\
        );

    \I__4433\ : LocalMux
    port map (
            O => \N__26991\,
            I => \current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0\
        );

    \I__4432\ : Odrv4
    port map (
            O => \N__26988\,
            I => \current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0\
        );

    \I__4431\ : LocalMux
    port map (
            O => \N__26985\,
            I => \current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0\
        );

    \I__4430\ : InMux
    port map (
            O => \N__26978\,
            I => \N__26975\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__26975\,
            I => \N__26972\
        );

    \I__4428\ : Span4Mux_v
    port map (
            O => \N__26972\,
            I => \N__26969\
        );

    \I__4427\ : Odrv4
    port map (
            O => \N__26969\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINKG81_27\
        );

    \I__4426\ : InMux
    port map (
            O => \N__26966\,
            I => \bfn_10_21_0_\
        );

    \I__4425\ : InMux
    port map (
            O => \N__26963\,
            I => \current_shift_inst.timer_s1.counter_cry_0\
        );

    \I__4424\ : CascadeMux
    port map (
            O => \N__26960\,
            I => \N__26956\
        );

    \I__4423\ : CascadeMux
    port map (
            O => \N__26959\,
            I => \N__26953\
        );

    \I__4422\ : InMux
    port map (
            O => \N__26956\,
            I => \N__26948\
        );

    \I__4421\ : InMux
    port map (
            O => \N__26953\,
            I => \N__26943\
        );

    \I__4420\ : InMux
    port map (
            O => \N__26952\,
            I => \N__26943\
        );

    \I__4419\ : CascadeMux
    port map (
            O => \N__26951\,
            I => \N__26940\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__26948\,
            I => \N__26937\
        );

    \I__4417\ : LocalMux
    port map (
            O => \N__26943\,
            I => \N__26934\
        );

    \I__4416\ : InMux
    port map (
            O => \N__26940\,
            I => \N__26931\
        );

    \I__4415\ : Odrv4
    port map (
            O => \N__26937\,
            I => \current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0\
        );

    \I__4414\ : Odrv4
    port map (
            O => \N__26934\,
            I => \current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0\
        );

    \I__4413\ : LocalMux
    port map (
            O => \N__26931\,
            I => \current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0\
        );

    \I__4412\ : InMux
    port map (
            O => \N__26924\,
            I => \current_shift_inst.un4_control_input_cry_17\
        );

    \I__4411\ : CascadeMux
    port map (
            O => \N__26921\,
            I => \N__26918\
        );

    \I__4410\ : InMux
    port map (
            O => \N__26918\,
            I => \N__26915\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__26915\,
            I => \N__26909\
        );

    \I__4408\ : InMux
    port map (
            O => \N__26914\,
            I => \N__26904\
        );

    \I__4407\ : InMux
    port map (
            O => \N__26913\,
            I => \N__26904\
        );

    \I__4406\ : CascadeMux
    port map (
            O => \N__26912\,
            I => \N__26901\
        );

    \I__4405\ : Span4Mux_v
    port map (
            O => \N__26909\,
            I => \N__26896\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__26904\,
            I => \N__26896\
        );

    \I__4403\ : InMux
    port map (
            O => \N__26901\,
            I => \N__26893\
        );

    \I__4402\ : Odrv4
    port map (
            O => \N__26896\,
            I => \current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__26893\,
            I => \current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0\
        );

    \I__4400\ : InMux
    port map (
            O => \N__26888\,
            I => \current_shift_inst.un4_control_input_cry_18\
        );

    \I__4399\ : CascadeMux
    port map (
            O => \N__26885\,
            I => \N__26882\
        );

    \I__4398\ : InMux
    port map (
            O => \N__26882\,
            I => \N__26879\
        );

    \I__4397\ : LocalMux
    port map (
            O => \N__26879\,
            I => \N__26874\
        );

    \I__4396\ : InMux
    port map (
            O => \N__26878\,
            I => \N__26869\
        );

    \I__4395\ : InMux
    port map (
            O => \N__26877\,
            I => \N__26869\
        );

    \I__4394\ : Span4Mux_v
    port map (
            O => \N__26874\,
            I => \N__26863\
        );

    \I__4393\ : LocalMux
    port map (
            O => \N__26869\,
            I => \N__26863\
        );

    \I__4392\ : CascadeMux
    port map (
            O => \N__26868\,
            I => \N__26860\
        );

    \I__4391\ : Span4Mux_h
    port map (
            O => \N__26863\,
            I => \N__26857\
        );

    \I__4390\ : InMux
    port map (
            O => \N__26860\,
            I => \N__26854\
        );

    \I__4389\ : Odrv4
    port map (
            O => \N__26857\,
            I => \current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__26854\,
            I => \current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0\
        );

    \I__4387\ : InMux
    port map (
            O => \N__26849\,
            I => \current_shift_inst.un4_control_input_cry_19\
        );

    \I__4386\ : CascadeMux
    port map (
            O => \N__26846\,
            I => \N__26843\
        );

    \I__4385\ : InMux
    port map (
            O => \N__26843\,
            I => \N__26837\
        );

    \I__4384\ : InMux
    port map (
            O => \N__26842\,
            I => \N__26832\
        );

    \I__4383\ : InMux
    port map (
            O => \N__26841\,
            I => \N__26832\
        );

    \I__4382\ : CascadeMux
    port map (
            O => \N__26840\,
            I => \N__26829\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__26837\,
            I => \N__26824\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__26832\,
            I => \N__26824\
        );

    \I__4379\ : InMux
    port map (
            O => \N__26829\,
            I => \N__26821\
        );

    \I__4378\ : Odrv4
    port map (
            O => \N__26824\,
            I => \current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0\
        );

    \I__4377\ : LocalMux
    port map (
            O => \N__26821\,
            I => \current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0\
        );

    \I__4376\ : InMux
    port map (
            O => \N__26816\,
            I => \current_shift_inst.un4_control_input_cry_20\
        );

    \I__4375\ : InMux
    port map (
            O => \N__26813\,
            I => \N__26807\
        );

    \I__4374\ : InMux
    port map (
            O => \N__26812\,
            I => \N__26807\
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__26807\,
            I => \N__26803\
        );

    \I__4372\ : InMux
    port map (
            O => \N__26806\,
            I => \N__26800\
        );

    \I__4371\ : Span4Mux_h
    port map (
            O => \N__26803\,
            I => \N__26794\
        );

    \I__4370\ : LocalMux
    port map (
            O => \N__26800\,
            I => \N__26794\
        );

    \I__4369\ : InMux
    port map (
            O => \N__26799\,
            I => \N__26791\
        );

    \I__4368\ : Odrv4
    port map (
            O => \N__26794\,
            I => \current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__26791\,
            I => \current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0\
        );

    \I__4366\ : InMux
    port map (
            O => \N__26786\,
            I => \current_shift_inst.un4_control_input_cry_21\
        );

    \I__4365\ : InMux
    port map (
            O => \N__26783\,
            I => \current_shift_inst.un4_control_input_cry_22\
        );

    \I__4364\ : InMux
    port map (
            O => \N__26780\,
            I => \current_shift_inst.un4_control_input_cry_23\
        );

    \I__4363\ : InMux
    port map (
            O => \N__26777\,
            I => \bfn_10_20_0_\
        );

    \I__4362\ : InMux
    port map (
            O => \N__26774\,
            I => \current_shift_inst.un4_control_input_cry_25\
        );

    \I__4361\ : InMux
    port map (
            O => \N__26771\,
            I => \N__26766\
        );

    \I__4360\ : InMux
    port map (
            O => \N__26770\,
            I => \N__26760\
        );

    \I__4359\ : InMux
    port map (
            O => \N__26769\,
            I => \N__26760\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__26766\,
            I => \N__26757\
        );

    \I__4357\ : CascadeMux
    port map (
            O => \N__26765\,
            I => \N__26754\
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__26760\,
            I => \N__26751\
        );

    \I__4355\ : Span4Mux_v
    port map (
            O => \N__26757\,
            I => \N__26748\
        );

    \I__4354\ : InMux
    port map (
            O => \N__26754\,
            I => \N__26745\
        );

    \I__4353\ : Odrv4
    port map (
            O => \N__26751\,
            I => \current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0\
        );

    \I__4352\ : Odrv4
    port map (
            O => \N__26748\,
            I => \current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0\
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__26745\,
            I => \current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0\
        );

    \I__4350\ : InMux
    port map (
            O => \N__26738\,
            I => \bfn_10_18_0_\
        );

    \I__4349\ : CascadeMux
    port map (
            O => \N__26735\,
            I => \N__26731\
        );

    \I__4348\ : InMux
    port map (
            O => \N__26734\,
            I => \N__26727\
        );

    \I__4347\ : InMux
    port map (
            O => \N__26731\,
            I => \N__26724\
        );

    \I__4346\ : InMux
    port map (
            O => \N__26730\,
            I => \N__26721\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__26727\,
            I => \N__26715\
        );

    \I__4344\ : LocalMux
    port map (
            O => \N__26724\,
            I => \N__26715\
        );

    \I__4343\ : LocalMux
    port map (
            O => \N__26721\,
            I => \N__26712\
        );

    \I__4342\ : CascadeMux
    port map (
            O => \N__26720\,
            I => \N__26709\
        );

    \I__4341\ : Span4Mux_v
    port map (
            O => \N__26715\,
            I => \N__26704\
        );

    \I__4340\ : Span4Mux_v
    port map (
            O => \N__26712\,
            I => \N__26704\
        );

    \I__4339\ : InMux
    port map (
            O => \N__26709\,
            I => \N__26701\
        );

    \I__4338\ : Odrv4
    port map (
            O => \N__26704\,
            I => \current_shift_inst.un4_control_input_cry_9_c_RNIALDJZ0\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__26701\,
            I => \current_shift_inst.un4_control_input_cry_9_c_RNIALDJZ0\
        );

    \I__4336\ : InMux
    port map (
            O => \N__26696\,
            I => \current_shift_inst.un4_control_input_cry_9\
        );

    \I__4335\ : CascadeMux
    port map (
            O => \N__26693\,
            I => \N__26690\
        );

    \I__4334\ : InMux
    port map (
            O => \N__26690\,
            I => \N__26685\
        );

    \I__4333\ : InMux
    port map (
            O => \N__26689\,
            I => \N__26682\
        );

    \I__4332\ : InMux
    port map (
            O => \N__26688\,
            I => \N__26678\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__26685\,
            I => \N__26673\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__26682\,
            I => \N__26673\
        );

    \I__4329\ : CascadeMux
    port map (
            O => \N__26681\,
            I => \N__26670\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__26678\,
            I => \N__26665\
        );

    \I__4327\ : Span4Mux_h
    port map (
            O => \N__26673\,
            I => \N__26665\
        );

    \I__4326\ : InMux
    port map (
            O => \N__26670\,
            I => \N__26662\
        );

    \I__4325\ : Odrv4
    port map (
            O => \N__26665\,
            I => \current_shift_inst.un4_control_input_cry_10_c_RNIJLTGZ0\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__26662\,
            I => \current_shift_inst.un4_control_input_cry_10_c_RNIJLTGZ0\
        );

    \I__4323\ : InMux
    port map (
            O => \N__26657\,
            I => \current_shift_inst.un4_control_input_cry_10\
        );

    \I__4322\ : InMux
    port map (
            O => \N__26654\,
            I => \current_shift_inst.un4_control_input_cry_11\
        );

    \I__4321\ : InMux
    port map (
            O => \N__26651\,
            I => \current_shift_inst.un4_control_input_cry_12\
        );

    \I__4320\ : CascadeMux
    port map (
            O => \N__26648\,
            I => \N__26644\
        );

    \I__4319\ : InMux
    port map (
            O => \N__26647\,
            I => \N__26640\
        );

    \I__4318\ : InMux
    port map (
            O => \N__26644\,
            I => \N__26635\
        );

    \I__4317\ : InMux
    port map (
            O => \N__26643\,
            I => \N__26635\
        );

    \I__4316\ : LocalMux
    port map (
            O => \N__26640\,
            I => \N__26631\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__26635\,
            I => \N__26628\
        );

    \I__4314\ : CascadeMux
    port map (
            O => \N__26634\,
            I => \N__26625\
        );

    \I__4313\ : Span4Mux_v
    port map (
            O => \N__26631\,
            I => \N__26622\
        );

    \I__4312\ : Span4Mux_h
    port map (
            O => \N__26628\,
            I => \N__26619\
        );

    \I__4311\ : InMux
    port map (
            O => \N__26625\,
            I => \N__26616\
        );

    \I__4310\ : Odrv4
    port map (
            O => \N__26622\,
            I => \current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0\
        );

    \I__4309\ : Odrv4
    port map (
            O => \N__26619\,
            I => \current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__26616\,
            I => \current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0\
        );

    \I__4307\ : InMux
    port map (
            O => \N__26609\,
            I => \current_shift_inst.un4_control_input_cry_13\
        );

    \I__4306\ : CascadeMux
    port map (
            O => \N__26606\,
            I => \N__26603\
        );

    \I__4305\ : InMux
    port map (
            O => \N__26603\,
            I => \N__26600\
        );

    \I__4304\ : LocalMux
    port map (
            O => \N__26600\,
            I => \N__26594\
        );

    \I__4303\ : InMux
    port map (
            O => \N__26599\,
            I => \N__26591\
        );

    \I__4302\ : InMux
    port map (
            O => \N__26598\,
            I => \N__26588\
        );

    \I__4301\ : CascadeMux
    port map (
            O => \N__26597\,
            I => \N__26585\
        );

    \I__4300\ : Sp12to4
    port map (
            O => \N__26594\,
            I => \N__26578\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__26591\,
            I => \N__26578\
        );

    \I__4298\ : LocalMux
    port map (
            O => \N__26588\,
            I => \N__26578\
        );

    \I__4297\ : InMux
    port map (
            O => \N__26585\,
            I => \N__26575\
        );

    \I__4296\ : Odrv12
    port map (
            O => \N__26578\,
            I => \current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0\
        );

    \I__4295\ : LocalMux
    port map (
            O => \N__26575\,
            I => \current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0\
        );

    \I__4294\ : InMux
    port map (
            O => \N__26570\,
            I => \current_shift_inst.un4_control_input_cry_14\
        );

    \I__4293\ : InMux
    port map (
            O => \N__26567\,
            I => \N__26562\
        );

    \I__4292\ : InMux
    port map (
            O => \N__26566\,
            I => \N__26557\
        );

    \I__4291\ : InMux
    port map (
            O => \N__26565\,
            I => \N__26557\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__26562\,
            I => \N__26551\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__26557\,
            I => \N__26551\
        );

    \I__4288\ : InMux
    port map (
            O => \N__26556\,
            I => \N__26548\
        );

    \I__4287\ : Odrv12
    port map (
            O => \N__26551\,
            I => \current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__26548\,
            I => \current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0\
        );

    \I__4285\ : InMux
    port map (
            O => \N__26543\,
            I => \current_shift_inst.un4_control_input_cry_15\
        );

    \I__4284\ : InMux
    port map (
            O => \N__26540\,
            I => \N__26535\
        );

    \I__4283\ : InMux
    port map (
            O => \N__26539\,
            I => \N__26530\
        );

    \I__4282\ : InMux
    port map (
            O => \N__26538\,
            I => \N__26530\
        );

    \I__4281\ : LocalMux
    port map (
            O => \N__26535\,
            I => \N__26525\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__26530\,
            I => \N__26525\
        );

    \I__4279\ : Span4Mux_v
    port map (
            O => \N__26525\,
            I => \N__26521\
        );

    \I__4278\ : InMux
    port map (
            O => \N__26524\,
            I => \N__26518\
        );

    \I__4277\ : Odrv4
    port map (
            O => \N__26521\,
            I => \current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0\
        );

    \I__4276\ : LocalMux
    port map (
            O => \N__26518\,
            I => \current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0\
        );

    \I__4275\ : InMux
    port map (
            O => \N__26513\,
            I => \bfn_10_19_0_\
        );

    \I__4274\ : CascadeMux
    port map (
            O => \N__26510\,
            I => \N__26507\
        );

    \I__4273\ : InMux
    port map (
            O => \N__26507\,
            I => \N__26504\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__26504\,
            I => \N__26501\
        );

    \I__4271\ : Span4Mux_h
    port map (
            O => \N__26501\,
            I => \N__26497\
        );

    \I__4270\ : InMux
    port map (
            O => \N__26500\,
            I => \N__26494\
        );

    \I__4269\ : Odrv4
    port map (
            O => \N__26497\,
            I => \current_shift_inst.un38_control_input_0\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__26494\,
            I => \current_shift_inst.un38_control_input_0\
        );

    \I__4267\ : InMux
    port map (
            O => \N__26489\,
            I => \N__26485\
        );

    \I__4266\ : InMux
    port map (
            O => \N__26488\,
            I => \N__26482\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__26485\,
            I => \N__26479\
        );

    \I__4264\ : LocalMux
    port map (
            O => \N__26482\,
            I => \N__26476\
        );

    \I__4263\ : Span4Mux_v
    port map (
            O => \N__26479\,
            I => \N__26472\
        );

    \I__4262\ : Span4Mux_h
    port map (
            O => \N__26476\,
            I => \N__26469\
        );

    \I__4261\ : InMux
    port map (
            O => \N__26475\,
            I => \N__26466\
        );

    \I__4260\ : Odrv4
    port map (
            O => \N__26472\,
            I => \current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0\
        );

    \I__4259\ : Odrv4
    port map (
            O => \N__26469\,
            I => \current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__26466\,
            I => \current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0\
        );

    \I__4257\ : InMux
    port map (
            O => \N__26459\,
            I => \current_shift_inst.un4_control_input_cry_1\
        );

    \I__4256\ : CascadeMux
    port map (
            O => \N__26456\,
            I => \N__26452\
        );

    \I__4255\ : InMux
    port map (
            O => \N__26455\,
            I => \N__26449\
        );

    \I__4254\ : InMux
    port map (
            O => \N__26452\,
            I => \N__26445\
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__26449\,
            I => \N__26442\
        );

    \I__4252\ : CascadeMux
    port map (
            O => \N__26448\,
            I => \N__26439\
        );

    \I__4251\ : LocalMux
    port map (
            O => \N__26445\,
            I => \N__26436\
        );

    \I__4250\ : Span4Mux_h
    port map (
            O => \N__26442\,
            I => \N__26433\
        );

    \I__4249\ : InMux
    port map (
            O => \N__26439\,
            I => \N__26430\
        );

    \I__4248\ : Odrv12
    port map (
            O => \N__26436\,
            I => \current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0\
        );

    \I__4247\ : Odrv4
    port map (
            O => \N__26433\,
            I => \current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0\
        );

    \I__4246\ : LocalMux
    port map (
            O => \N__26430\,
            I => \current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0\
        );

    \I__4245\ : InMux
    port map (
            O => \N__26423\,
            I => \current_shift_inst.un4_control_input_cry_2\
        );

    \I__4244\ : InMux
    port map (
            O => \N__26420\,
            I => \N__26417\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__26417\,
            I => \N__26414\
        );

    \I__4242\ : Span4Mux_h
    port map (
            O => \N__26414\,
            I => \N__26410\
        );

    \I__4241\ : InMux
    port map (
            O => \N__26413\,
            I => \N__26407\
        );

    \I__4240\ : Odrv4
    port map (
            O => \N__26410\,
            I => \current_shift_inst.un4_control_input_cry_3_c_RNINL4GZ0\
        );

    \I__4239\ : LocalMux
    port map (
            O => \N__26407\,
            I => \current_shift_inst.un4_control_input_cry_3_c_RNINL4GZ0\
        );

    \I__4238\ : InMux
    port map (
            O => \N__26402\,
            I => \current_shift_inst.un4_control_input_cry_3\
        );

    \I__4237\ : InMux
    port map (
            O => \N__26399\,
            I => \N__26394\
        );

    \I__4236\ : InMux
    port map (
            O => \N__26398\,
            I => \N__26389\
        );

    \I__4235\ : InMux
    port map (
            O => \N__26397\,
            I => \N__26389\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__26394\,
            I => \N__26383\
        );

    \I__4233\ : LocalMux
    port map (
            O => \N__26389\,
            I => \N__26383\
        );

    \I__4232\ : InMux
    port map (
            O => \N__26388\,
            I => \N__26380\
        );

    \I__4231\ : Odrv12
    port map (
            O => \N__26383\,
            I => \current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0\
        );

    \I__4230\ : LocalMux
    port map (
            O => \N__26380\,
            I => \current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0\
        );

    \I__4229\ : InMux
    port map (
            O => \N__26375\,
            I => \current_shift_inst.un4_control_input_cry_4\
        );

    \I__4228\ : CascadeMux
    port map (
            O => \N__26372\,
            I => \N__26369\
        );

    \I__4227\ : InMux
    port map (
            O => \N__26369\,
            I => \N__26359\
        );

    \I__4226\ : InMux
    port map (
            O => \N__26368\,
            I => \N__26359\
        );

    \I__4225\ : InMux
    port map (
            O => \N__26367\,
            I => \N__26359\
        );

    \I__4224\ : CascadeMux
    port map (
            O => \N__26366\,
            I => \N__26356\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__26359\,
            I => \N__26353\
        );

    \I__4222\ : InMux
    port map (
            O => \N__26356\,
            I => \N__26350\
        );

    \I__4221\ : Odrv12
    port map (
            O => \N__26353\,
            I => \current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0\
        );

    \I__4220\ : LocalMux
    port map (
            O => \N__26350\,
            I => \current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0\
        );

    \I__4219\ : InMux
    port map (
            O => \N__26345\,
            I => \current_shift_inst.un4_control_input_cry_5\
        );

    \I__4218\ : CascadeMux
    port map (
            O => \N__26342\,
            I => \N__26339\
        );

    \I__4217\ : InMux
    port map (
            O => \N__26339\,
            I => \N__26331\
        );

    \I__4216\ : InMux
    port map (
            O => \N__26338\,
            I => \N__26331\
        );

    \I__4215\ : InMux
    port map (
            O => \N__26337\,
            I => \N__26328\
        );

    \I__4214\ : CascadeMux
    port map (
            O => \N__26336\,
            I => \N__26325\
        );

    \I__4213\ : LocalMux
    port map (
            O => \N__26331\,
            I => \N__26320\
        );

    \I__4212\ : LocalMux
    port map (
            O => \N__26328\,
            I => \N__26320\
        );

    \I__4211\ : InMux
    port map (
            O => \N__26325\,
            I => \N__26317\
        );

    \I__4210\ : Odrv12
    port map (
            O => \N__26320\,
            I => \current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__26317\,
            I => \current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0\
        );

    \I__4208\ : InMux
    port map (
            O => \N__26312\,
            I => \current_shift_inst.un4_control_input_cry_6\
        );

    \I__4207\ : CascadeMux
    port map (
            O => \N__26309\,
            I => \N__26306\
        );

    \I__4206\ : InMux
    port map (
            O => \N__26306\,
            I => \N__26300\
        );

    \I__4205\ : InMux
    port map (
            O => \N__26305\,
            I => \N__26295\
        );

    \I__4204\ : InMux
    port map (
            O => \N__26304\,
            I => \N__26295\
        );

    \I__4203\ : CascadeMux
    port map (
            O => \N__26303\,
            I => \N__26292\
        );

    \I__4202\ : LocalMux
    port map (
            O => \N__26300\,
            I => \N__26287\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__26295\,
            I => \N__26287\
        );

    \I__4200\ : InMux
    port map (
            O => \N__26292\,
            I => \N__26284\
        );

    \I__4199\ : Odrv12
    port map (
            O => \N__26287\,
            I => \current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__26284\,
            I => \current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0\
        );

    \I__4197\ : InMux
    port map (
            O => \N__26279\,
            I => \current_shift_inst.un4_control_input_cry_7\
        );

    \I__4196\ : CascadeMux
    port map (
            O => \N__26276\,
            I => \N__26273\
        );

    \I__4195\ : InMux
    port map (
            O => \N__26273\,
            I => \N__26270\
        );

    \I__4194\ : LocalMux
    port map (
            O => \N__26270\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIOV0K_21\
        );

    \I__4193\ : CascadeMux
    port map (
            O => \N__26267\,
            I => \N__26264\
        );

    \I__4192\ : InMux
    port map (
            O => \N__26264\,
            I => \N__26261\
        );

    \I__4191\ : LocalMux
    port map (
            O => \N__26261\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIAL3J_18\
        );

    \I__4190\ : CascadeMux
    port map (
            O => \N__26258\,
            I => \N__26255\
        );

    \I__4189\ : InMux
    port map (
            O => \N__26255\,
            I => \N__26252\
        );

    \I__4188\ : LocalMux
    port map (
            O => \N__26252\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI7H2J_17\
        );

    \I__4187\ : CascadeMux
    port map (
            O => \N__26249\,
            I => \N__26246\
        );

    \I__4186\ : InMux
    port map (
            O => \N__26246\,
            I => \N__26243\
        );

    \I__4185\ : LocalMux
    port map (
            O => \N__26243\,
            I => \current_shift_inst.elapsed_time_ns_1_RNILRVJ_20\
        );

    \I__4184\ : InMux
    port map (
            O => \N__26240\,
            I => \N__26236\
        );

    \I__4183\ : CascadeMux
    port map (
            O => \N__26239\,
            I => \N__26233\
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__26236\,
            I => \N__26229\
        );

    \I__4181\ : InMux
    port map (
            O => \N__26233\,
            I => \N__26224\
        );

    \I__4180\ : InMux
    port map (
            O => \N__26232\,
            I => \N__26224\
        );

    \I__4179\ : Span4Mux_v
    port map (
            O => \N__26229\,
            I => \N__26219\
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__26224\,
            I => \N__26219\
        );

    \I__4177\ : Span4Mux_h
    port map (
            O => \N__26219\,
            I => \N__26215\
        );

    \I__4176\ : InMux
    port map (
            O => \N__26218\,
            I => \N__26212\
        );

    \I__4175\ : Span4Mux_v
    port map (
            O => \N__26215\,
            I => \N__26209\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__26212\,
            I => \N__26206\
        );

    \I__4173\ : Odrv4
    port map (
            O => \N__26209\,
            I => \current_shift_inst.elapsed_time_ns_phase_19\
        );

    \I__4172\ : Odrv4
    port map (
            O => \N__26206\,
            I => \current_shift_inst.elapsed_time_ns_phase_19\
        );

    \I__4171\ : InMux
    port map (
            O => \N__26201\,
            I => \N__26198\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__26198\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPC571_19\
        );

    \I__4169\ : InMux
    port map (
            O => \N__26195\,
            I => \N__26189\
        );

    \I__4168\ : InMux
    port map (
            O => \N__26194\,
            I => \N__26189\
        );

    \I__4167\ : LocalMux
    port map (
            O => \N__26189\,
            I => \N__26184\
        );

    \I__4166\ : InMux
    port map (
            O => \N__26188\,
            I => \N__26181\
        );

    \I__4165\ : CascadeMux
    port map (
            O => \N__26187\,
            I => \N__26178\
        );

    \I__4164\ : Span4Mux_h
    port map (
            O => \N__26184\,
            I => \N__26175\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__26181\,
            I => \N__26172\
        );

    \I__4162\ : InMux
    port map (
            O => \N__26178\,
            I => \N__26169\
        );

    \I__4161\ : Span4Mux_v
    port map (
            O => \N__26175\,
            I => \N__26166\
        );

    \I__4160\ : Span4Mux_h
    port map (
            O => \N__26172\,
            I => \N__26161\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__26169\,
            I => \N__26161\
        );

    \I__4158\ : Odrv4
    port map (
            O => \N__26166\,
            I => \current_shift_inst.elapsed_time_ns_phase_16\
        );

    \I__4157\ : Odrv4
    port map (
            O => \N__26161\,
            I => \current_shift_inst.elapsed_time_ns_phase_16\
        );

    \I__4156\ : InMux
    port map (
            O => \N__26156\,
            I => \N__26153\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__26153\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIBU361_16\
        );

    \I__4154\ : CascadeMux
    port map (
            O => \N__26150\,
            I => \N__26147\
        );

    \I__4153\ : InMux
    port map (
            O => \N__26147\,
            I => \N__26141\
        );

    \I__4152\ : InMux
    port map (
            O => \N__26146\,
            I => \N__26141\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__26141\,
            I => \N__26136\
        );

    \I__4150\ : InMux
    port map (
            O => \N__26140\,
            I => \N__26133\
        );

    \I__4149\ : CascadeMux
    port map (
            O => \N__26139\,
            I => \N__26130\
        );

    \I__4148\ : Span4Mux_h
    port map (
            O => \N__26136\,
            I => \N__26127\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__26133\,
            I => \N__26124\
        );

    \I__4146\ : InMux
    port map (
            O => \N__26130\,
            I => \N__26121\
        );

    \I__4145\ : Span4Mux_v
    port map (
            O => \N__26127\,
            I => \N__26118\
        );

    \I__4144\ : Span4Mux_h
    port map (
            O => \N__26124\,
            I => \N__26113\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__26121\,
            I => \N__26113\
        );

    \I__4142\ : Odrv4
    port map (
            O => \N__26118\,
            I => \current_shift_inst.elapsed_time_ns_phase_15\
        );

    \I__4141\ : Odrv4
    port map (
            O => \N__26113\,
            I => \current_shift_inst.elapsed_time_ns_phase_15\
        );

    \I__4140\ : InMux
    port map (
            O => \N__26108\,
            I => \N__26105\
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__26105\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI190J_15\
        );

    \I__4138\ : CascadeMux
    port map (
            O => \N__26102\,
            I => \N__26098\
        );

    \I__4137\ : InMux
    port map (
            O => \N__26101\,
            I => \N__26090\
        );

    \I__4136\ : InMux
    port map (
            O => \N__26098\,
            I => \N__26090\
        );

    \I__4135\ : InMux
    port map (
            O => \N__26097\,
            I => \N__26090\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__26090\,
            I => \N__26087\
        );

    \I__4133\ : Span4Mux_v
    port map (
            O => \N__26087\,
            I => \N__26083\
        );

    \I__4132\ : InMux
    port map (
            O => \N__26086\,
            I => \N__26080\
        );

    \I__4131\ : Span4Mux_h
    port map (
            O => \N__26083\,
            I => \N__26077\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__26080\,
            I => \N__26074\
        );

    \I__4129\ : Odrv4
    port map (
            O => \N__26077\,
            I => \current_shift_inst.elapsed_time_ns_phase_20\
        );

    \I__4128\ : Odrv4
    port map (
            O => \N__26074\,
            I => \current_shift_inst.elapsed_time_ns_phase_20\
        );

    \I__4127\ : InMux
    port map (
            O => \N__26069\,
            I => \N__26062\
        );

    \I__4126\ : InMux
    port map (
            O => \N__26068\,
            I => \N__26062\
        );

    \I__4125\ : InMux
    port map (
            O => \N__26067\,
            I => \N__26059\
        );

    \I__4124\ : LocalMux
    port map (
            O => \N__26062\,
            I => \N__26056\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__26059\,
            I => \N__26053\
        );

    \I__4122\ : Span4Mux_v
    port map (
            O => \N__26056\,
            I => \N__26050\
        );

    \I__4121\ : Span4Mux_v
    port map (
            O => \N__26053\,
            I => \N__26044\
        );

    \I__4120\ : Span4Mux_h
    port map (
            O => \N__26050\,
            I => \N__26044\
        );

    \I__4119\ : InMux
    port map (
            O => \N__26049\,
            I => \N__26041\
        );

    \I__4118\ : Span4Mux_h
    port map (
            O => \N__26044\,
            I => \N__26038\
        );

    \I__4117\ : LocalMux
    port map (
            O => \N__26041\,
            I => \N__26035\
        );

    \I__4116\ : Odrv4
    port map (
            O => \N__26038\,
            I => \current_shift_inst.elapsed_time_ns_phase_21\
        );

    \I__4115\ : Odrv4
    port map (
            O => \N__26035\,
            I => \current_shift_inst.elapsed_time_ns_phase_21\
        );

    \I__4114\ : InMux
    port map (
            O => \N__26030\,
            I => \N__26027\
        );

    \I__4113\ : LocalMux
    port map (
            O => \N__26027\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIDR081_20\
        );

    \I__4112\ : CascadeMux
    port map (
            O => \N__26024\,
            I => \N__26020\
        );

    \I__4111\ : InMux
    port map (
            O => \N__26023\,
            I => \N__26012\
        );

    \I__4110\ : InMux
    port map (
            O => \N__26020\,
            I => \N__26012\
        );

    \I__4109\ : InMux
    port map (
            O => \N__26019\,
            I => \N__26012\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__26012\,
            I => \N__26009\
        );

    \I__4107\ : Span4Mux_h
    port map (
            O => \N__26009\,
            I => \N__26006\
        );

    \I__4106\ : Span4Mux_v
    port map (
            O => \N__26006\,
            I => \N__26002\
        );

    \I__4105\ : InMux
    port map (
            O => \N__26005\,
            I => \N__25999\
        );

    \I__4104\ : Odrv4
    port map (
            O => \N__26002\,
            I => \current_shift_inst.elapsed_time_ns_phase_17\
        );

    \I__4103\ : LocalMux
    port map (
            O => \N__25999\,
            I => \current_shift_inst.elapsed_time_ns_phase_17\
        );

    \I__4102\ : CascadeMux
    port map (
            O => \N__25994\,
            I => \N__25991\
        );

    \I__4101\ : InMux
    port map (
            O => \N__25991\,
            I => \N__25984\
        );

    \I__4100\ : InMux
    port map (
            O => \N__25990\,
            I => \N__25984\
        );

    \I__4099\ : InMux
    port map (
            O => \N__25989\,
            I => \N__25981\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__25984\,
            I => \N__25978\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__25981\,
            I => \N__25975\
        );

    \I__4096\ : Span4Mux_h
    port map (
            O => \N__25978\,
            I => \N__25972\
        );

    \I__4095\ : Span12Mux_h
    port map (
            O => \N__25975\,
            I => \N__25968\
        );

    \I__4094\ : Span4Mux_v
    port map (
            O => \N__25972\,
            I => \N__25965\
        );

    \I__4093\ : InMux
    port map (
            O => \N__25971\,
            I => \N__25962\
        );

    \I__4092\ : Odrv12
    port map (
            O => \N__25968\,
            I => \current_shift_inst.elapsed_time_ns_phase_18\
        );

    \I__4091\ : Odrv4
    port map (
            O => \N__25965\,
            I => \current_shift_inst.elapsed_time_ns_phase_18\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__25962\,
            I => \current_shift_inst.elapsed_time_ns_phase_18\
        );

    \I__4089\ : InMux
    port map (
            O => \N__25955\,
            I => \N__25952\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__25952\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIH6661_17\
        );

    \I__4087\ : InMux
    port map (
            O => \N__25949\,
            I => \N__25946\
        );

    \I__4086\ : LocalMux
    port map (
            O => \N__25946\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI7DM51_10\
        );

    \I__4085\ : CascadeMux
    port map (
            O => \N__25943\,
            I => \N__25940\
        );

    \I__4084\ : InMux
    port map (
            O => \N__25940\,
            I => \N__25937\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__25937\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI4H5J_19\
        );

    \I__4082\ : InMux
    port map (
            O => \N__25934\,
            I => \N__25929\
        );

    \I__4081\ : InMux
    port map (
            O => \N__25933\,
            I => \N__25926\
        );

    \I__4080\ : InMux
    port map (
            O => \N__25932\,
            I => \N__25923\
        );

    \I__4079\ : LocalMux
    port map (
            O => \N__25929\,
            I => \N__25918\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__25926\,
            I => \N__25918\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__25923\,
            I => \N__25915\
        );

    \I__4076\ : Span4Mux_v
    port map (
            O => \N__25918\,
            I => \N__25910\
        );

    \I__4075\ : Span4Mux_h
    port map (
            O => \N__25915\,
            I => \N__25910\
        );

    \I__4074\ : Span4Mux_v
    port map (
            O => \N__25910\,
            I => \N__25906\
        );

    \I__4073\ : InMux
    port map (
            O => \N__25909\,
            I => \N__25903\
        );

    \I__4072\ : Odrv4
    port map (
            O => \N__25906\,
            I => \current_shift_inst.elapsed_time_ns_phase_10\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__25903\,
            I => \current_shift_inst.elapsed_time_ns_phase_10\
        );

    \I__4070\ : InMux
    port map (
            O => \N__25898\,
            I => \N__25895\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__25895\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJDBL1_10\
        );

    \I__4068\ : InMux
    port map (
            O => \N__25892\,
            I => \N__25887\
        );

    \I__4067\ : InMux
    port map (
            O => \N__25891\,
            I => \N__25884\
        );

    \I__4066\ : InMux
    port map (
            O => \N__25890\,
            I => \N__25881\
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__25887\,
            I => \N__25877\
        );

    \I__4064\ : LocalMux
    port map (
            O => \N__25884\,
            I => \N__25872\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__25881\,
            I => \N__25872\
        );

    \I__4062\ : CascadeMux
    port map (
            O => \N__25880\,
            I => \N__25869\
        );

    \I__4061\ : Span4Mux_v
    port map (
            O => \N__25877\,
            I => \N__25866\
        );

    \I__4060\ : Span4Mux_h
    port map (
            O => \N__25872\,
            I => \N__25863\
        );

    \I__4059\ : InMux
    port map (
            O => \N__25869\,
            I => \N__25860\
        );

    \I__4058\ : Span4Mux_h
    port map (
            O => \N__25866\,
            I => \N__25855\
        );

    \I__4057\ : Span4Mux_v
    port map (
            O => \N__25863\,
            I => \N__25855\
        );

    \I__4056\ : LocalMux
    port map (
            O => \N__25860\,
            I => \N__25852\
        );

    \I__4055\ : Odrv4
    port map (
            O => \N__25855\,
            I => \current_shift_inst.elapsed_time_ns_phase_7\
        );

    \I__4054\ : Odrv4
    port map (
            O => \N__25852\,
            I => \current_shift_inst.elapsed_time_ns_phase_7\
        );

    \I__4053\ : InMux
    port map (
            O => \N__25847\,
            I => \N__25844\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__25844\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIBBPU1_7\
        );

    \I__4051\ : InMux
    port map (
            O => \N__25841\,
            I => \N__25838\
        );

    \I__4050\ : LocalMux
    port map (
            O => \N__25838\,
            I => \N__25833\
        );

    \I__4049\ : InMux
    port map (
            O => \N__25837\,
            I => \N__25830\
        );

    \I__4048\ : InMux
    port map (
            O => \N__25836\,
            I => \N__25827\
        );

    \I__4047\ : Span4Mux_v
    port map (
            O => \N__25833\,
            I => \N__25821\
        );

    \I__4046\ : LocalMux
    port map (
            O => \N__25830\,
            I => \N__25821\
        );

    \I__4045\ : LocalMux
    port map (
            O => \N__25827\,
            I => \N__25818\
        );

    \I__4044\ : CascadeMux
    port map (
            O => \N__25826\,
            I => \N__25815\
        );

    \I__4043\ : Span4Mux_h
    port map (
            O => \N__25821\,
            I => \N__25812\
        );

    \I__4042\ : Span4Mux_h
    port map (
            O => \N__25818\,
            I => \N__25809\
        );

    \I__4041\ : InMux
    port map (
            O => \N__25815\,
            I => \N__25806\
        );

    \I__4040\ : Span4Mux_v
    port map (
            O => \N__25812\,
            I => \N__25803\
        );

    \I__4039\ : Span4Mux_v
    port map (
            O => \N__25809\,
            I => \N__25798\
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__25806\,
            I => \N__25798\
        );

    \I__4037\ : Odrv4
    port map (
            O => \N__25803\,
            I => \current_shift_inst.elapsed_time_ns_phase_14\
        );

    \I__4036\ : Odrv4
    port map (
            O => \N__25798\,
            I => \current_shift_inst.elapsed_time_ns_phase_14\
        );

    \I__4035\ : CascadeMux
    port map (
            O => \N__25793\,
            I => \N__25790\
        );

    \I__4034\ : InMux
    port map (
            O => \N__25790\,
            I => \N__25787\
        );

    \I__4033\ : LocalMux
    port map (
            O => \N__25787\,
            I => \N__25784\
        );

    \I__4032\ : Odrv4
    port map (
            O => \N__25784\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIU4VI_14\
        );

    \I__4031\ : CascadeMux
    port map (
            O => \N__25781\,
            I => \N__25778\
        );

    \I__4030\ : InMux
    port map (
            O => \N__25778\,
            I => \N__25774\
        );

    \I__4029\ : InMux
    port map (
            O => \N__25777\,
            I => \N__25771\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__25774\,
            I => \N__25765\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__25771\,
            I => \N__25765\
        );

    \I__4026\ : InMux
    port map (
            O => \N__25770\,
            I => \N__25762\
        );

    \I__4025\ : Span4Mux_v
    port map (
            O => \N__25765\,
            I => \N__25757\
        );

    \I__4024\ : LocalMux
    port map (
            O => \N__25762\,
            I => \N__25757\
        );

    \I__4023\ : Span4Mux_h
    port map (
            O => \N__25757\,
            I => \N__25754\
        );

    \I__4022\ : Span4Mux_v
    port map (
            O => \N__25754\,
            I => \N__25750\
        );

    \I__4021\ : InMux
    port map (
            O => \N__25753\,
            I => \N__25747\
        );

    \I__4020\ : Odrv4
    port map (
            O => \N__25750\,
            I => \current_shift_inst.elapsed_time_ns_phase_9\
        );

    \I__4019\ : LocalMux
    port map (
            O => \N__25747\,
            I => \current_shift_inst.elapsed_time_ns_phase_9\
        );

    \I__4018\ : InMux
    port map (
            O => \N__25742\,
            I => \N__25736\
        );

    \I__4017\ : InMux
    port map (
            O => \N__25741\,
            I => \N__25731\
        );

    \I__4016\ : InMux
    port map (
            O => \N__25740\,
            I => \N__25731\
        );

    \I__4015\ : CascadeMux
    port map (
            O => \N__25739\,
            I => \N__25728\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__25736\,
            I => \N__25725\
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__25731\,
            I => \N__25722\
        );

    \I__4012\ : InMux
    port map (
            O => \N__25728\,
            I => \N__25719\
        );

    \I__4011\ : Span12Mux_v
    port map (
            O => \N__25725\,
            I => \N__25716\
        );

    \I__4010\ : Span4Mux_h
    port map (
            O => \N__25722\,
            I => \N__25711\
        );

    \I__4009\ : LocalMux
    port map (
            O => \N__25719\,
            I => \N__25711\
        );

    \I__4008\ : Odrv12
    port map (
            O => \N__25716\,
            I => \current_shift_inst.elapsed_time_ns_phase_8\
        );

    \I__4007\ : Odrv4
    port map (
            O => \N__25711\,
            I => \current_shift_inst.elapsed_time_ns_phase_8\
        );

    \I__4006\ : InMux
    port map (
            O => \N__25706\,
            I => \N__25703\
        );

    \I__4005\ : LocalMux
    port map (
            O => \N__25703\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIO0U12_8\
        );

    \I__4004\ : InMux
    port map (
            O => \N__25700\,
            I => \N__25697\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__25697\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIE6961_18\
        );

    \I__4002\ : InMux
    port map (
            O => \N__25694\,
            I => \N__25691\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__25691\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJ3381_21\
        );

    \I__4000\ : CascadeMux
    port map (
            O => \N__25688\,
            I => \N__25685\
        );

    \I__3999\ : InMux
    port map (
            O => \N__25685\,
            I => \N__25682\
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__25682\,
            I => \N__25677\
        );

    \I__3997\ : InMux
    port map (
            O => \N__25681\,
            I => \N__25671\
        );

    \I__3996\ : InMux
    port map (
            O => \N__25680\,
            I => \N__25671\
        );

    \I__3995\ : Span4Mux_h
    port map (
            O => \N__25677\,
            I => \N__25668\
        );

    \I__3994\ : InMux
    port map (
            O => \N__25676\,
            I => \N__25665\
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__25671\,
            I => \N__25662\
        );

    \I__3992\ : Span4Mux_v
    port map (
            O => \N__25668\,
            I => \N__25657\
        );

    \I__3991\ : LocalMux
    port map (
            O => \N__25665\,
            I => \N__25657\
        );

    \I__3990\ : Odrv4
    port map (
            O => \N__25662\,
            I => \current_shift_inst.elapsed_time_ns_phase_13\
        );

    \I__3989\ : Odrv4
    port map (
            O => \N__25657\,
            I => \current_shift_inst.elapsed_time_ns_phase_13\
        );

    \I__3988\ : CascadeMux
    port map (
            O => \N__25652\,
            I => \N__25649\
        );

    \I__3987\ : InMux
    port map (
            O => \N__25649\,
            I => \N__25646\
        );

    \I__3986\ : LocalMux
    port map (
            O => \N__25646\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP5T51_13\
        );

    \I__3985\ : InMux
    port map (
            O => \N__25643\,
            I => \N__25634\
        );

    \I__3984\ : InMux
    port map (
            O => \N__25642\,
            I => \N__25634\
        );

    \I__3983\ : InMux
    port map (
            O => \N__25641\,
            I => \N__25634\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__25634\,
            I => \N__25631\
        );

    \I__3981\ : Span4Mux_v
    port map (
            O => \N__25631\,
            I => \N__25627\
        );

    \I__3980\ : InMux
    port map (
            O => \N__25630\,
            I => \N__25624\
        );

    \I__3979\ : Span4Mux_h
    port map (
            O => \N__25627\,
            I => \N__25621\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__25624\,
            I => \N__25618\
        );

    \I__3977\ : Odrv4
    port map (
            O => \N__25621\,
            I => \current_shift_inst.elapsed_time_ns_phase_5\
        );

    \I__3976\ : Odrv4
    port map (
            O => \N__25618\,
            I => \current_shift_inst.elapsed_time_ns_phase_5\
        );

    \I__3975\ : CascadeMux
    port map (
            O => \N__25613\,
            I => \N__25609\
        );

    \I__3974\ : CascadeMux
    port map (
            O => \N__25612\,
            I => \N__25606\
        );

    \I__3973\ : InMux
    port map (
            O => \N__25609\,
            I => \N__25602\
        );

    \I__3972\ : InMux
    port map (
            O => \N__25606\,
            I => \N__25597\
        );

    \I__3971\ : InMux
    port map (
            O => \N__25605\,
            I => \N__25597\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__25602\,
            I => \N__25594\
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__25597\,
            I => \N__25591\
        );

    \I__3968\ : Span4Mux_v
    port map (
            O => \N__25594\,
            I => \N__25587\
        );

    \I__3967\ : Span4Mux_h
    port map (
            O => \N__25591\,
            I => \N__25584\
        );

    \I__3966\ : InMux
    port map (
            O => \N__25590\,
            I => \N__25581\
        );

    \I__3965\ : Span4Mux_v
    port map (
            O => \N__25587\,
            I => \N__25578\
        );

    \I__3964\ : Span4Mux_v
    port map (
            O => \N__25584\,
            I => \N__25573\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__25581\,
            I => \N__25573\
        );

    \I__3962\ : Odrv4
    port map (
            O => \N__25578\,
            I => \current_shift_inst.elapsed_time_ns_phase_4\
        );

    \I__3961\ : Odrv4
    port map (
            O => \N__25573\,
            I => \current_shift_inst.elapsed_time_ns_phase_4\
        );

    \I__3960\ : InMux
    port map (
            O => \N__25568\,
            I => \N__25565\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__25565\,
            I => \N__25562\
        );

    \I__3958\ : Odrv4
    port map (
            O => \N__25562\,
            I => \current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0\
        );

    \I__3957\ : CascadeMux
    port map (
            O => \N__25559\,
            I => \N__25556\
        );

    \I__3956\ : InMux
    port map (
            O => \N__25556\,
            I => \N__25553\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__25553\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5M161_15\
        );

    \I__3954\ : CascadeMux
    port map (
            O => \N__25550\,
            I => \N__25547\
        );

    \I__3953\ : InMux
    port map (
            O => \N__25547\,
            I => \N__25544\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__25544\,
            I => \N__25541\
        );

    \I__3951\ : Odrv4
    port map (
            O => \N__25541\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIIKQI_10\
        );

    \I__3950\ : CascadeMux
    port map (
            O => \N__25538\,
            I => \N__25535\
        );

    \I__3949\ : InMux
    port map (
            O => \N__25535\,
            I => \N__25532\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__25532\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI4D1J_16\
        );

    \I__3947\ : InMux
    port map (
            O => \N__25529\,
            I => \N__25526\
        );

    \I__3946\ : LocalMux
    port map (
            O => \N__25526\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIVDV51_14\
        );

    \I__3945\ : CascadeMux
    port map (
            O => \N__25523\,
            I => \N__25520\
        );

    \I__3944\ : InMux
    port map (
            O => \N__25520\,
            I => \N__25517\
        );

    \I__3943\ : LocalMux
    port map (
            O => \N__25517\,
            I => \N__25514\
        );

    \I__3942\ : Odrv4
    port map (
            O => \N__25514\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIK3CV_7\
        );

    \I__3941\ : InMux
    port map (
            O => \N__25511\,
            I => \N__25508\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__25508\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI53NU1_6\
        );

    \I__3939\ : InMux
    port map (
            O => \N__25505\,
            I => \N__25498\
        );

    \I__3938\ : InMux
    port map (
            O => \N__25504\,
            I => \N__25498\
        );

    \I__3937\ : InMux
    port map (
            O => \N__25503\,
            I => \N__25495\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__25498\,
            I => \N__25492\
        );

    \I__3935\ : LocalMux
    port map (
            O => \N__25495\,
            I => \N__25489\
        );

    \I__3934\ : Span4Mux_v
    port map (
            O => \N__25492\,
            I => \N__25483\
        );

    \I__3933\ : Span4Mux_v
    port map (
            O => \N__25489\,
            I => \N__25483\
        );

    \I__3932\ : InMux
    port map (
            O => \N__25488\,
            I => \N__25480\
        );

    \I__3931\ : Span4Mux_h
    port map (
            O => \N__25483\,
            I => \N__25477\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__25480\,
            I => \N__25474\
        );

    \I__3929\ : Odrv4
    port map (
            O => \N__25477\,
            I => \current_shift_inst.elapsed_time_ns_phase_6\
        );

    \I__3928\ : Odrv4
    port map (
            O => \N__25474\,
            I => \current_shift_inst.elapsed_time_ns_phase_6\
        );

    \I__3927\ : CascadeMux
    port map (
            O => \N__25469\,
            I => \N__25466\
        );

    \I__3926\ : InMux
    port map (
            O => \N__25466\,
            I => \N__25463\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__25463\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIHVAV_6\
        );

    \I__3924\ : InMux
    port map (
            O => \N__25460\,
            I => \N__25456\
        );

    \I__3923\ : CascadeMux
    port map (
            O => \N__25459\,
            I => \N__25453\
        );

    \I__3922\ : LocalMux
    port map (
            O => \N__25456\,
            I => \N__25450\
        );

    \I__3921\ : InMux
    port map (
            O => \N__25453\,
            I => \N__25447\
        );

    \I__3920\ : Span4Mux_v
    port map (
            O => \N__25450\,
            I => \N__25442\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__25447\,
            I => \N__25442\
        );

    \I__3918\ : Span4Mux_h
    port map (
            O => \N__25442\,
            I => \N__25439\
        );

    \I__3917\ : Span4Mux_v
    port map (
            O => \N__25439\,
            I => \N__25436\
        );

    \I__3916\ : Odrv4
    port map (
            O => \N__25436\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3\
        );

    \I__3915\ : InMux
    port map (
            O => \N__25433\,
            I => \N__25430\
        );

    \I__3914\ : LocalMux
    port map (
            O => \N__25430\,
            I => \current_shift_inst.un38_control_input_0_cry_4_c_RNOZ0\
        );

    \I__3913\ : CascadeMux
    port map (
            O => \N__25427\,
            I => \N__25424\
        );

    \I__3912\ : InMux
    port map (
            O => \N__25424\,
            I => \N__25421\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__25421\,
            I => \N__25418\
        );

    \I__3910\ : Odrv4
    port map (
            O => \N__25418\,
            I => \current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0Z_0\
        );

    \I__3909\ : InMux
    port map (
            O => \N__25415\,
            I => \N__25412\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__25412\,
            I => \N__25409\
        );

    \I__3907\ : Odrv4
    port map (
            O => \N__25409\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIVQKU1_5\
        );

    \I__3906\ : CascadeMux
    port map (
            O => \N__25406\,
            I => \N__25403\
        );

    \I__3905\ : InMux
    port map (
            O => \N__25403\,
            I => \N__25400\
        );

    \I__3904\ : LocalMux
    port map (
            O => \N__25400\,
            I => \current_shift_inst.elapsed_time_ns_1_RNILORI_11\
        );

    \I__3903\ : CascadeMux
    port map (
            O => \N__25397\,
            I => \N__25394\
        );

    \I__3902\ : InMux
    port map (
            O => \N__25394\,
            I => \N__25391\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__25391\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIN7DV_8\
        );

    \I__3900\ : CascadeMux
    port map (
            O => \N__25388\,
            I => \N__25385\
        );

    \I__3899\ : InMux
    port map (
            O => \N__25385\,
            I => \N__25382\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__25382\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIOSSI_12\
        );

    \I__3897\ : CascadeMux
    port map (
            O => \N__25379\,
            I => \N__25376\
        );

    \I__3896\ : InMux
    port map (
            O => \N__25376\,
            I => \N__25373\
        );

    \I__3895\ : LocalMux
    port map (
            O => \N__25373\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI1PG21_9\
        );

    \I__3894\ : CascadeMux
    port map (
            O => \N__25370\,
            I => \N__25367\
        );

    \I__3893\ : InMux
    port map (
            O => \N__25367\,
            I => \N__25364\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__25364\,
            I => \N__25361\
        );

    \I__3891\ : Odrv4
    port map (
            O => \N__25361\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIER9V_5\
        );

    \I__3890\ : InMux
    port map (
            O => \N__25358\,
            I => \N__25355\
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__25355\,
            I => \N__25352\
        );

    \I__3888\ : Odrv4
    port map (
            O => \N__25352\,
            I => \il_max_comp1_D1\
        );

    \I__3887\ : CascadeMux
    port map (
            O => \N__25349\,
            I => \N__25346\
        );

    \I__3886\ : InMux
    port map (
            O => \N__25346\,
            I => \N__25343\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__25343\,
            I => \N__25340\
        );

    \I__3884\ : Span4Mux_h
    port map (
            O => \N__25340\,
            I => \N__25337\
        );

    \I__3883\ : Odrv4
    port map (
            O => \N__25337\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\
        );

    \I__3882\ : CascadeMux
    port map (
            O => \N__25334\,
            I => \N__25331\
        );

    \I__3881\ : InMux
    port map (
            O => \N__25331\,
            I => \N__25328\
        );

    \I__3880\ : LocalMux
    port map (
            O => \N__25328\,
            I => \N__25325\
        );

    \I__3879\ : Span4Mux_h
    port map (
            O => \N__25325\,
            I => \N__25322\
        );

    \I__3878\ : Span4Mux_h
    port map (
            O => \N__25322\,
            I => \N__25319\
        );

    \I__3877\ : Odrv4
    port map (
            O => \N__25319\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\
        );

    \I__3876\ : CascadeMux
    port map (
            O => \N__25316\,
            I => \N__25313\
        );

    \I__3875\ : InMux
    port map (
            O => \N__25313\,
            I => \N__25310\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__25310\,
            I => \current_shift_inst.z_5_30\
        );

    \I__3873\ : InMux
    port map (
            O => \N__25307\,
            I => \N__25304\
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__25304\,
            I => \current_shift_inst.z_5_cry_30_THRU_CO\
        );

    \I__3871\ : CascadeMux
    port map (
            O => \N__25301\,
            I => \N__25298\
        );

    \I__3870\ : InMux
    port map (
            O => \N__25298\,
            I => \N__25294\
        );

    \I__3869\ : InMux
    port map (
            O => \N__25297\,
            I => \N__25291\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__25294\,
            I => \N__25288\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__25291\,
            I => \N__25285\
        );

    \I__3866\ : Span4Mux_h
    port map (
            O => \N__25288\,
            I => \N__25282\
        );

    \I__3865\ : Odrv12
    port map (
            O => \N__25285\,
            I => \current_shift_inst.elapsed_time_ns_phase_31\
        );

    \I__3864\ : Odrv4
    port map (
            O => \N__25282\,
            I => \current_shift_inst.elapsed_time_ns_phase_31\
        );

    \I__3863\ : InMux
    port map (
            O => \N__25277\,
            I => \current_shift_inst.z_cry_30\
        );

    \I__3862\ : InMux
    port map (
            O => \N__25274\,
            I => \N__25271\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__25271\,
            I => \N__25268\
        );

    \I__3860\ : Odrv4
    port map (
            O => \N__25268\,
            I => \current_shift_inst.stop_timer_s1_RNOZ0Z_0\
        );

    \I__3859\ : InMux
    port map (
            O => \N__25265\,
            I => \N__25260\
        );

    \I__3858\ : InMux
    port map (
            O => \N__25264\,
            I => \N__25257\
        );

    \I__3857\ : InMux
    port map (
            O => \N__25263\,
            I => \N__25254\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__25260\,
            I => \current_shift_inst.start_timer_phaseZ0\
        );

    \I__3855\ : LocalMux
    port map (
            O => \N__25257\,
            I => \current_shift_inst.start_timer_phaseZ0\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__25254\,
            I => \current_shift_inst.start_timer_phaseZ0\
        );

    \I__3853\ : CascadeMux
    port map (
            O => \N__25247\,
            I => \N__25244\
        );

    \I__3852\ : InMux
    port map (
            O => \N__25244\,
            I => \N__25241\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__25241\,
            I => \current_shift_inst.z_5_21\
        );

    \I__3850\ : InMux
    port map (
            O => \N__25238\,
            I => \N__25235\
        );

    \I__3849\ : LocalMux
    port map (
            O => \N__25235\,
            I => \current_shift_inst.z_5_22\
        );

    \I__3848\ : InMux
    port map (
            O => \N__25232\,
            I => \N__25229\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__25229\,
            I => \current_shift_inst.z_5_23\
        );

    \I__3846\ : InMux
    port map (
            O => \N__25226\,
            I => \N__25223\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__25223\,
            I => \N__25220\
        );

    \I__3844\ : Odrv4
    port map (
            O => \N__25220\,
            I => \current_shift_inst.z_5_24\
        );

    \I__3843\ : InMux
    port map (
            O => \N__25217\,
            I => \N__25214\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__25214\,
            I => \current_shift_inst.z_5_25\
        );

    \I__3841\ : InMux
    port map (
            O => \N__25211\,
            I => \N__25208\
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__25208\,
            I => \current_shift_inst.z_5_26\
        );

    \I__3839\ : InMux
    port map (
            O => \N__25205\,
            I => \N__25202\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__25202\,
            I => \current_shift_inst.z_5_27\
        );

    \I__3837\ : InMux
    port map (
            O => \N__25199\,
            I => \N__25196\
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__25196\,
            I => \current_shift_inst.z_5_28\
        );

    \I__3835\ : CascadeMux
    port map (
            O => \N__25193\,
            I => \N__25190\
        );

    \I__3834\ : InMux
    port map (
            O => \N__25190\,
            I => \N__25187\
        );

    \I__3833\ : LocalMux
    port map (
            O => \N__25187\,
            I => \current_shift_inst.z_5_29\
        );

    \I__3832\ : InMux
    port map (
            O => \N__25184\,
            I => \N__25181\
        );

    \I__3831\ : LocalMux
    port map (
            O => \N__25181\,
            I => \current_shift_inst.z_5_13\
        );

    \I__3830\ : InMux
    port map (
            O => \N__25178\,
            I => \N__25175\
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__25175\,
            I => \current_shift_inst.z_5_14\
        );

    \I__3828\ : CascadeMux
    port map (
            O => \N__25172\,
            I => \N__25169\
        );

    \I__3827\ : InMux
    port map (
            O => \N__25169\,
            I => \N__25166\
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__25166\,
            I => \current_shift_inst.z_5_15\
        );

    \I__3825\ : CascadeMux
    port map (
            O => \N__25163\,
            I => \N__25160\
        );

    \I__3824\ : InMux
    port map (
            O => \N__25160\,
            I => \N__25157\
        );

    \I__3823\ : LocalMux
    port map (
            O => \N__25157\,
            I => \N__25154\
        );

    \I__3822\ : Span4Mux_v
    port map (
            O => \N__25154\,
            I => \N__25151\
        );

    \I__3821\ : Odrv4
    port map (
            O => \N__25151\,
            I => \current_shift_inst.z_5_16\
        );

    \I__3820\ : InMux
    port map (
            O => \N__25148\,
            I => \N__25145\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__25145\,
            I => \current_shift_inst.z_5_17\
        );

    \I__3818\ : InMux
    port map (
            O => \N__25142\,
            I => \N__25139\
        );

    \I__3817\ : LocalMux
    port map (
            O => \N__25139\,
            I => \current_shift_inst.z_5_18\
        );

    \I__3816\ : InMux
    port map (
            O => \N__25136\,
            I => \N__25133\
        );

    \I__3815\ : LocalMux
    port map (
            O => \N__25133\,
            I => \current_shift_inst.z_5_19\
        );

    \I__3814\ : InMux
    port map (
            O => \N__25130\,
            I => \N__25127\
        );

    \I__3813\ : LocalMux
    port map (
            O => \N__25127\,
            I => \current_shift_inst.z_5_20\
        );

    \I__3812\ : InMux
    port map (
            O => \N__25124\,
            I => \N__25121\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__25121\,
            I => \current_shift_inst.z_5_5\
        );

    \I__3810\ : InMux
    port map (
            O => \N__25118\,
            I => \N__25115\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__25115\,
            I => \current_shift_inst.z_5_6\
        );

    \I__3808\ : InMux
    port map (
            O => \N__25112\,
            I => \N__25109\
        );

    \I__3807\ : LocalMux
    port map (
            O => \N__25109\,
            I => \current_shift_inst.z_5_7\
        );

    \I__3806\ : InMux
    port map (
            O => \N__25106\,
            I => \N__25103\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__25103\,
            I => \N__25100\
        );

    \I__3804\ : Odrv4
    port map (
            O => \N__25100\,
            I => \current_shift_inst.z_5_8\
        );

    \I__3803\ : InMux
    port map (
            O => \N__25097\,
            I => \N__25094\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__25094\,
            I => \current_shift_inst.z_5_9\
        );

    \I__3801\ : InMux
    port map (
            O => \N__25091\,
            I => \N__25088\
        );

    \I__3800\ : LocalMux
    port map (
            O => \N__25088\,
            I => \current_shift_inst.z_5_10\
        );

    \I__3799\ : InMux
    port map (
            O => \N__25085\,
            I => \N__25082\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__25082\,
            I => \current_shift_inst.z_5_11\
        );

    \I__3797\ : CascadeMux
    port map (
            O => \N__25079\,
            I => \N__25076\
        );

    \I__3796\ : InMux
    port map (
            O => \N__25076\,
            I => \N__25073\
        );

    \I__3795\ : LocalMux
    port map (
            O => \N__25073\,
            I => \current_shift_inst.z_5_12\
        );

    \I__3794\ : InMux
    port map (
            O => \N__25070\,
            I => \N__25067\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__25067\,
            I => \N__25064\
        );

    \I__3792\ : Odrv4
    port map (
            O => \N__25064\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIDS8K_28\
        );

    \I__3791\ : CascadeMux
    port map (
            O => \N__25061\,
            I => \N__25058\
        );

    \I__3790\ : InMux
    port map (
            O => \N__25058\,
            I => \N__25055\
        );

    \I__3789\ : LocalMux
    port map (
            O => \N__25055\,
            I => \N__25052\
        );

    \I__3788\ : Odrv4
    port map (
            O => \N__25052\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIKKJ81_29\
        );

    \I__3787\ : InMux
    port map (
            O => \N__25049\,
            I => \N__25046\
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__25046\,
            I => \current_shift_inst.control_input_1_axb_23\
        );

    \I__3785\ : InMux
    port map (
            O => \N__25043\,
            I => \current_shift_inst.un38_control_input_0_cry_28\
        );

    \I__3784\ : InMux
    port map (
            O => \N__25040\,
            I => \N__25037\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__25037\,
            I => \N__25034\
        );

    \I__3782\ : Span4Mux_v
    port map (
            O => \N__25034\,
            I => \N__25031\
        );

    \I__3781\ : Odrv4
    port map (
            O => \N__25031\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIVQF91_30\
        );

    \I__3780\ : CascadeMux
    port map (
            O => \N__25028\,
            I => \N__25024\
        );

    \I__3779\ : InMux
    port map (
            O => \N__25027\,
            I => \N__25021\
        );

    \I__3778\ : InMux
    port map (
            O => \N__25024\,
            I => \N__25018\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__25021\,
            I => \N__25015\
        );

    \I__3776\ : LocalMux
    port map (
            O => \N__25018\,
            I => \N__25012\
        );

    \I__3775\ : Span4Mux_h
    port map (
            O => \N__25015\,
            I => \N__25009\
        );

    \I__3774\ : Span4Mux_h
    port map (
            O => \N__25012\,
            I => \N__25006\
        );

    \I__3773\ : Odrv4
    port map (
            O => \N__25009\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI7OAK_29\
        );

    \I__3772\ : Odrv4
    port map (
            O => \N__25006\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI7OAK_29\
        );

    \I__3771\ : InMux
    port map (
            O => \N__25001\,
            I => \N__24998\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__24998\,
            I => \current_shift_inst.control_input_1_axb_24\
        );

    \I__3769\ : InMux
    port map (
            O => \N__24995\,
            I => \current_shift_inst.un38_control_input_0_cry_29\
        );

    \I__3768\ : InMux
    port map (
            O => \N__24992\,
            I => \N__24989\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__24989\,
            I => \N__24986\
        );

    \I__3766\ : Span4Mux_h
    port map (
            O => \N__24986\,
            I => \N__24983\
        );

    \I__3765\ : Odrv4
    port map (
            O => \N__24983\,
            I => \current_shift_inst.un38_control_input_0_axb_31\
        );

    \I__3764\ : CascadeMux
    port map (
            O => \N__24980\,
            I => \N__24977\
        );

    \I__3763\ : InMux
    port map (
            O => \N__24977\,
            I => \N__24974\
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__24974\,
            I => \current_shift_inst.control_input_1_cry_24_THRU_CO\
        );

    \I__3761\ : InMux
    port map (
            O => \N__24971\,
            I => \bfn_9_17_0_\
        );

    \I__3760\ : CEMux
    port map (
            O => \N__24968\,
            I => \N__24963\
        );

    \I__3759\ : CEMux
    port map (
            O => \N__24967\,
            I => \N__24960\
        );

    \I__3758\ : CEMux
    port map (
            O => \N__24966\,
            I => \N__24956\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__24963\,
            I => \N__24953\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__24960\,
            I => \N__24949\
        );

    \I__3755\ : CEMux
    port map (
            O => \N__24959\,
            I => \N__24946\
        );

    \I__3754\ : LocalMux
    port map (
            O => \N__24956\,
            I => \N__24941\
        );

    \I__3753\ : Span4Mux_v
    port map (
            O => \N__24953\,
            I => \N__24941\
        );

    \I__3752\ : CEMux
    port map (
            O => \N__24952\,
            I => \N__24938\
        );

    \I__3751\ : Span4Mux_v
    port map (
            O => \N__24949\,
            I => \N__24935\
        );

    \I__3750\ : LocalMux
    port map (
            O => \N__24946\,
            I => \N__24928\
        );

    \I__3749\ : Span4Mux_v
    port map (
            O => \N__24941\,
            I => \N__24928\
        );

    \I__3748\ : LocalMux
    port map (
            O => \N__24938\,
            I => \N__24928\
        );

    \I__3747\ : Odrv4
    port map (
            O => \N__24935\,
            I => \current_shift_inst.phase_valid_RNISLORZ0Z2\
        );

    \I__3746\ : Odrv4
    port map (
            O => \N__24928\,
            I => \current_shift_inst.phase_valid_RNISLORZ0Z2\
        );

    \I__3745\ : CascadeMux
    port map (
            O => \N__24923\,
            I => \N__24920\
        );

    \I__3744\ : InMux
    port map (
            O => \N__24920\,
            I => \N__24917\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__24917\,
            I => \G_406\
        );

    \I__3742\ : InMux
    port map (
            O => \N__24914\,
            I => \N__24910\
        );

    \I__3741\ : InMux
    port map (
            O => \N__24913\,
            I => \N__24904\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__24910\,
            I => \N__24901\
        );

    \I__3739\ : InMux
    port map (
            O => \N__24909\,
            I => \N__24897\
        );

    \I__3738\ : InMux
    port map (
            O => \N__24908\,
            I => \N__24892\
        );

    \I__3737\ : InMux
    port map (
            O => \N__24907\,
            I => \N__24892\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__24904\,
            I => \N__24887\
        );

    \I__3735\ : Span4Mux_h
    port map (
            O => \N__24901\,
            I => \N__24887\
        );

    \I__3734\ : InMux
    port map (
            O => \N__24900\,
            I => \N__24884\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__24897\,
            I => \current_shift_inst.elapsed_time_ns_phase_1\
        );

    \I__3732\ : LocalMux
    port map (
            O => \N__24892\,
            I => \current_shift_inst.elapsed_time_ns_phase_1\
        );

    \I__3731\ : Odrv4
    port map (
            O => \N__24887\,
            I => \current_shift_inst.elapsed_time_ns_phase_1\
        );

    \I__3730\ : LocalMux
    port map (
            O => \N__24884\,
            I => \current_shift_inst.elapsed_time_ns_phase_1\
        );

    \I__3729\ : CascadeMux
    port map (
            O => \N__24875\,
            I => \N__24872\
        );

    \I__3728\ : InMux
    port map (
            O => \N__24872\,
            I => \N__24869\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__24869\,
            I => \G_405\
        );

    \I__3726\ : InMux
    port map (
            O => \N__24866\,
            I => \N__24863\
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__24863\,
            I => \N__24860\
        );

    \I__3724\ : Odrv4
    port map (
            O => \N__24860\,
            I => \current_shift_inst.z_5_2\
        );

    \I__3723\ : CascadeMux
    port map (
            O => \N__24857\,
            I => \N__24854\
        );

    \I__3722\ : InMux
    port map (
            O => \N__24854\,
            I => \N__24851\
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__24851\,
            I => \current_shift_inst.z_5_3\
        );

    \I__3720\ : CascadeMux
    port map (
            O => \N__24848\,
            I => \N__24845\
        );

    \I__3719\ : InMux
    port map (
            O => \N__24845\,
            I => \N__24842\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__24842\,
            I => \current_shift_inst.z_5_4\
        );

    \I__3717\ : InMux
    port map (
            O => \N__24839\,
            I => \N__24836\
        );

    \I__3716\ : LocalMux
    port map (
            O => \N__24836\,
            I => \current_shift_inst.control_input_1_axb_15\
        );

    \I__3715\ : InMux
    port map (
            O => \N__24833\,
            I => \current_shift_inst.un38_control_input_0_cry_20\
        );

    \I__3714\ : InMux
    port map (
            O => \N__24830\,
            I => \N__24827\
        );

    \I__3713\ : LocalMux
    port map (
            O => \N__24827\,
            I => \current_shift_inst.control_input_1_axb_16\
        );

    \I__3712\ : InMux
    port map (
            O => \N__24824\,
            I => \current_shift_inst.un38_control_input_0_cry_21\
        );

    \I__3711\ : InMux
    port map (
            O => \N__24821\,
            I => \N__24818\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__24818\,
            I => \current_shift_inst.control_input_1_axb_17\
        );

    \I__3709\ : InMux
    port map (
            O => \N__24815\,
            I => \bfn_9_16_0_\
        );

    \I__3708\ : InMux
    port map (
            O => \N__24812\,
            I => \N__24809\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__24809\,
            I => \N__24806\
        );

    \I__3706\ : Odrv4
    port map (
            O => \N__24806\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIU73K_23\
        );

    \I__3705\ : CascadeMux
    port map (
            O => \N__24803\,
            I => \N__24800\
        );

    \I__3704\ : InMux
    port map (
            O => \N__24800\,
            I => \N__24797\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__24797\,
            I => \N__24794\
        );

    \I__3702\ : Odrv4
    port map (
            O => \N__24794\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIVJ781_23\
        );

    \I__3701\ : InMux
    port map (
            O => \N__24791\,
            I => \N__24788\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__24788\,
            I => \current_shift_inst.control_input_1_axb_18\
        );

    \I__3699\ : InMux
    port map (
            O => \N__24785\,
            I => \current_shift_inst.un38_control_input_0_cry_23\
        );

    \I__3698\ : InMux
    port map (
            O => \N__24782\,
            I => \N__24779\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__24779\,
            I => \current_shift_inst.control_input_1_axb_19\
        );

    \I__3696\ : InMux
    port map (
            O => \N__24776\,
            I => \current_shift_inst.un38_control_input_0_cry_24\
        );

    \I__3695\ : InMux
    port map (
            O => \N__24773\,
            I => \N__24770\
        );

    \I__3694\ : LocalMux
    port map (
            O => \N__24770\,
            I => \N__24767\
        );

    \I__3693\ : Odrv4
    port map (
            O => \N__24767\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIB4C81_25\
        );

    \I__3692\ : CascadeMux
    port map (
            O => \N__24764\,
            I => \N__24761\
        );

    \I__3691\ : InMux
    port map (
            O => \N__24761\,
            I => \N__24758\
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__24758\,
            I => \N__24755\
        );

    \I__3689\ : Odrv4
    port map (
            O => \N__24755\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI4G5K_25\
        );

    \I__3688\ : InMux
    port map (
            O => \N__24752\,
            I => \N__24749\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__24749\,
            I => \current_shift_inst.control_input_1_axb_20\
        );

    \I__3686\ : InMux
    port map (
            O => \N__24746\,
            I => \current_shift_inst.un38_control_input_0_cry_25\
        );

    \I__3685\ : InMux
    port map (
            O => \N__24743\,
            I => \N__24740\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__24740\,
            I => \current_shift_inst.control_input_1_axb_21\
        );

    \I__3683\ : InMux
    port map (
            O => \N__24737\,
            I => \current_shift_inst.un38_control_input_0_cry_26\
        );

    \I__3682\ : CascadeMux
    port map (
            O => \N__24734\,
            I => \N__24731\
        );

    \I__3681\ : InMux
    port map (
            O => \N__24731\,
            I => \N__24728\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__24728\,
            I => \N__24725\
        );

    \I__3679\ : Odrv4
    port map (
            O => \N__24725\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIAO7K_27\
        );

    \I__3678\ : InMux
    port map (
            O => \N__24722\,
            I => \N__24719\
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__24719\,
            I => \current_shift_inst.control_input_1_axb_22\
        );

    \I__3676\ : InMux
    port map (
            O => \N__24716\,
            I => \current_shift_inst.un38_control_input_0_cry_27\
        );

    \I__3675\ : InMux
    port map (
            O => \N__24713\,
            I => \N__24710\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__24710\,
            I => \current_shift_inst.control_input_1_axb_6\
        );

    \I__3673\ : InMux
    port map (
            O => \N__24707\,
            I => \current_shift_inst.un38_control_input_0_cry_11\
        );

    \I__3672\ : InMux
    port map (
            O => \N__24704\,
            I => \N__24701\
        );

    \I__3671\ : LocalMux
    port map (
            O => \N__24701\,
            I => \N__24698\
        );

    \I__3670\ : Span4Mux_h
    port map (
            O => \N__24698\,
            I => \N__24695\
        );

    \I__3669\ : Odrv4
    port map (
            O => \N__24695\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJTQ51_12\
        );

    \I__3668\ : InMux
    port map (
            O => \N__24692\,
            I => \N__24689\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__24689\,
            I => \current_shift_inst.control_input_1_axb_7\
        );

    \I__3666\ : InMux
    port map (
            O => \N__24686\,
            I => \current_shift_inst.un38_control_input_0_cry_12\
        );

    \I__3665\ : InMux
    port map (
            O => \N__24683\,
            I => \N__24680\
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__24680\,
            I => \N__24677\
        );

    \I__3663\ : Span4Mux_h
    port map (
            O => \N__24677\,
            I => \N__24674\
        );

    \I__3662\ : Odrv4
    port map (
            O => \N__24674\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIR0UI_13\
        );

    \I__3661\ : InMux
    port map (
            O => \N__24671\,
            I => \N__24668\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__24668\,
            I => \current_shift_inst.control_input_1_axb_8\
        );

    \I__3659\ : InMux
    port map (
            O => \N__24665\,
            I => \current_shift_inst.un38_control_input_0_cry_13\
        );

    \I__3658\ : InMux
    port map (
            O => \N__24662\,
            I => \N__24659\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__24659\,
            I => \current_shift_inst.control_input_1_axb_9\
        );

    \I__3656\ : InMux
    port map (
            O => \N__24656\,
            I => \bfn_9_15_0_\
        );

    \I__3655\ : InMux
    port map (
            O => \N__24653\,
            I => \N__24650\
        );

    \I__3654\ : LocalMux
    port map (
            O => \N__24650\,
            I => \current_shift_inst.control_input_1_axb_10\
        );

    \I__3653\ : InMux
    port map (
            O => \N__24647\,
            I => \current_shift_inst.un38_control_input_0_cry_15\
        );

    \I__3652\ : InMux
    port map (
            O => \N__24644\,
            I => \N__24641\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__24641\,
            I => \current_shift_inst.control_input_1_axb_11\
        );

    \I__3650\ : InMux
    port map (
            O => \N__24638\,
            I => \current_shift_inst.un38_control_input_0_cry_16\
        );

    \I__3649\ : InMux
    port map (
            O => \N__24635\,
            I => \N__24632\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__24632\,
            I => \current_shift_inst.control_input_1_axb_12\
        );

    \I__3647\ : InMux
    port map (
            O => \N__24629\,
            I => \current_shift_inst.un38_control_input_0_cry_17\
        );

    \I__3646\ : InMux
    port map (
            O => \N__24626\,
            I => \N__24623\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__24623\,
            I => \current_shift_inst.control_input_1_axb_13\
        );

    \I__3644\ : InMux
    port map (
            O => \N__24620\,
            I => \current_shift_inst.un38_control_input_0_cry_18\
        );

    \I__3643\ : InMux
    port map (
            O => \N__24617\,
            I => \N__24614\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__24614\,
            I => \current_shift_inst.control_input_1_axb_14\
        );

    \I__3641\ : InMux
    port map (
            O => \N__24611\,
            I => \current_shift_inst.un38_control_input_0_cry_19\
        );

    \I__3640\ : InMux
    port map (
            O => \N__24608\,
            I => \N__24605\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__24605\,
            I => \current_shift_inst.control_input_1_axb_0\
        );

    \I__3638\ : InMux
    port map (
            O => \N__24602\,
            I => \current_shift_inst.un38_control_input_0_cry_5\
        );

    \I__3637\ : InMux
    port map (
            O => \N__24599\,
            I => \N__24596\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__24596\,
            I => \current_shift_inst.control_input_1_axb_1\
        );

    \I__3635\ : InMux
    port map (
            O => \N__24593\,
            I => \bfn_9_14_0_\
        );

    \I__3634\ : InMux
    port map (
            O => \N__24590\,
            I => \N__24587\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__24587\,
            I => \current_shift_inst.control_input_1_axb_2\
        );

    \I__3632\ : InMux
    port map (
            O => \N__24584\,
            I => \current_shift_inst.un38_control_input_0_cry_7\
        );

    \I__3631\ : InMux
    port map (
            O => \N__24581\,
            I => \N__24578\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__24578\,
            I => \current_shift_inst.control_input_1_axb_3\
        );

    \I__3629\ : InMux
    port map (
            O => \N__24575\,
            I => \current_shift_inst.un38_control_input_0_cry_8\
        );

    \I__3628\ : InMux
    port map (
            O => \N__24572\,
            I => \N__24569\
        );

    \I__3627\ : LocalMux
    port map (
            O => \N__24569\,
            I => \current_shift_inst.control_input_1_axb_4\
        );

    \I__3626\ : InMux
    port map (
            O => \N__24566\,
            I => \current_shift_inst.un38_control_input_0_cry_9\
        );

    \I__3625\ : InMux
    port map (
            O => \N__24563\,
            I => \N__24560\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__24560\,
            I => \current_shift_inst.control_input_1_axb_5\
        );

    \I__3623\ : InMux
    port map (
            O => \N__24557\,
            I => \current_shift_inst.un38_control_input_0_cry_10\
        );

    \I__3622\ : InMux
    port map (
            O => \N__24554\,
            I => \N__24551\
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__24551\,
            I => \current_shift_inst.z_i_0_31\
        );

    \I__3620\ : CascadeMux
    port map (
            O => \N__24548\,
            I => \N__24545\
        );

    \I__3619\ : InMux
    port map (
            O => \N__24545\,
            I => \N__24542\
        );

    \I__3618\ : LocalMux
    port map (
            O => \N__24542\,
            I => \N__24539\
        );

    \I__3617\ : Span4Mux_v
    port map (
            O => \N__24539\,
            I => \N__24536\
        );

    \I__3616\ : Odrv4
    port map (
            O => \N__24536\,
            I => \current_shift_inst.un38_control_input_0_cry_1_c_RNOZ0\
        );

    \I__3615\ : CascadeMux
    port map (
            O => \N__24533\,
            I => \N__24530\
        );

    \I__3614\ : InMux
    port map (
            O => \N__24530\,
            I => \N__24527\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__24527\,
            I => \N__24524\
        );

    \I__3612\ : Span4Mux_h
    port map (
            O => \N__24524\,
            I => \N__24521\
        );

    \I__3611\ : Odrv4
    port map (
            O => \N__24521\,
            I => \current_shift_inst.un38_control_input_0_cry_2_c_RNOZ0\
        );

    \I__3610\ : InMux
    port map (
            O => \N__24518\,
            I => \N__24515\
        );

    \I__3609\ : LocalMux
    port map (
            O => \N__24515\,
            I => \N__24512\
        );

    \I__3608\ : Span12Mux_v
    port map (
            O => \N__24512\,
            I => \N__24509\
        );

    \I__3607\ : Odrv12
    port map (
            O => \N__24509\,
            I => \current_shift_inst.N_1620_i\
        );

    \I__3606\ : CascadeMux
    port map (
            O => \N__24506\,
            I => \N__24503\
        );

    \I__3605\ : InMux
    port map (
            O => \N__24503\,
            I => \N__24500\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__24500\,
            I => \current_shift_inst.un38_control_input_0_cry_3_c_invZ0\
        );

    \I__3603\ : InMux
    port map (
            O => \N__24497\,
            I => \N__24494\
        );

    \I__3602\ : LocalMux
    port map (
            O => \N__24494\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12\
        );

    \I__3601\ : InMux
    port map (
            O => \N__24491\,
            I => \N__24486\
        );

    \I__3600\ : InMux
    port map (
            O => \N__24490\,
            I => \N__24483\
        );

    \I__3599\ : InMux
    port map (
            O => \N__24489\,
            I => \N__24480\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__24486\,
            I => \N__24477\
        );

    \I__3597\ : LocalMux
    port map (
            O => \N__24483\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__3596\ : LocalMux
    port map (
            O => \N__24480\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__3595\ : Odrv4
    port map (
            O => \N__24477\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__3594\ : InMux
    port map (
            O => \N__24470\,
            I => \N__24465\
        );

    \I__3593\ : InMux
    port map (
            O => \N__24469\,
            I => \N__24462\
        );

    \I__3592\ : InMux
    port map (
            O => \N__24468\,
            I => \N__24459\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__24465\,
            I => \N__24456\
        );

    \I__3590\ : LocalMux
    port map (
            O => \N__24462\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__24459\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__3588\ : Odrv12
    port map (
            O => \N__24456\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__3587\ : InMux
    port map (
            O => \N__24449\,
            I => \N__24446\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__24446\,
            I => \pwm_generator_inst.un1_counterlto2_0\
        );

    \I__3585\ : CascadeMux
    port map (
            O => \N__24443\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_11_cascade_\
        );

    \I__3584\ : InMux
    port map (
            O => \N__24440\,
            I => \N__24437\
        );

    \I__3583\ : LocalMux
    port map (
            O => \N__24437\,
            I => \current_shift_inst.PI_CTRL.N_44\
        );

    \I__3582\ : InMux
    port map (
            O => \N__24434\,
            I => \N__24431\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__24431\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\
        );

    \I__3580\ : InMux
    port map (
            O => \N__24428\,
            I => \N__24425\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__24425\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\
        );

    \I__3578\ : CascadeMux
    port map (
            O => \N__24422\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15_cascade_\
        );

    \I__3577\ : InMux
    port map (
            O => \N__24419\,
            I => \N__24416\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__24416\,
            I => \current_shift_inst.PI_CTRL.N_43\
        );

    \I__3575\ : InMux
    port map (
            O => \N__24413\,
            I => \pwm_generator_inst.counter_cry_8\
        );

    \I__3574\ : InMux
    port map (
            O => \N__24410\,
            I => \N__24406\
        );

    \I__3573\ : InMux
    port map (
            O => \N__24409\,
            I => \N__24402\
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__24406\,
            I => \N__24399\
        );

    \I__3571\ : InMux
    port map (
            O => \N__24405\,
            I => \N__24396\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__24402\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__3569\ : Odrv4
    port map (
            O => \N__24399\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__3568\ : LocalMux
    port map (
            O => \N__24396\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__3567\ : InMux
    port map (
            O => \N__24389\,
            I => \N__24385\
        );

    \I__3566\ : InMux
    port map (
            O => \N__24388\,
            I => \N__24381\
        );

    \I__3565\ : LocalMux
    port map (
            O => \N__24385\,
            I => \N__24378\
        );

    \I__3564\ : InMux
    port map (
            O => \N__24384\,
            I => \N__24375\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__24381\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__3562\ : Odrv4
    port map (
            O => \N__24378\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__24375\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__3560\ : CascadeMux
    port map (
            O => \N__24368\,
            I => \N__24365\
        );

    \I__3559\ : InMux
    port map (
            O => \N__24365\,
            I => \N__24361\
        );

    \I__3558\ : InMux
    port map (
            O => \N__24364\,
            I => \N__24357\
        );

    \I__3557\ : LocalMux
    port map (
            O => \N__24361\,
            I => \N__24354\
        );

    \I__3556\ : InMux
    port map (
            O => \N__24360\,
            I => \N__24351\
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__24357\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__3554\ : Odrv4
    port map (
            O => \N__24354\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__24351\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__3552\ : InMux
    port map (
            O => \N__24344\,
            I => \N__24341\
        );

    \I__3551\ : LocalMux
    port map (
            O => \N__24341\,
            I => \N__24336\
        );

    \I__3550\ : InMux
    port map (
            O => \N__24340\,
            I => \N__24333\
        );

    \I__3549\ : InMux
    port map (
            O => \N__24339\,
            I => \N__24330\
        );

    \I__3548\ : Odrv4
    port map (
            O => \N__24336\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__24333\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__24330\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__3545\ : CascadeMux
    port map (
            O => \N__24323\,
            I => \pwm_generator_inst.un1_counterlt9_cascade_\
        );

    \I__3544\ : InMux
    port map (
            O => \N__24320\,
            I => \N__24317\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__24317\,
            I => \N__24312\
        );

    \I__3542\ : InMux
    port map (
            O => \N__24316\,
            I => \N__24309\
        );

    \I__3541\ : InMux
    port map (
            O => \N__24315\,
            I => \N__24306\
        );

    \I__3540\ : Odrv4
    port map (
            O => \N__24312\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__24309\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__24306\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__3537\ : InMux
    port map (
            O => \N__24299\,
            I => \N__24281\
        );

    \I__3536\ : InMux
    port map (
            O => \N__24298\,
            I => \N__24281\
        );

    \I__3535\ : InMux
    port map (
            O => \N__24297\,
            I => \N__24281\
        );

    \I__3534\ : InMux
    port map (
            O => \N__24296\,
            I => \N__24281\
        );

    \I__3533\ : InMux
    port map (
            O => \N__24295\,
            I => \N__24272\
        );

    \I__3532\ : InMux
    port map (
            O => \N__24294\,
            I => \N__24272\
        );

    \I__3531\ : InMux
    port map (
            O => \N__24293\,
            I => \N__24272\
        );

    \I__3530\ : InMux
    port map (
            O => \N__24292\,
            I => \N__24272\
        );

    \I__3529\ : InMux
    port map (
            O => \N__24291\,
            I => \N__24267\
        );

    \I__3528\ : InMux
    port map (
            O => \N__24290\,
            I => \N__24267\
        );

    \I__3527\ : LocalMux
    port map (
            O => \N__24281\,
            I => \N__24262\
        );

    \I__3526\ : LocalMux
    port map (
            O => \N__24272\,
            I => \N__24262\
        );

    \I__3525\ : LocalMux
    port map (
            O => \N__24267\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__3524\ : Odrv4
    port map (
            O => \N__24262\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__3523\ : InMux
    port map (
            O => \N__24257\,
            I => \N__24252\
        );

    \I__3522\ : InMux
    port map (
            O => \N__24256\,
            I => \N__24249\
        );

    \I__3521\ : InMux
    port map (
            O => \N__24255\,
            I => \N__24246\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__24252\,
            I => \N__24243\
        );

    \I__3519\ : LocalMux
    port map (
            O => \N__24249\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__24246\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__3517\ : Odrv4
    port map (
            O => \N__24243\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__3516\ : InMux
    port map (
            O => \N__24236\,
            I => \N__24231\
        );

    \I__3515\ : InMux
    port map (
            O => \N__24235\,
            I => \N__24228\
        );

    \I__3514\ : InMux
    port map (
            O => \N__24234\,
            I => \N__24225\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__24231\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__24228\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__24225\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__3510\ : InMux
    port map (
            O => \N__24218\,
            I => \N__24214\
        );

    \I__3509\ : InMux
    port map (
            O => \N__24217\,
            I => \N__24210\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__24214\,
            I => \N__24207\
        );

    \I__3507\ : InMux
    port map (
            O => \N__24213\,
            I => \N__24204\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__24210\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__3505\ : Odrv4
    port map (
            O => \N__24207\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__24204\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__3503\ : InMux
    port map (
            O => \N__24197\,
            I => \N__24194\
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__24194\,
            I => \pwm_generator_inst.un1_counterlto9_2\
        );

    \I__3501\ : InMux
    port map (
            O => \N__24191\,
            I => \N__24188\
        );

    \I__3500\ : LocalMux
    port map (
            O => \N__24188\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\
        );

    \I__3499\ : CascadeMux
    port map (
            O => \N__24185\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_\
        );

    \I__3498\ : InMux
    port map (
            O => \N__24182\,
            I => \N__24179\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__24179\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_10\
        );

    \I__3496\ : InMux
    port map (
            O => \N__24176\,
            I => \bfn_9_7_0_\
        );

    \I__3495\ : InMux
    port map (
            O => \N__24173\,
            I => \pwm_generator_inst.counter_cry_0\
        );

    \I__3494\ : InMux
    port map (
            O => \N__24170\,
            I => \pwm_generator_inst.counter_cry_1\
        );

    \I__3493\ : InMux
    port map (
            O => \N__24167\,
            I => \pwm_generator_inst.counter_cry_2\
        );

    \I__3492\ : InMux
    port map (
            O => \N__24164\,
            I => \pwm_generator_inst.counter_cry_3\
        );

    \I__3491\ : InMux
    port map (
            O => \N__24161\,
            I => \pwm_generator_inst.counter_cry_4\
        );

    \I__3490\ : InMux
    port map (
            O => \N__24158\,
            I => \pwm_generator_inst.counter_cry_5\
        );

    \I__3489\ : InMux
    port map (
            O => \N__24155\,
            I => \pwm_generator_inst.counter_cry_6\
        );

    \I__3488\ : InMux
    port map (
            O => \N__24152\,
            I => \bfn_9_8_0_\
        );

    \I__3487\ : CascadeMux
    port map (
            O => \N__24149\,
            I => \N__24145\
        );

    \I__3486\ : CascadeMux
    port map (
            O => \N__24148\,
            I => \N__24142\
        );

    \I__3485\ : InMux
    port map (
            O => \N__24145\,
            I => \N__24139\
        );

    \I__3484\ : InMux
    port map (
            O => \N__24142\,
            I => \N__24136\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__24139\,
            I => \N__24132\
        );

    \I__3482\ : LocalMux
    port map (
            O => \N__24136\,
            I => \N__24129\
        );

    \I__3481\ : InMux
    port map (
            O => \N__24135\,
            I => \N__24126\
        );

    \I__3480\ : Span4Mux_h
    port map (
            O => \N__24132\,
            I => \N__24123\
        );

    \I__3479\ : Odrv4
    port map (
            O => \N__24129\,
            I => \current_shift_inst.timer_phase.counterZ0Z_25\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__24126\,
            I => \current_shift_inst.timer_phase.counterZ0Z_25\
        );

    \I__3477\ : Odrv4
    port map (
            O => \N__24123\,
            I => \current_shift_inst.timer_phase.counterZ0Z_25\
        );

    \I__3476\ : InMux
    port map (
            O => \N__24116\,
            I => \current_shift_inst.timer_phase.counter_cry_24\
        );

    \I__3475\ : CascadeMux
    port map (
            O => \N__24113\,
            I => \N__24109\
        );

    \I__3474\ : InMux
    port map (
            O => \N__24112\,
            I => \N__24105\
        );

    \I__3473\ : InMux
    port map (
            O => \N__24109\,
            I => \N__24102\
        );

    \I__3472\ : InMux
    port map (
            O => \N__24108\,
            I => \N__24099\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__24105\,
            I => \N__24094\
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__24102\,
            I => \N__24094\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__24099\,
            I => \N__24089\
        );

    \I__3468\ : Span4Mux_v
    port map (
            O => \N__24094\,
            I => \N__24089\
        );

    \I__3467\ : Odrv4
    port map (
            O => \N__24089\,
            I => \current_shift_inst.timer_phase.counterZ0Z_26\
        );

    \I__3466\ : InMux
    port map (
            O => \N__24086\,
            I => \current_shift_inst.timer_phase.counter_cry_25\
        );

    \I__3465\ : InMux
    port map (
            O => \N__24083\,
            I => \N__24076\
        );

    \I__3464\ : InMux
    port map (
            O => \N__24082\,
            I => \N__24076\
        );

    \I__3463\ : InMux
    port map (
            O => \N__24081\,
            I => \N__24073\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__24076\,
            I => \N__24070\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__24073\,
            I => \current_shift_inst.timer_phase.counterZ0Z_27\
        );

    \I__3460\ : Odrv4
    port map (
            O => \N__24070\,
            I => \current_shift_inst.timer_phase.counterZ0Z_27\
        );

    \I__3459\ : InMux
    port map (
            O => \N__24065\,
            I => \current_shift_inst.timer_phase.counter_cry_26\
        );

    \I__3458\ : CascadeMux
    port map (
            O => \N__24062\,
            I => \N__24059\
        );

    \I__3457\ : InMux
    port map (
            O => \N__24059\,
            I => \N__24055\
        );

    \I__3456\ : InMux
    port map (
            O => \N__24058\,
            I => \N__24052\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__24055\,
            I => \N__24049\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__24052\,
            I => \current_shift_inst.timer_phase.counterZ0Z_28\
        );

    \I__3453\ : Odrv4
    port map (
            O => \N__24049\,
            I => \current_shift_inst.timer_phase.counterZ0Z_28\
        );

    \I__3452\ : InMux
    port map (
            O => \N__24044\,
            I => \current_shift_inst.timer_phase.counter_cry_27\
        );

    \I__3451\ : InMux
    port map (
            O => \N__24041\,
            I => \current_shift_inst.timer_phase.counter_cry_28\
        );

    \I__3450\ : CascadeMux
    port map (
            O => \N__24038\,
            I => \N__24035\
        );

    \I__3449\ : InMux
    port map (
            O => \N__24035\,
            I => \N__24031\
        );

    \I__3448\ : InMux
    port map (
            O => \N__24034\,
            I => \N__24028\
        );

    \I__3447\ : LocalMux
    port map (
            O => \N__24031\,
            I => \N__24025\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__24028\,
            I => \current_shift_inst.timer_phase.counterZ0Z_29\
        );

    \I__3445\ : Odrv4
    port map (
            O => \N__24025\,
            I => \current_shift_inst.timer_phase.counterZ0Z_29\
        );

    \I__3444\ : IoInMux
    port map (
            O => \N__24020\,
            I => \N__24017\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__24017\,
            I => \N__24014\
        );

    \I__3442\ : Span4Mux_s1_v
    port map (
            O => \N__24014\,
            I => \N__24011\
        );

    \I__3441\ : Span4Mux_v
    port map (
            O => \N__24011\,
            I => \N__24008\
        );

    \I__3440\ : Odrv4
    port map (
            O => \N__24008\,
            I => \current_shift_inst.timer_s1.N_187_i\
        );

    \I__3439\ : CEMux
    port map (
            O => \N__24005\,
            I => \N__24002\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__24002\,
            I => \N__23997\
        );

    \I__3437\ : CEMux
    port map (
            O => \N__24001\,
            I => \N__23994\
        );

    \I__3436\ : CEMux
    port map (
            O => \N__24000\,
            I => \N__23991\
        );

    \I__3435\ : Span4Mux_h
    port map (
            O => \N__23997\,
            I => \N__23986\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__23994\,
            I => \N__23986\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__23991\,
            I => \N__23982\
        );

    \I__3432\ : Sp12to4
    port map (
            O => \N__23986\,
            I => \N__23979\
        );

    \I__3431\ : CEMux
    port map (
            O => \N__23985\,
            I => \N__23976\
        );

    \I__3430\ : Odrv12
    port map (
            O => \N__23982\,
            I => \current_shift_inst.timer_phase.N_193_i\
        );

    \I__3429\ : Odrv12
    port map (
            O => \N__23979\,
            I => \current_shift_inst.timer_phase.N_193_i\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__23976\,
            I => \current_shift_inst.timer_phase.N_193_i\
        );

    \I__3427\ : InMux
    port map (
            O => \N__23969\,
            I => \N__23931\
        );

    \I__3426\ : InMux
    port map (
            O => \N__23968\,
            I => \N__23931\
        );

    \I__3425\ : InMux
    port map (
            O => \N__23967\,
            I => \N__23931\
        );

    \I__3424\ : InMux
    port map (
            O => \N__23966\,
            I => \N__23931\
        );

    \I__3423\ : InMux
    port map (
            O => \N__23965\,
            I => \N__23922\
        );

    \I__3422\ : InMux
    port map (
            O => \N__23964\,
            I => \N__23922\
        );

    \I__3421\ : InMux
    port map (
            O => \N__23963\,
            I => \N__23922\
        );

    \I__3420\ : InMux
    port map (
            O => \N__23962\,
            I => \N__23922\
        );

    \I__3419\ : InMux
    port map (
            O => \N__23961\,
            I => \N__23913\
        );

    \I__3418\ : InMux
    port map (
            O => \N__23960\,
            I => \N__23913\
        );

    \I__3417\ : InMux
    port map (
            O => \N__23959\,
            I => \N__23913\
        );

    \I__3416\ : InMux
    port map (
            O => \N__23958\,
            I => \N__23913\
        );

    \I__3415\ : InMux
    port map (
            O => \N__23957\,
            I => \N__23904\
        );

    \I__3414\ : InMux
    port map (
            O => \N__23956\,
            I => \N__23904\
        );

    \I__3413\ : InMux
    port map (
            O => \N__23955\,
            I => \N__23904\
        );

    \I__3412\ : InMux
    port map (
            O => \N__23954\,
            I => \N__23904\
        );

    \I__3411\ : InMux
    port map (
            O => \N__23953\,
            I => \N__23895\
        );

    \I__3410\ : InMux
    port map (
            O => \N__23952\,
            I => \N__23895\
        );

    \I__3409\ : InMux
    port map (
            O => \N__23951\,
            I => \N__23895\
        );

    \I__3408\ : InMux
    port map (
            O => \N__23950\,
            I => \N__23895\
        );

    \I__3407\ : InMux
    port map (
            O => \N__23949\,
            I => \N__23886\
        );

    \I__3406\ : InMux
    port map (
            O => \N__23948\,
            I => \N__23886\
        );

    \I__3405\ : InMux
    port map (
            O => \N__23947\,
            I => \N__23886\
        );

    \I__3404\ : InMux
    port map (
            O => \N__23946\,
            I => \N__23886\
        );

    \I__3403\ : InMux
    port map (
            O => \N__23945\,
            I => \N__23881\
        );

    \I__3402\ : InMux
    port map (
            O => \N__23944\,
            I => \N__23881\
        );

    \I__3401\ : InMux
    port map (
            O => \N__23943\,
            I => \N__23872\
        );

    \I__3400\ : InMux
    port map (
            O => \N__23942\,
            I => \N__23872\
        );

    \I__3399\ : InMux
    port map (
            O => \N__23941\,
            I => \N__23872\
        );

    \I__3398\ : InMux
    port map (
            O => \N__23940\,
            I => \N__23872\
        );

    \I__3397\ : LocalMux
    port map (
            O => \N__23931\,
            I => \N__23867\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__23922\,
            I => \N__23867\
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__23913\,
            I => \N__23858\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__23904\,
            I => \N__23858\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__23895\,
            I => \N__23858\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__23886\,
            I => \N__23858\
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__23881\,
            I => \current_shift_inst.timer_phase.running_i\
        );

    \I__3390\ : LocalMux
    port map (
            O => \N__23872\,
            I => \current_shift_inst.timer_phase.running_i\
        );

    \I__3389\ : Odrv4
    port map (
            O => \N__23867\,
            I => \current_shift_inst.timer_phase.running_i\
        );

    \I__3388\ : Odrv12
    port map (
            O => \N__23858\,
            I => \current_shift_inst.timer_phase.running_i\
        );

    \I__3387\ : InMux
    port map (
            O => \N__23849\,
            I => \N__23846\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__23846\,
            I => \N__23843\
        );

    \I__3385\ : Span4Mux_h
    port map (
            O => \N__23843\,
            I => \N__23840\
        );

    \I__3384\ : Odrv4
    port map (
            O => \N__23840\,
            I => il_max_comp1_c
        );

    \I__3383\ : CascadeMux
    port map (
            O => \N__23837\,
            I => \N__23833\
        );

    \I__3382\ : CascadeMux
    port map (
            O => \N__23836\,
            I => \N__23830\
        );

    \I__3381\ : InMux
    port map (
            O => \N__23833\,
            I => \N__23827\
        );

    \I__3380\ : InMux
    port map (
            O => \N__23830\,
            I => \N__23823\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__23827\,
            I => \N__23820\
        );

    \I__3378\ : InMux
    port map (
            O => \N__23826\,
            I => \N__23817\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__23823\,
            I => \N__23812\
        );

    \I__3376\ : Span4Mux_h
    port map (
            O => \N__23820\,
            I => \N__23812\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__23817\,
            I => \current_shift_inst.timer_phase.counterZ0Z_17\
        );

    \I__3374\ : Odrv4
    port map (
            O => \N__23812\,
            I => \current_shift_inst.timer_phase.counterZ0Z_17\
        );

    \I__3373\ : InMux
    port map (
            O => \N__23807\,
            I => \current_shift_inst.timer_phase.counter_cry_16\
        );

    \I__3372\ : CascadeMux
    port map (
            O => \N__23804\,
            I => \N__23801\
        );

    \I__3371\ : InMux
    port map (
            O => \N__23801\,
            I => \N__23796\
        );

    \I__3370\ : InMux
    port map (
            O => \N__23800\,
            I => \N__23793\
        );

    \I__3369\ : InMux
    port map (
            O => \N__23799\,
            I => \N__23790\
        );

    \I__3368\ : LocalMux
    port map (
            O => \N__23796\,
            I => \N__23787\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__23793\,
            I => \N__23784\
        );

    \I__3366\ : LocalMux
    port map (
            O => \N__23790\,
            I => \N__23779\
        );

    \I__3365\ : Span4Mux_v
    port map (
            O => \N__23787\,
            I => \N__23779\
        );

    \I__3364\ : Odrv4
    port map (
            O => \N__23784\,
            I => \current_shift_inst.timer_phase.counterZ0Z_18\
        );

    \I__3363\ : Odrv4
    port map (
            O => \N__23779\,
            I => \current_shift_inst.timer_phase.counterZ0Z_18\
        );

    \I__3362\ : InMux
    port map (
            O => \N__23774\,
            I => \current_shift_inst.timer_phase.counter_cry_17\
        );

    \I__3361\ : InMux
    port map (
            O => \N__23771\,
            I => \N__23764\
        );

    \I__3360\ : InMux
    port map (
            O => \N__23770\,
            I => \N__23764\
        );

    \I__3359\ : InMux
    port map (
            O => \N__23769\,
            I => \N__23761\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__23764\,
            I => \N__23758\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__23761\,
            I => \N__23753\
        );

    \I__3356\ : Span4Mux_v
    port map (
            O => \N__23758\,
            I => \N__23753\
        );

    \I__3355\ : Odrv4
    port map (
            O => \N__23753\,
            I => \current_shift_inst.timer_phase.counterZ0Z_19\
        );

    \I__3354\ : InMux
    port map (
            O => \N__23750\,
            I => \current_shift_inst.timer_phase.counter_cry_18\
        );

    \I__3353\ : CascadeMux
    port map (
            O => \N__23747\,
            I => \N__23743\
        );

    \I__3352\ : CascadeMux
    port map (
            O => \N__23746\,
            I => \N__23740\
        );

    \I__3351\ : InMux
    port map (
            O => \N__23743\,
            I => \N__23735\
        );

    \I__3350\ : InMux
    port map (
            O => \N__23740\,
            I => \N__23735\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__23735\,
            I => \N__23731\
        );

    \I__3348\ : InMux
    port map (
            O => \N__23734\,
            I => \N__23728\
        );

    \I__3347\ : Span4Mux_h
    port map (
            O => \N__23731\,
            I => \N__23725\
        );

    \I__3346\ : LocalMux
    port map (
            O => \N__23728\,
            I => \current_shift_inst.timer_phase.counterZ0Z_20\
        );

    \I__3345\ : Odrv4
    port map (
            O => \N__23725\,
            I => \current_shift_inst.timer_phase.counterZ0Z_20\
        );

    \I__3344\ : InMux
    port map (
            O => \N__23720\,
            I => \current_shift_inst.timer_phase.counter_cry_19\
        );

    \I__3343\ : CascadeMux
    port map (
            O => \N__23717\,
            I => \N__23713\
        );

    \I__3342\ : CascadeMux
    port map (
            O => \N__23716\,
            I => \N__23710\
        );

    \I__3341\ : InMux
    port map (
            O => \N__23713\,
            I => \N__23705\
        );

    \I__3340\ : InMux
    port map (
            O => \N__23710\,
            I => \N__23705\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__23705\,
            I => \N__23701\
        );

    \I__3338\ : InMux
    port map (
            O => \N__23704\,
            I => \N__23698\
        );

    \I__3337\ : Span4Mux_h
    port map (
            O => \N__23701\,
            I => \N__23695\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__23698\,
            I => \current_shift_inst.timer_phase.counterZ0Z_21\
        );

    \I__3335\ : Odrv4
    port map (
            O => \N__23695\,
            I => \current_shift_inst.timer_phase.counterZ0Z_21\
        );

    \I__3334\ : InMux
    port map (
            O => \N__23690\,
            I => \current_shift_inst.timer_phase.counter_cry_20\
        );

    \I__3333\ : InMux
    port map (
            O => \N__23687\,
            I => \N__23681\
        );

    \I__3332\ : InMux
    port map (
            O => \N__23686\,
            I => \N__23681\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__23681\,
            I => \N__23677\
        );

    \I__3330\ : InMux
    port map (
            O => \N__23680\,
            I => \N__23674\
        );

    \I__3329\ : Span4Mux_h
    port map (
            O => \N__23677\,
            I => \N__23671\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__23674\,
            I => \current_shift_inst.timer_phase.counterZ0Z_22\
        );

    \I__3327\ : Odrv4
    port map (
            O => \N__23671\,
            I => \current_shift_inst.timer_phase.counterZ0Z_22\
        );

    \I__3326\ : InMux
    port map (
            O => \N__23666\,
            I => \current_shift_inst.timer_phase.counter_cry_21\
        );

    \I__3325\ : InMux
    port map (
            O => \N__23663\,
            I => \N__23656\
        );

    \I__3324\ : InMux
    port map (
            O => \N__23662\,
            I => \N__23656\
        );

    \I__3323\ : InMux
    port map (
            O => \N__23661\,
            I => \N__23653\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__23656\,
            I => \N__23650\
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__23653\,
            I => \current_shift_inst.timer_phase.counterZ0Z_23\
        );

    \I__3320\ : Odrv4
    port map (
            O => \N__23650\,
            I => \current_shift_inst.timer_phase.counterZ0Z_23\
        );

    \I__3319\ : InMux
    port map (
            O => \N__23645\,
            I => \current_shift_inst.timer_phase.counter_cry_22\
        );

    \I__3318\ : CascadeMux
    port map (
            O => \N__23642\,
            I => \N__23639\
        );

    \I__3317\ : InMux
    port map (
            O => \N__23639\,
            I => \N__23635\
        );

    \I__3316\ : InMux
    port map (
            O => \N__23638\,
            I => \N__23631\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__23635\,
            I => \N__23628\
        );

    \I__3314\ : InMux
    port map (
            O => \N__23634\,
            I => \N__23625\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__23631\,
            I => \N__23620\
        );

    \I__3312\ : Span4Mux_h
    port map (
            O => \N__23628\,
            I => \N__23620\
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__23625\,
            I => \current_shift_inst.timer_phase.counterZ0Z_24\
        );

    \I__3310\ : Odrv4
    port map (
            O => \N__23620\,
            I => \current_shift_inst.timer_phase.counterZ0Z_24\
        );

    \I__3309\ : InMux
    port map (
            O => \N__23615\,
            I => \bfn_8_24_0_\
        );

    \I__3308\ : CascadeMux
    port map (
            O => \N__23612\,
            I => \N__23608\
        );

    \I__3307\ : CascadeMux
    port map (
            O => \N__23611\,
            I => \N__23605\
        );

    \I__3306\ : InMux
    port map (
            O => \N__23608\,
            I => \N__23602\
        );

    \I__3305\ : InMux
    port map (
            O => \N__23605\,
            I => \N__23598\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__23602\,
            I => \N__23595\
        );

    \I__3303\ : InMux
    port map (
            O => \N__23601\,
            I => \N__23592\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__23598\,
            I => \N__23589\
        );

    \I__3301\ : Span4Mux_h
    port map (
            O => \N__23595\,
            I => \N__23586\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__23592\,
            I => \current_shift_inst.timer_phase.counterZ0Z_8\
        );

    \I__3299\ : Odrv4
    port map (
            O => \N__23589\,
            I => \current_shift_inst.timer_phase.counterZ0Z_8\
        );

    \I__3298\ : Odrv4
    port map (
            O => \N__23586\,
            I => \current_shift_inst.timer_phase.counterZ0Z_8\
        );

    \I__3297\ : InMux
    port map (
            O => \N__23579\,
            I => \bfn_8_22_0_\
        );

    \I__3296\ : CascadeMux
    port map (
            O => \N__23576\,
            I => \N__23572\
        );

    \I__3295\ : InMux
    port map (
            O => \N__23575\,
            I => \N__23568\
        );

    \I__3294\ : InMux
    port map (
            O => \N__23572\,
            I => \N__23565\
        );

    \I__3293\ : InMux
    port map (
            O => \N__23571\,
            I => \N__23562\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__23568\,
            I => \N__23557\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__23565\,
            I => \N__23557\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__23562\,
            I => \current_shift_inst.timer_phase.counterZ0Z_9\
        );

    \I__3289\ : Odrv4
    port map (
            O => \N__23557\,
            I => \current_shift_inst.timer_phase.counterZ0Z_9\
        );

    \I__3288\ : InMux
    port map (
            O => \N__23552\,
            I => \current_shift_inst.timer_phase.counter_cry_8\
        );

    \I__3287\ : InMux
    port map (
            O => \N__23549\,
            I => \N__23542\
        );

    \I__3286\ : InMux
    port map (
            O => \N__23548\,
            I => \N__23542\
        );

    \I__3285\ : InMux
    port map (
            O => \N__23547\,
            I => \N__23539\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__23542\,
            I => \N__23536\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__23539\,
            I => \current_shift_inst.timer_phase.counterZ0Z_10\
        );

    \I__3282\ : Odrv4
    port map (
            O => \N__23536\,
            I => \current_shift_inst.timer_phase.counterZ0Z_10\
        );

    \I__3281\ : InMux
    port map (
            O => \N__23531\,
            I => \current_shift_inst.timer_phase.counter_cry_9\
        );

    \I__3280\ : CascadeMux
    port map (
            O => \N__23528\,
            I => \N__23524\
        );

    \I__3279\ : CascadeMux
    port map (
            O => \N__23527\,
            I => \N__23521\
        );

    \I__3278\ : InMux
    port map (
            O => \N__23524\,
            I => \N__23515\
        );

    \I__3277\ : InMux
    port map (
            O => \N__23521\,
            I => \N__23515\
        );

    \I__3276\ : InMux
    port map (
            O => \N__23520\,
            I => \N__23512\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__23515\,
            I => \N__23509\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__23512\,
            I => \current_shift_inst.timer_phase.counterZ0Z_11\
        );

    \I__3273\ : Odrv4
    port map (
            O => \N__23509\,
            I => \current_shift_inst.timer_phase.counterZ0Z_11\
        );

    \I__3272\ : InMux
    port map (
            O => \N__23504\,
            I => \current_shift_inst.timer_phase.counter_cry_10\
        );

    \I__3271\ : CascadeMux
    port map (
            O => \N__23501\,
            I => \N__23497\
        );

    \I__3270\ : CascadeMux
    port map (
            O => \N__23500\,
            I => \N__23494\
        );

    \I__3269\ : InMux
    port map (
            O => \N__23497\,
            I => \N__23489\
        );

    \I__3268\ : InMux
    port map (
            O => \N__23494\,
            I => \N__23489\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__23489\,
            I => \N__23485\
        );

    \I__3266\ : InMux
    port map (
            O => \N__23488\,
            I => \N__23482\
        );

    \I__3265\ : Span4Mux_h
    port map (
            O => \N__23485\,
            I => \N__23479\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__23482\,
            I => \current_shift_inst.timer_phase.counterZ0Z_12\
        );

    \I__3263\ : Odrv4
    port map (
            O => \N__23479\,
            I => \current_shift_inst.timer_phase.counterZ0Z_12\
        );

    \I__3262\ : InMux
    port map (
            O => \N__23474\,
            I => \current_shift_inst.timer_phase.counter_cry_11\
        );

    \I__3261\ : CascadeMux
    port map (
            O => \N__23471\,
            I => \N__23468\
        );

    \I__3260\ : InMux
    port map (
            O => \N__23468\,
            I => \N__23464\
        );

    \I__3259\ : InMux
    port map (
            O => \N__23467\,
            I => \N__23461\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__23464\,
            I => \N__23455\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__23461\,
            I => \N__23455\
        );

    \I__3256\ : InMux
    port map (
            O => \N__23460\,
            I => \N__23452\
        );

    \I__3255\ : Span4Mux_h
    port map (
            O => \N__23455\,
            I => \N__23449\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__23452\,
            I => \current_shift_inst.timer_phase.counterZ0Z_13\
        );

    \I__3253\ : Odrv4
    port map (
            O => \N__23449\,
            I => \current_shift_inst.timer_phase.counterZ0Z_13\
        );

    \I__3252\ : InMux
    port map (
            O => \N__23444\,
            I => \current_shift_inst.timer_phase.counter_cry_12\
        );

    \I__3251\ : InMux
    port map (
            O => \N__23441\,
            I => \N__23435\
        );

    \I__3250\ : InMux
    port map (
            O => \N__23440\,
            I => \N__23435\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__23435\,
            I => \N__23431\
        );

    \I__3248\ : InMux
    port map (
            O => \N__23434\,
            I => \N__23428\
        );

    \I__3247\ : Span4Mux_h
    port map (
            O => \N__23431\,
            I => \N__23425\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__23428\,
            I => \current_shift_inst.timer_phase.counterZ0Z_14\
        );

    \I__3245\ : Odrv4
    port map (
            O => \N__23425\,
            I => \current_shift_inst.timer_phase.counterZ0Z_14\
        );

    \I__3244\ : InMux
    port map (
            O => \N__23420\,
            I => \current_shift_inst.timer_phase.counter_cry_13\
        );

    \I__3243\ : InMux
    port map (
            O => \N__23417\,
            I => \N__23410\
        );

    \I__3242\ : InMux
    port map (
            O => \N__23416\,
            I => \N__23410\
        );

    \I__3241\ : InMux
    port map (
            O => \N__23415\,
            I => \N__23407\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__23410\,
            I => \N__23404\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__23407\,
            I => \current_shift_inst.timer_phase.counterZ0Z_15\
        );

    \I__3238\ : Odrv4
    port map (
            O => \N__23404\,
            I => \current_shift_inst.timer_phase.counterZ0Z_15\
        );

    \I__3237\ : InMux
    port map (
            O => \N__23399\,
            I => \current_shift_inst.timer_phase.counter_cry_14\
        );

    \I__3236\ : CascadeMux
    port map (
            O => \N__23396\,
            I => \N__23393\
        );

    \I__3235\ : InMux
    port map (
            O => \N__23393\,
            I => \N__23389\
        );

    \I__3234\ : InMux
    port map (
            O => \N__23392\,
            I => \N__23385\
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__23389\,
            I => \N__23382\
        );

    \I__3232\ : InMux
    port map (
            O => \N__23388\,
            I => \N__23379\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__23385\,
            I => \N__23374\
        );

    \I__3230\ : Span4Mux_h
    port map (
            O => \N__23382\,
            I => \N__23374\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__23379\,
            I => \current_shift_inst.timer_phase.counterZ0Z_16\
        );

    \I__3228\ : Odrv4
    port map (
            O => \N__23374\,
            I => \current_shift_inst.timer_phase.counterZ0Z_16\
        );

    \I__3227\ : InMux
    port map (
            O => \N__23369\,
            I => \bfn_8_23_0_\
        );

    \I__3226\ : InMux
    port map (
            O => \N__23366\,
            I => \N__23363\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__23363\,
            I => \N__23359\
        );

    \I__3224\ : InMux
    port map (
            O => \N__23362\,
            I => \N__23356\
        );

    \I__3223\ : Span4Mux_v
    port map (
            O => \N__23359\,
            I => \N__23350\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__23356\,
            I => \N__23350\
        );

    \I__3221\ : InMux
    port map (
            O => \N__23355\,
            I => \N__23347\
        );

    \I__3220\ : Odrv4
    port map (
            O => \N__23350\,
            I => \current_shift_inst.timer_phase.counterZ0Z_0\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__23347\,
            I => \current_shift_inst.timer_phase.counterZ0Z_0\
        );

    \I__3218\ : InMux
    port map (
            O => \N__23342\,
            I => \bfn_8_21_0_\
        );

    \I__3217\ : InMux
    port map (
            O => \N__23339\,
            I => \N__23336\
        );

    \I__3216\ : LocalMux
    port map (
            O => \N__23336\,
            I => \N__23332\
        );

    \I__3215\ : InMux
    port map (
            O => \N__23335\,
            I => \N__23329\
        );

    \I__3214\ : Span4Mux_h
    port map (
            O => \N__23332\,
            I => \N__23323\
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__23329\,
            I => \N__23323\
        );

    \I__3212\ : InMux
    port map (
            O => \N__23328\,
            I => \N__23320\
        );

    \I__3211\ : Odrv4
    port map (
            O => \N__23323\,
            I => \current_shift_inst.timer_phase.counterZ0Z_1\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__23320\,
            I => \current_shift_inst.timer_phase.counterZ0Z_1\
        );

    \I__3209\ : InMux
    port map (
            O => \N__23315\,
            I => \current_shift_inst.timer_phase.counter_cry_0\
        );

    \I__3208\ : CascadeMux
    port map (
            O => \N__23312\,
            I => \N__23308\
        );

    \I__3207\ : InMux
    port map (
            O => \N__23311\,
            I => \N__23304\
        );

    \I__3206\ : InMux
    port map (
            O => \N__23308\,
            I => \N__23301\
        );

    \I__3205\ : InMux
    port map (
            O => \N__23307\,
            I => \N__23298\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__23304\,
            I => \N__23293\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__23301\,
            I => \N__23293\
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__23298\,
            I => \N__23288\
        );

    \I__3201\ : Span4Mux_v
    port map (
            O => \N__23293\,
            I => \N__23288\
        );

    \I__3200\ : Odrv4
    port map (
            O => \N__23288\,
            I => \current_shift_inst.timer_phase.counterZ0Z_2\
        );

    \I__3199\ : InMux
    port map (
            O => \N__23285\,
            I => \current_shift_inst.timer_phase.counter_cry_1\
        );

    \I__3198\ : CascadeMux
    port map (
            O => \N__23282\,
            I => \N__23278\
        );

    \I__3197\ : CascadeMux
    port map (
            O => \N__23281\,
            I => \N__23275\
        );

    \I__3196\ : InMux
    port map (
            O => \N__23278\,
            I => \N__23269\
        );

    \I__3195\ : InMux
    port map (
            O => \N__23275\,
            I => \N__23269\
        );

    \I__3194\ : InMux
    port map (
            O => \N__23274\,
            I => \N__23266\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__23269\,
            I => \N__23263\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__23266\,
            I => \current_shift_inst.timer_phase.counterZ0Z_3\
        );

    \I__3191\ : Odrv4
    port map (
            O => \N__23263\,
            I => \current_shift_inst.timer_phase.counterZ0Z_3\
        );

    \I__3190\ : InMux
    port map (
            O => \N__23258\,
            I => \current_shift_inst.timer_phase.counter_cry_2\
        );

    \I__3189\ : CascadeMux
    port map (
            O => \N__23255\,
            I => \N__23251\
        );

    \I__3188\ : CascadeMux
    port map (
            O => \N__23254\,
            I => \N__23248\
        );

    \I__3187\ : InMux
    port map (
            O => \N__23251\,
            I => \N__23243\
        );

    \I__3186\ : InMux
    port map (
            O => \N__23248\,
            I => \N__23243\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__23243\,
            I => \N__23239\
        );

    \I__3184\ : InMux
    port map (
            O => \N__23242\,
            I => \N__23236\
        );

    \I__3183\ : Span4Mux_h
    port map (
            O => \N__23239\,
            I => \N__23233\
        );

    \I__3182\ : LocalMux
    port map (
            O => \N__23236\,
            I => \current_shift_inst.timer_phase.counterZ0Z_4\
        );

    \I__3181\ : Odrv4
    port map (
            O => \N__23233\,
            I => \current_shift_inst.timer_phase.counterZ0Z_4\
        );

    \I__3180\ : InMux
    port map (
            O => \N__23228\,
            I => \current_shift_inst.timer_phase.counter_cry_3\
        );

    \I__3179\ : InMux
    port map (
            O => \N__23225\,
            I => \N__23219\
        );

    \I__3178\ : InMux
    port map (
            O => \N__23224\,
            I => \N__23219\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__23219\,
            I => \N__23215\
        );

    \I__3176\ : InMux
    port map (
            O => \N__23218\,
            I => \N__23212\
        );

    \I__3175\ : Span4Mux_h
    port map (
            O => \N__23215\,
            I => \N__23209\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__23212\,
            I => \current_shift_inst.timer_phase.counterZ0Z_5\
        );

    \I__3173\ : Odrv4
    port map (
            O => \N__23209\,
            I => \current_shift_inst.timer_phase.counterZ0Z_5\
        );

    \I__3172\ : InMux
    port map (
            O => \N__23204\,
            I => \current_shift_inst.timer_phase.counter_cry_4\
        );

    \I__3171\ : InMux
    port map (
            O => \N__23201\,
            I => \N__23195\
        );

    \I__3170\ : InMux
    port map (
            O => \N__23200\,
            I => \N__23195\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__23195\,
            I => \N__23191\
        );

    \I__3168\ : InMux
    port map (
            O => \N__23194\,
            I => \N__23188\
        );

    \I__3167\ : Span4Mux_h
    port map (
            O => \N__23191\,
            I => \N__23185\
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__23188\,
            I => \current_shift_inst.timer_phase.counterZ0Z_6\
        );

    \I__3165\ : Odrv4
    port map (
            O => \N__23185\,
            I => \current_shift_inst.timer_phase.counterZ0Z_6\
        );

    \I__3164\ : InMux
    port map (
            O => \N__23180\,
            I => \current_shift_inst.timer_phase.counter_cry_5\
        );

    \I__3163\ : CascadeMux
    port map (
            O => \N__23177\,
            I => \N__23173\
        );

    \I__3162\ : InMux
    port map (
            O => \N__23176\,
            I => \N__23170\
        );

    \I__3161\ : InMux
    port map (
            O => \N__23173\,
            I => \N__23167\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__23170\,
            I => \N__23162\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__23167\,
            I => \N__23162\
        );

    \I__3158\ : Span4Mux_h
    port map (
            O => \N__23162\,
            I => \N__23158\
        );

    \I__3157\ : InMux
    port map (
            O => \N__23161\,
            I => \N__23155\
        );

    \I__3156\ : Span4Mux_h
    port map (
            O => \N__23158\,
            I => \N__23152\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__23155\,
            I => \current_shift_inst.timer_phase.counterZ0Z_7\
        );

    \I__3154\ : Odrv4
    port map (
            O => \N__23152\,
            I => \current_shift_inst.timer_phase.counterZ0Z_7\
        );

    \I__3153\ : InMux
    port map (
            O => \N__23147\,
            I => \current_shift_inst.timer_phase.counter_cry_6\
        );

    \I__3152\ : InMux
    port map (
            O => \N__23144\,
            I => \current_shift_inst.z_5_cry_22\
        );

    \I__3151\ : InMux
    port map (
            O => \N__23141\,
            I => \current_shift_inst.z_5_cry_23\
        );

    \I__3150\ : InMux
    port map (
            O => \N__23138\,
            I => \bfn_8_20_0_\
        );

    \I__3149\ : InMux
    port map (
            O => \N__23135\,
            I => \current_shift_inst.z_5_cry_25\
        );

    \I__3148\ : InMux
    port map (
            O => \N__23132\,
            I => \current_shift_inst.z_5_cry_26\
        );

    \I__3147\ : InMux
    port map (
            O => \N__23129\,
            I => \current_shift_inst.z_5_cry_27\
        );

    \I__3146\ : CascadeMux
    port map (
            O => \N__23126\,
            I => \N__23123\
        );

    \I__3145\ : InMux
    port map (
            O => \N__23123\,
            I => \N__23116\
        );

    \I__3144\ : InMux
    port map (
            O => \N__23122\,
            I => \N__23116\
        );

    \I__3143\ : InMux
    port map (
            O => \N__23121\,
            I => \N__23113\
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__23116\,
            I => \N__23110\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__23113\,
            I => \N__23107\
        );

    \I__3140\ : Odrv12
    port map (
            O => \N__23110\,
            I => \current_shift_inst.elapsed_time_ns_phase_29\
        );

    \I__3139\ : Odrv4
    port map (
            O => \N__23107\,
            I => \current_shift_inst.elapsed_time_ns_phase_29\
        );

    \I__3138\ : InMux
    port map (
            O => \N__23102\,
            I => \current_shift_inst.z_5_cry_28\
        );

    \I__3137\ : InMux
    port map (
            O => \N__23099\,
            I => \N__23096\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__23096\,
            I => \N__23081\
        );

    \I__3135\ : InMux
    port map (
            O => \N__23095\,
            I => \N__23074\
        );

    \I__3134\ : InMux
    port map (
            O => \N__23094\,
            I => \N__23074\
        );

    \I__3133\ : InMux
    port map (
            O => \N__23093\,
            I => \N__23074\
        );

    \I__3132\ : InMux
    port map (
            O => \N__23092\,
            I => \N__23065\
        );

    \I__3131\ : InMux
    port map (
            O => \N__23091\,
            I => \N__23065\
        );

    \I__3130\ : InMux
    port map (
            O => \N__23090\,
            I => \N__23065\
        );

    \I__3129\ : InMux
    port map (
            O => \N__23089\,
            I => \N__23065\
        );

    \I__3128\ : CascadeMux
    port map (
            O => \N__23088\,
            I => \N__23052\
        );

    \I__3127\ : CascadeMux
    port map (
            O => \N__23087\,
            I => \N__23047\
        );

    \I__3126\ : CascadeMux
    port map (
            O => \N__23086\,
            I => \N__23044\
        );

    \I__3125\ : CascadeMux
    port map (
            O => \N__23085\,
            I => \N__23040\
        );

    \I__3124\ : CascadeMux
    port map (
            O => \N__23084\,
            I => \N__23037\
        );

    \I__3123\ : Span4Mux_v
    port map (
            O => \N__23081\,
            I => \N__23020\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__23074\,
            I => \N__23020\
        );

    \I__3121\ : LocalMux
    port map (
            O => \N__23065\,
            I => \N__23020\
        );

    \I__3120\ : InMux
    port map (
            O => \N__23064\,
            I => \N__23017\
        );

    \I__3119\ : InMux
    port map (
            O => \N__23063\,
            I => \N__23010\
        );

    \I__3118\ : InMux
    port map (
            O => \N__23062\,
            I => \N__23010\
        );

    \I__3117\ : InMux
    port map (
            O => \N__23061\,
            I => \N__23010\
        );

    \I__3116\ : InMux
    port map (
            O => \N__23060\,
            I => \N__23001\
        );

    \I__3115\ : InMux
    port map (
            O => \N__23059\,
            I => \N__23001\
        );

    \I__3114\ : InMux
    port map (
            O => \N__23058\,
            I => \N__23001\
        );

    \I__3113\ : InMux
    port map (
            O => \N__23057\,
            I => \N__23001\
        );

    \I__3112\ : CascadeMux
    port map (
            O => \N__23056\,
            I => \N__22998\
        );

    \I__3111\ : CascadeMux
    port map (
            O => \N__23055\,
            I => \N__22995\
        );

    \I__3110\ : InMux
    port map (
            O => \N__23052\,
            I => \N__22982\
        );

    \I__3109\ : InMux
    port map (
            O => \N__23051\,
            I => \N__22982\
        );

    \I__3108\ : InMux
    port map (
            O => \N__23050\,
            I => \N__22982\
        );

    \I__3107\ : InMux
    port map (
            O => \N__23047\,
            I => \N__22982\
        );

    \I__3106\ : InMux
    port map (
            O => \N__23044\,
            I => \N__22982\
        );

    \I__3105\ : InMux
    port map (
            O => \N__23043\,
            I => \N__22975\
        );

    \I__3104\ : InMux
    port map (
            O => \N__23040\,
            I => \N__22975\
        );

    \I__3103\ : InMux
    port map (
            O => \N__23037\,
            I => \N__22975\
        );

    \I__3102\ : CascadeMux
    port map (
            O => \N__23036\,
            I => \N__22971\
        );

    \I__3101\ : CascadeMux
    port map (
            O => \N__23035\,
            I => \N__22968\
        );

    \I__3100\ : CascadeMux
    port map (
            O => \N__23034\,
            I => \N__22964\
        );

    \I__3099\ : CascadeMux
    port map (
            O => \N__23033\,
            I => \N__22961\
        );

    \I__3098\ : CascadeMux
    port map (
            O => \N__23032\,
            I => \N__22958\
        );

    \I__3097\ : CascadeMux
    port map (
            O => \N__23031\,
            I => \N__22954\
        );

    \I__3096\ : CascadeMux
    port map (
            O => \N__23030\,
            I => \N__22951\
        );

    \I__3095\ : CascadeMux
    port map (
            O => \N__23029\,
            I => \N__22946\
        );

    \I__3094\ : CascadeMux
    port map (
            O => \N__23028\,
            I => \N__22943\
        );

    \I__3093\ : CascadeMux
    port map (
            O => \N__23027\,
            I => \N__22940\
        );

    \I__3092\ : Span4Mux_s1_h
    port map (
            O => \N__23020\,
            I => \N__22937\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__23017\,
            I => \N__22932\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__23010\,
            I => \N__22932\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__23001\,
            I => \N__22929\
        );

    \I__3088\ : InMux
    port map (
            O => \N__22998\,
            I => \N__22926\
        );

    \I__3087\ : InMux
    port map (
            O => \N__22995\,
            I => \N__22921\
        );

    \I__3086\ : InMux
    port map (
            O => \N__22994\,
            I => \N__22921\
        );

    \I__3085\ : InMux
    port map (
            O => \N__22993\,
            I => \N__22918\
        );

    \I__3084\ : LocalMux
    port map (
            O => \N__22982\,
            I => \N__22913\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__22975\,
            I => \N__22913\
        );

    \I__3082\ : InMux
    port map (
            O => \N__22974\,
            I => \N__22906\
        );

    \I__3081\ : InMux
    port map (
            O => \N__22971\,
            I => \N__22906\
        );

    \I__3080\ : InMux
    port map (
            O => \N__22968\,
            I => \N__22906\
        );

    \I__3079\ : InMux
    port map (
            O => \N__22967\,
            I => \N__22897\
        );

    \I__3078\ : InMux
    port map (
            O => \N__22964\,
            I => \N__22897\
        );

    \I__3077\ : InMux
    port map (
            O => \N__22961\,
            I => \N__22897\
        );

    \I__3076\ : InMux
    port map (
            O => \N__22958\,
            I => \N__22897\
        );

    \I__3075\ : InMux
    port map (
            O => \N__22957\,
            I => \N__22890\
        );

    \I__3074\ : InMux
    port map (
            O => \N__22954\,
            I => \N__22890\
        );

    \I__3073\ : InMux
    port map (
            O => \N__22951\,
            I => \N__22890\
        );

    \I__3072\ : InMux
    port map (
            O => \N__22950\,
            I => \N__22879\
        );

    \I__3071\ : InMux
    port map (
            O => \N__22949\,
            I => \N__22879\
        );

    \I__3070\ : InMux
    port map (
            O => \N__22946\,
            I => \N__22879\
        );

    \I__3069\ : InMux
    port map (
            O => \N__22943\,
            I => \N__22879\
        );

    \I__3068\ : InMux
    port map (
            O => \N__22940\,
            I => \N__22879\
        );

    \I__3067\ : Span4Mux_v
    port map (
            O => \N__22937\,
            I => \N__22863\
        );

    \I__3066\ : Span4Mux_v
    port map (
            O => \N__22932\,
            I => \N__22863\
        );

    \I__3065\ : Span4Mux_v
    port map (
            O => \N__22929\,
            I => \N__22863\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__22926\,
            I => \N__22863\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__22921\,
            I => \N__22863\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__22918\,
            I => \N__22860\
        );

    \I__3061\ : Span4Mux_v
    port map (
            O => \N__22913\,
            I => \N__22854\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__22906\,
            I => \N__22845\
        );

    \I__3059\ : LocalMux
    port map (
            O => \N__22897\,
            I => \N__22845\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__22890\,
            I => \N__22845\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__22879\,
            I => \N__22845\
        );

    \I__3056\ : CascadeMux
    port map (
            O => \N__22878\,
            I => \N__22842\
        );

    \I__3055\ : CascadeMux
    port map (
            O => \N__22877\,
            I => \N__22839\
        );

    \I__3054\ : CascadeMux
    port map (
            O => \N__22876\,
            I => \N__22835\
        );

    \I__3053\ : CascadeMux
    port map (
            O => \N__22875\,
            I => \N__22832\
        );

    \I__3052\ : CascadeMux
    port map (
            O => \N__22874\,
            I => \N__22829\
        );

    \I__3051\ : Span4Mux_h
    port map (
            O => \N__22863\,
            I => \N__22826\
        );

    \I__3050\ : IoSpan4Mux
    port map (
            O => \N__22860\,
            I => \N__22823\
        );

    \I__3049\ : InMux
    port map (
            O => \N__22859\,
            I => \N__22820\
        );

    \I__3048\ : InMux
    port map (
            O => \N__22858\,
            I => \N__22817\
        );

    \I__3047\ : InMux
    port map (
            O => \N__22857\,
            I => \N__22814\
        );

    \I__3046\ : Span4Mux_h
    port map (
            O => \N__22854\,
            I => \N__22809\
        );

    \I__3045\ : Span4Mux_v
    port map (
            O => \N__22845\,
            I => \N__22809\
        );

    \I__3044\ : InMux
    port map (
            O => \N__22842\,
            I => \N__22804\
        );

    \I__3043\ : InMux
    port map (
            O => \N__22839\,
            I => \N__22804\
        );

    \I__3042\ : InMux
    port map (
            O => \N__22838\,
            I => \N__22795\
        );

    \I__3041\ : InMux
    port map (
            O => \N__22835\,
            I => \N__22795\
        );

    \I__3040\ : InMux
    port map (
            O => \N__22832\,
            I => \N__22795\
        );

    \I__3039\ : InMux
    port map (
            O => \N__22829\,
            I => \N__22795\
        );

    \I__3038\ : Span4Mux_v
    port map (
            O => \N__22826\,
            I => \N__22792\
        );

    \I__3037\ : Span4Mux_s2_v
    port map (
            O => \N__22823\,
            I => \N__22789\
        );

    \I__3036\ : LocalMux
    port map (
            O => \N__22820\,
            I => \N__22786\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__22817\,
            I => \N__22781\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__22814\,
            I => \N__22781\
        );

    \I__3033\ : Sp12to4
    port map (
            O => \N__22809\,
            I => \N__22774\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__22804\,
            I => \N__22774\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__22795\,
            I => \N__22774\
        );

    \I__3030\ : Sp12to4
    port map (
            O => \N__22792\,
            I => \N__22771\
        );

    \I__3029\ : Span4Mux_h
    port map (
            O => \N__22789\,
            I => \N__22768\
        );

    \I__3028\ : Span4Mux_s2_v
    port map (
            O => \N__22786\,
            I => \N__22765\
        );

    \I__3027\ : Span4Mux_s2_v
    port map (
            O => \N__22781\,
            I => \N__22762\
        );

    \I__3026\ : Span12Mux_h
    port map (
            O => \N__22774\,
            I => \N__22759\
        );

    \I__3025\ : Span12Mux_v
    port map (
            O => \N__22771\,
            I => \N__22754\
        );

    \I__3024\ : Sp12to4
    port map (
            O => \N__22768\,
            I => \N__22754\
        );

    \I__3023\ : Span4Mux_h
    port map (
            O => \N__22765\,
            I => \N__22749\
        );

    \I__3022\ : Span4Mux_h
    port map (
            O => \N__22762\,
            I => \N__22749\
        );

    \I__3021\ : Odrv12
    port map (
            O => \N__22759\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3020\ : Odrv12
    port map (
            O => \N__22754\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3019\ : Odrv4
    port map (
            O => \N__22749\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3018\ : CascadeMux
    port map (
            O => \N__22742\,
            I => \N__22737\
        );

    \I__3017\ : InMux
    port map (
            O => \N__22741\,
            I => \N__22734\
        );

    \I__3016\ : InMux
    port map (
            O => \N__22740\,
            I => \N__22731\
        );

    \I__3015\ : InMux
    port map (
            O => \N__22737\,
            I => \N__22728\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__22734\,
            I => \N__22723\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__22731\,
            I => \N__22723\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__22728\,
            I => \N__22720\
        );

    \I__3011\ : Odrv12
    port map (
            O => \N__22723\,
            I => \current_shift_inst.elapsed_time_ns_phase_30\
        );

    \I__3010\ : Odrv4
    port map (
            O => \N__22720\,
            I => \current_shift_inst.elapsed_time_ns_phase_30\
        );

    \I__3009\ : InMux
    port map (
            O => \N__22715\,
            I => \current_shift_inst.z_5_cry_29\
        );

    \I__3008\ : InMux
    port map (
            O => \N__22712\,
            I => \current_shift_inst.z_5_cry_30\
        );

    \I__3007\ : InMux
    port map (
            O => \N__22709\,
            I => \current_shift_inst.z_5_cry_13\
        );

    \I__3006\ : InMux
    port map (
            O => \N__22706\,
            I => \current_shift_inst.z_5_cry_14\
        );

    \I__3005\ : InMux
    port map (
            O => \N__22703\,
            I => \current_shift_inst.z_5_cry_15\
        );

    \I__3004\ : InMux
    port map (
            O => \N__22700\,
            I => \bfn_8_19_0_\
        );

    \I__3003\ : InMux
    port map (
            O => \N__22697\,
            I => \current_shift_inst.z_5_cry_17\
        );

    \I__3002\ : InMux
    port map (
            O => \N__22694\,
            I => \current_shift_inst.z_5_cry_18\
        );

    \I__3001\ : InMux
    port map (
            O => \N__22691\,
            I => \current_shift_inst.z_5_cry_19\
        );

    \I__3000\ : InMux
    port map (
            O => \N__22688\,
            I => \current_shift_inst.z_5_cry_20\
        );

    \I__2999\ : InMux
    port map (
            O => \N__22685\,
            I => \current_shift_inst.z_5_cry_21\
        );

    \I__2998\ : InMux
    port map (
            O => \N__22682\,
            I => \current_shift_inst.z_5_cry_4\
        );

    \I__2997\ : InMux
    port map (
            O => \N__22679\,
            I => \current_shift_inst.z_5_cry_5\
        );

    \I__2996\ : InMux
    port map (
            O => \N__22676\,
            I => \current_shift_inst.z_5_cry_6\
        );

    \I__2995\ : InMux
    port map (
            O => \N__22673\,
            I => \current_shift_inst.z_5_cry_7\
        );

    \I__2994\ : InMux
    port map (
            O => \N__22670\,
            I => \bfn_8_18_0_\
        );

    \I__2993\ : InMux
    port map (
            O => \N__22667\,
            I => \current_shift_inst.z_5_cry_9\
        );

    \I__2992\ : InMux
    port map (
            O => \N__22664\,
            I => \current_shift_inst.z_5_cry_10\
        );

    \I__2991\ : InMux
    port map (
            O => \N__22661\,
            I => \current_shift_inst.z_5_cry_11\
        );

    \I__2990\ : InMux
    port map (
            O => \N__22658\,
            I => \current_shift_inst.z_5_cry_12\
        );

    \I__2989\ : InMux
    port map (
            O => \N__22655\,
            I => \current_shift_inst.control_input_1_cry_20\
        );

    \I__2988\ : InMux
    port map (
            O => \N__22652\,
            I => \current_shift_inst.control_input_1_cry_21\
        );

    \I__2987\ : InMux
    port map (
            O => \N__22649\,
            I => \current_shift_inst.control_input_1_cry_22\
        );

    \I__2986\ : InMux
    port map (
            O => \N__22646\,
            I => \bfn_8_16_0_\
        );

    \I__2985\ : InMux
    port map (
            O => \N__22643\,
            I => \current_shift_inst.control_input_1_cry_24\
        );

    \I__2984\ : CascadeMux
    port map (
            O => \N__22640\,
            I => \N__22636\
        );

    \I__2983\ : InMux
    port map (
            O => \N__22639\,
            I => \N__22631\
        );

    \I__2982\ : InMux
    port map (
            O => \N__22636\,
            I => \N__22626\
        );

    \I__2981\ : InMux
    port map (
            O => \N__22635\,
            I => \N__22626\
        );

    \I__2980\ : InMux
    port map (
            O => \N__22634\,
            I => \N__22623\
        );

    \I__2979\ : LocalMux
    port map (
            O => \N__22631\,
            I => \current_shift_inst.elapsed_time_ns_phase_2\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__22626\,
            I => \current_shift_inst.elapsed_time_ns_phase_2\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__22623\,
            I => \current_shift_inst.elapsed_time_ns_phase_2\
        );

    \I__2976\ : InMux
    port map (
            O => \N__22616\,
            I => \current_shift_inst.z_5_cry_1\
        );

    \I__2975\ : InMux
    port map (
            O => \N__22613\,
            I => \N__22608\
        );

    \I__2974\ : InMux
    port map (
            O => \N__22612\,
            I => \N__22603\
        );

    \I__2973\ : InMux
    port map (
            O => \N__22611\,
            I => \N__22603\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__22608\,
            I => \N__22600\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__22603\,
            I => \current_shift_inst.elapsed_time_ns_phase_3\
        );

    \I__2970\ : Odrv4
    port map (
            O => \N__22600\,
            I => \current_shift_inst.elapsed_time_ns_phase_3\
        );

    \I__2969\ : InMux
    port map (
            O => \N__22595\,
            I => \current_shift_inst.z_5_cry_2\
        );

    \I__2968\ : InMux
    port map (
            O => \N__22592\,
            I => \current_shift_inst.z_5_cry_3\
        );

    \I__2967\ : InMux
    port map (
            O => \N__22589\,
            I => \current_shift_inst.control_input_1_cry_11\
        );

    \I__2966\ : InMux
    port map (
            O => \N__22586\,
            I => \current_shift_inst.control_input_1_cry_12\
        );

    \I__2965\ : InMux
    port map (
            O => \N__22583\,
            I => \current_shift_inst.control_input_1_cry_13\
        );

    \I__2964\ : InMux
    port map (
            O => \N__22580\,
            I => \current_shift_inst.control_input_1_cry_14\
        );

    \I__2963\ : InMux
    port map (
            O => \N__22577\,
            I => \bfn_8_15_0_\
        );

    \I__2962\ : InMux
    port map (
            O => \N__22574\,
            I => \current_shift_inst.control_input_1_cry_16\
        );

    \I__2961\ : InMux
    port map (
            O => \N__22571\,
            I => \current_shift_inst.control_input_1_cry_17\
        );

    \I__2960\ : InMux
    port map (
            O => \N__22568\,
            I => \current_shift_inst.control_input_1_cry_18\
        );

    \I__2959\ : InMux
    port map (
            O => \N__22565\,
            I => \current_shift_inst.control_input_1_cry_19\
        );

    \I__2958\ : InMux
    port map (
            O => \N__22562\,
            I => \current_shift_inst.control_input_1_cry_2\
        );

    \I__2957\ : InMux
    port map (
            O => \N__22559\,
            I => \current_shift_inst.control_input_1_cry_3\
        );

    \I__2956\ : InMux
    port map (
            O => \N__22556\,
            I => \current_shift_inst.control_input_1_cry_4\
        );

    \I__2955\ : InMux
    port map (
            O => \N__22553\,
            I => \current_shift_inst.control_input_1_cry_5\
        );

    \I__2954\ : InMux
    port map (
            O => \N__22550\,
            I => \current_shift_inst.control_input_1_cry_6\
        );

    \I__2953\ : InMux
    port map (
            O => \N__22547\,
            I => \bfn_8_14_0_\
        );

    \I__2952\ : InMux
    port map (
            O => \N__22544\,
            I => \current_shift_inst.control_input_1_cry_8\
        );

    \I__2951\ : InMux
    port map (
            O => \N__22541\,
            I => \current_shift_inst.control_input_1_cry_9\
        );

    \I__2950\ : InMux
    port map (
            O => \N__22538\,
            I => \current_shift_inst.control_input_1_cry_10\
        );

    \I__2949\ : InMux
    port map (
            O => \N__22535\,
            I => \N__22532\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__22532\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_15\
        );

    \I__2947\ : InMux
    port map (
            O => \N__22529\,
            I => \N__22526\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__22526\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_14\
        );

    \I__2945\ : CascadeMux
    port map (
            O => \N__22523\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_12_cascade_\
        );

    \I__2944\ : InMux
    port map (
            O => \N__22520\,
            I => \N__22517\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__22517\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\
        );

    \I__2942\ : CascadeMux
    port map (
            O => \N__22514\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\
        );

    \I__2941\ : InMux
    port map (
            O => \N__22511\,
            I => \N__22508\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__22508\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0\
        );

    \I__2939\ : InMux
    port map (
            O => \N__22505\,
            I => \N__22502\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__22502\,
            I => \current_shift_inst.PI_CTRL.un1_enablelt3_0\
        );

    \I__2937\ : CascadeMux
    port map (
            O => \N__22499\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_3_cascade_\
        );

    \I__2936\ : InMux
    port map (
            O => \N__22496\,
            I => \N__22493\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__22493\,
            I => \N__22490\
        );

    \I__2934\ : Odrv4
    port map (
            O => \N__22490\,
            I => \delay_measurement_inst.delay_hc_reg3lto31_5_0\
        );

    \I__2933\ : InMux
    port map (
            O => \N__22487\,
            I => \current_shift_inst.control_input_1_cry_0\
        );

    \I__2932\ : InMux
    port map (
            O => \N__22484\,
            I => \current_shift_inst.control_input_1_cry_1\
        );

    \I__2931\ : InMux
    port map (
            O => \N__22481\,
            I => \N__22478\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__22478\,
            I => \pwm_generator_inst.thresholdZ0Z_6\
        );

    \I__2929\ : CascadeMux
    port map (
            O => \N__22475\,
            I => \N__22472\
        );

    \I__2928\ : InMux
    port map (
            O => \N__22472\,
            I => \N__22469\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__22469\,
            I => \pwm_generator_inst.counter_i_6\
        );

    \I__2926\ : CascadeMux
    port map (
            O => \N__22466\,
            I => \N__22463\
        );

    \I__2925\ : InMux
    port map (
            O => \N__22463\,
            I => \N__22460\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__22460\,
            I => \pwm_generator_inst.thresholdZ0Z_7\
        );

    \I__2923\ : InMux
    port map (
            O => \N__22457\,
            I => \N__22454\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__22454\,
            I => \pwm_generator_inst.counter_i_7\
        );

    \I__2921\ : CascadeMux
    port map (
            O => \N__22451\,
            I => \N__22448\
        );

    \I__2920\ : InMux
    port map (
            O => \N__22448\,
            I => \N__22445\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__22445\,
            I => \pwm_generator_inst.thresholdZ0Z_8\
        );

    \I__2918\ : InMux
    port map (
            O => \N__22442\,
            I => \N__22439\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__22439\,
            I => \pwm_generator_inst.counter_i_8\
        );

    \I__2916\ : CascadeMux
    port map (
            O => \N__22436\,
            I => \N__22433\
        );

    \I__2915\ : InMux
    port map (
            O => \N__22433\,
            I => \N__22430\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__22430\,
            I => \pwm_generator_inst.thresholdZ0Z_9\
        );

    \I__2913\ : InMux
    port map (
            O => \N__22427\,
            I => \N__22424\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__22424\,
            I => \pwm_generator_inst.counter_i_9\
        );

    \I__2911\ : InMux
    port map (
            O => \N__22421\,
            I => \pwm_generator_inst.un14_counter_cry_9\
        );

    \I__2910\ : IoInMux
    port map (
            O => \N__22418\,
            I => \N__22415\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__22415\,
            I => \N__22412\
        );

    \I__2908\ : IoSpan4Mux
    port map (
            O => \N__22412\,
            I => \N__22409\
        );

    \I__2907\ : Span4Mux_s2_v
    port map (
            O => \N__22409\,
            I => \N__22406\
        );

    \I__2906\ : Span4Mux_v
    port map (
            O => \N__22406\,
            I => \N__22403\
        );

    \I__2905\ : Sp12to4
    port map (
            O => \N__22403\,
            I => \N__22400\
        );

    \I__2904\ : Span12Mux_h
    port map (
            O => \N__22400\,
            I => \N__22397\
        );

    \I__2903\ : Odrv12
    port map (
            O => \N__22397\,
            I => pwm_output_c
        );

    \I__2902\ : InMux
    port map (
            O => \N__22394\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_28\
        );

    \I__2901\ : InMux
    port map (
            O => \N__22391\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_29\
        );

    \I__2900\ : CEMux
    port map (
            O => \N__22388\,
            I => \N__22373\
        );

    \I__2899\ : CEMux
    port map (
            O => \N__22387\,
            I => \N__22373\
        );

    \I__2898\ : CEMux
    port map (
            O => \N__22386\,
            I => \N__22373\
        );

    \I__2897\ : CEMux
    port map (
            O => \N__22385\,
            I => \N__22373\
        );

    \I__2896\ : CEMux
    port map (
            O => \N__22384\,
            I => \N__22373\
        );

    \I__2895\ : GlobalMux
    port map (
            O => \N__22373\,
            I => \N__22370\
        );

    \I__2894\ : gio2CtrlBuf
    port map (
            O => \N__22370\,
            I => \current_shift_inst.timer_phase.N_188_i_g\
        );

    \I__2893\ : InMux
    port map (
            O => \N__22367\,
            I => \N__22364\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__22364\,
            I => \pwm_generator_inst.thresholdZ0Z_0\
        );

    \I__2891\ : CascadeMux
    port map (
            O => \N__22361\,
            I => \N__22358\
        );

    \I__2890\ : InMux
    port map (
            O => \N__22358\,
            I => \N__22355\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__22355\,
            I => \pwm_generator_inst.counter_i_0\
        );

    \I__2888\ : InMux
    port map (
            O => \N__22352\,
            I => \N__22349\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__22349\,
            I => \pwm_generator_inst.thresholdZ0Z_1\
        );

    \I__2886\ : CascadeMux
    port map (
            O => \N__22346\,
            I => \N__22343\
        );

    \I__2885\ : InMux
    port map (
            O => \N__22343\,
            I => \N__22340\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__22340\,
            I => \pwm_generator_inst.counter_i_1\
        );

    \I__2883\ : CascadeMux
    port map (
            O => \N__22337\,
            I => \N__22334\
        );

    \I__2882\ : InMux
    port map (
            O => \N__22334\,
            I => \N__22331\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__22331\,
            I => \pwm_generator_inst.thresholdZ0Z_2\
        );

    \I__2880\ : InMux
    port map (
            O => \N__22328\,
            I => \N__22325\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__22325\,
            I => \pwm_generator_inst.counter_i_2\
        );

    \I__2878\ : CascadeMux
    port map (
            O => \N__22322\,
            I => \N__22319\
        );

    \I__2877\ : InMux
    port map (
            O => \N__22319\,
            I => \N__22316\
        );

    \I__2876\ : LocalMux
    port map (
            O => \N__22316\,
            I => \N__22313\
        );

    \I__2875\ : Span4Mux_v
    port map (
            O => \N__22313\,
            I => \N__22310\
        );

    \I__2874\ : Odrv4
    port map (
            O => \N__22310\,
            I => \pwm_generator_inst.thresholdZ0Z_3\
        );

    \I__2873\ : InMux
    port map (
            O => \N__22307\,
            I => \N__22304\
        );

    \I__2872\ : LocalMux
    port map (
            O => \N__22304\,
            I => \pwm_generator_inst.counter_i_3\
        );

    \I__2871\ : InMux
    port map (
            O => \N__22301\,
            I => \N__22298\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__22298\,
            I => \pwm_generator_inst.thresholdZ0Z_4\
        );

    \I__2869\ : CascadeMux
    port map (
            O => \N__22295\,
            I => \N__22292\
        );

    \I__2868\ : InMux
    port map (
            O => \N__22292\,
            I => \N__22289\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__22289\,
            I => \pwm_generator_inst.counter_i_4\
        );

    \I__2866\ : InMux
    port map (
            O => \N__22286\,
            I => \N__22283\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__22283\,
            I => \pwm_generator_inst.thresholdZ0Z_5\
        );

    \I__2864\ : CascadeMux
    port map (
            O => \N__22280\,
            I => \N__22277\
        );

    \I__2863\ : InMux
    port map (
            O => \N__22277\,
            I => \N__22274\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__22274\,
            I => \pwm_generator_inst.counter_i_5\
        );

    \I__2861\ : InMux
    port map (
            O => \N__22271\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_19\
        );

    \I__2860\ : InMux
    port map (
            O => \N__22268\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_20\
        );

    \I__2859\ : InMux
    port map (
            O => \N__22265\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_21\
        );

    \I__2858\ : InMux
    port map (
            O => \N__22262\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_22\
        );

    \I__2857\ : InMux
    port map (
            O => \N__22259\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_23\
        );

    \I__2856\ : InMux
    port map (
            O => \N__22256\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_24\
        );

    \I__2855\ : InMux
    port map (
            O => \N__22253\,
            I => \bfn_7_22_0_\
        );

    \I__2854\ : InMux
    port map (
            O => \N__22250\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_26\
        );

    \I__2853\ : InMux
    port map (
            O => \N__22247\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_27\
        );

    \I__2852\ : InMux
    port map (
            O => \N__22244\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_10\
        );

    \I__2851\ : InMux
    port map (
            O => \N__22241\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_11\
        );

    \I__2850\ : InMux
    port map (
            O => \N__22238\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_12\
        );

    \I__2849\ : InMux
    port map (
            O => \N__22235\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_13\
        );

    \I__2848\ : InMux
    port map (
            O => \N__22232\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_14\
        );

    \I__2847\ : InMux
    port map (
            O => \N__22229\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_15\
        );

    \I__2846\ : InMux
    port map (
            O => \N__22226\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_16\
        );

    \I__2845\ : InMux
    port map (
            O => \N__22223\,
            I => \bfn_7_21_0_\
        );

    \I__2844\ : InMux
    port map (
            O => \N__22220\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_18\
        );

    \I__2843\ : InMux
    port map (
            O => \N__22217\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_2\
        );

    \I__2842\ : InMux
    port map (
            O => \N__22214\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_3\
        );

    \I__2841\ : InMux
    port map (
            O => \N__22211\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_4\
        );

    \I__2840\ : InMux
    port map (
            O => \N__22208\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_5\
        );

    \I__2839\ : InMux
    port map (
            O => \N__22205\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_6\
        );

    \I__2838\ : InMux
    port map (
            O => \N__22202\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_7\
        );

    \I__2837\ : InMux
    port map (
            O => \N__22199\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_8\
        );

    \I__2836\ : InMux
    port map (
            O => \N__22196\,
            I => \bfn_7_20_0_\
        );

    \I__2835\ : InMux
    port map (
            O => \N__22193\,
            I => \N__22190\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__22190\,
            I => \N__22187\
        );

    \I__2833\ : Odrv4
    port map (
            O => \N__22187\,
            I => \delay_measurement_inst.delay_hc_reg3lt19_0\
        );

    \I__2832\ : CascadeMux
    port map (
            O => \N__22184\,
            I => \delay_measurement_inst.delay_hc_reg3lt19_0_cascade_\
        );

    \I__2831\ : CascadeMux
    port map (
            O => \N__22181\,
            I => \N__22178\
        );

    \I__2830\ : InMux
    port map (
            O => \N__22178\,
            I => \N__22175\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__22175\,
            I => \N__22172\
        );

    \I__2828\ : Span4Mux_v
    port map (
            O => \N__22172\,
            I => \N__22169\
        );

    \I__2827\ : Odrv4
    port map (
            O => \N__22169\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_22\
        );

    \I__2826\ : CascadeMux
    port map (
            O => \N__22166\,
            I => \N__22163\
        );

    \I__2825\ : InMux
    port map (
            O => \N__22163\,
            I => \N__22160\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__22160\,
            I => \N__22157\
        );

    \I__2823\ : Span4Mux_v
    port map (
            O => \N__22157\,
            I => \N__22154\
        );

    \I__2822\ : Odrv4
    port map (
            O => \N__22154\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_17\
        );

    \I__2821\ : CascadeMux
    port map (
            O => \N__22151\,
            I => \N__22144\
        );

    \I__2820\ : CascadeMux
    port map (
            O => \N__22150\,
            I => \N__22140\
        );

    \I__2819\ : CascadeMux
    port map (
            O => \N__22149\,
            I => \N__22136\
        );

    \I__2818\ : InMux
    port map (
            O => \N__22148\,
            I => \N__22121\
        );

    \I__2817\ : InMux
    port map (
            O => \N__22147\,
            I => \N__22121\
        );

    \I__2816\ : InMux
    port map (
            O => \N__22144\,
            I => \N__22121\
        );

    \I__2815\ : InMux
    port map (
            O => \N__22143\,
            I => \N__22121\
        );

    \I__2814\ : InMux
    port map (
            O => \N__22140\,
            I => \N__22121\
        );

    \I__2813\ : InMux
    port map (
            O => \N__22139\,
            I => \N__22121\
        );

    \I__2812\ : InMux
    port map (
            O => \N__22136\,
            I => \N__22121\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__22121\,
            I => \N__22118\
        );

    \I__2810\ : Odrv12
    port map (
            O => \N__22118\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_25\
        );

    \I__2809\ : CascadeMux
    port map (
            O => \N__22115\,
            I => \N__22112\
        );

    \I__2808\ : InMux
    port map (
            O => \N__22112\,
            I => \N__22109\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__22109\,
            I => \N__22106\
        );

    \I__2806\ : Span4Mux_h
    port map (
            O => \N__22106\,
            I => \N__22103\
        );

    \I__2805\ : Odrv4
    port map (
            O => \N__22103\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_23\
        );

    \I__2804\ : InMux
    port map (
            O => \N__22100\,
            I => \N__22097\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__22097\,
            I => \N__22093\
        );

    \I__2802\ : CascadeMux
    port map (
            O => \N__22096\,
            I => \N__22089\
        );

    \I__2801\ : Span4Mux_h
    port map (
            O => \N__22093\,
            I => \N__22086\
        );

    \I__2800\ : CascadeMux
    port map (
            O => \N__22092\,
            I => \N__22082\
        );

    \I__2799\ : InMux
    port map (
            O => \N__22089\,
            I => \N__22079\
        );

    \I__2798\ : Span4Mux_v
    port map (
            O => \N__22086\,
            I => \N__22076\
        );

    \I__2797\ : InMux
    port map (
            O => \N__22085\,
            I => \N__22071\
        );

    \I__2796\ : InMux
    port map (
            O => \N__22082\,
            I => \N__22071\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__22079\,
            I => clk_10khz_i
        );

    \I__2794\ : Odrv4
    port map (
            O => \N__22076\,
            I => clk_10khz_i
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__22071\,
            I => clk_10khz_i
        );

    \I__2792\ : InMux
    port map (
            O => \N__22064\,
            I => \N__22061\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__22061\,
            I => \N__22058\
        );

    \I__2790\ : Span4Mux_h
    port map (
            O => \N__22058\,
            I => \N__22055\
        );

    \I__2789\ : Span4Mux_v
    port map (
            O => \N__22055\,
            I => \N__22052\
        );

    \I__2788\ : Odrv4
    port map (
            O => \N__22052\,
            I => \clk_10khz_RNIIENAZ0Z2\
        );

    \I__2787\ : InMux
    port map (
            O => \N__22049\,
            I => \N__22046\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__22046\,
            I => \N__22043\
        );

    \I__2785\ : Odrv4
    port map (
            O => \N__22043\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_1\
        );

    \I__2784\ : InMux
    port map (
            O => \N__22040\,
            I => \N__22037\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__22037\,
            I => \N__22034\
        );

    \I__2782\ : Odrv4
    port map (
            O => \N__22034\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_4\
        );

    \I__2781\ : InMux
    port map (
            O => \N__22031\,
            I => \N__22028\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__22028\,
            I => \N__22025\
        );

    \I__2779\ : Span4Mux_v
    port map (
            O => \N__22025\,
            I => \N__22022\
        );

    \I__2778\ : Span4Mux_h
    port map (
            O => \N__22022\,
            I => \N__22019\
        );

    \I__2777\ : Odrv4
    port map (
            O => \N__22019\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_9\
        );

    \I__2776\ : InMux
    port map (
            O => \N__22016\,
            I => \N__22013\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__22013\,
            I => \N__22010\
        );

    \I__2774\ : Span4Mux_v
    port map (
            O => \N__22010\,
            I => \N__22007\
        );

    \I__2773\ : Span4Mux_h
    port map (
            O => \N__22007\,
            I => \N__22004\
        );

    \I__2772\ : Odrv4
    port map (
            O => \N__22004\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_8\
        );

    \I__2771\ : InMux
    port map (
            O => \N__22001\,
            I => \N__21998\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__21998\,
            I => \N__21995\
        );

    \I__2769\ : Span4Mux_v
    port map (
            O => \N__21995\,
            I => \N__21992\
        );

    \I__2768\ : Odrv4
    port map (
            O => \N__21992\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\
        );

    \I__2767\ : CascadeMux
    port map (
            O => \N__21989\,
            I => \N__21986\
        );

    \I__2766\ : InMux
    port map (
            O => \N__21986\,
            I => \N__21983\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__21983\,
            I => \N__21980\
        );

    \I__2764\ : Odrv4
    port map (
            O => \N__21980\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\
        );

    \I__2763\ : CascadeMux
    port map (
            O => \N__21977\,
            I => \N__21974\
        );

    \I__2762\ : InMux
    port map (
            O => \N__21974\,
            I => \N__21971\
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__21971\,
            I => \N__21968\
        );

    \I__2760\ : Span4Mux_h
    port map (
            O => \N__21968\,
            I => \N__21965\
        );

    \I__2759\ : Span4Mux_h
    port map (
            O => \N__21965\,
            I => \N__21962\
        );

    \I__2758\ : Odrv4
    port map (
            O => \N__21962\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\
        );

    \I__2757\ : CascadeMux
    port map (
            O => \N__21959\,
            I => \N__21956\
        );

    \I__2756\ : InMux
    port map (
            O => \N__21956\,
            I => \N__21953\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__21953\,
            I => \N__21950\
        );

    \I__2754\ : Odrv12
    port map (
            O => \N__21950\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\
        );

    \I__2753\ : CascadeMux
    port map (
            O => \N__21947\,
            I => \N__21944\
        );

    \I__2752\ : InMux
    port map (
            O => \N__21944\,
            I => \N__21941\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__21941\,
            I => \N__21938\
        );

    \I__2750\ : Span4Mux_v
    port map (
            O => \N__21938\,
            I => \N__21935\
        );

    \I__2749\ : Odrv4
    port map (
            O => \N__21935\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\
        );

    \I__2748\ : CascadeMux
    port map (
            O => \N__21932\,
            I => \N__21928\
        );

    \I__2747\ : CascadeMux
    port map (
            O => \N__21931\,
            I => \N__21925\
        );

    \I__2746\ : InMux
    port map (
            O => \N__21928\,
            I => \N__21922\
        );

    \I__2745\ : InMux
    port map (
            O => \N__21925\,
            I => \N__21919\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__21922\,
            I => \N__21916\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__21919\,
            I => \N__21913\
        );

    \I__2742\ : Span4Mux_h
    port map (
            O => \N__21916\,
            I => \N__21910\
        );

    \I__2741\ : Span4Mux_h
    port map (
            O => \N__21913\,
            I => \N__21907\
        );

    \I__2740\ : Odrv4
    port map (
            O => \N__21910\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__2739\ : Odrv4
    port map (
            O => \N__21907\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__2738\ : InMux
    port map (
            O => \N__21902\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\
        );

    \I__2737\ : InMux
    port map (
            O => \N__21899\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\
        );

    \I__2736\ : CascadeMux
    port map (
            O => \N__21896\,
            I => \N__21887\
        );

    \I__2735\ : CascadeMux
    port map (
            O => \N__21895\,
            I => \N__21884\
        );

    \I__2734\ : CascadeMux
    port map (
            O => \N__21894\,
            I => \N__21881\
        );

    \I__2733\ : CascadeMux
    port map (
            O => \N__21893\,
            I => \N__21878\
        );

    \I__2732\ : CascadeMux
    port map (
            O => \N__21892\,
            I => \N__21875\
        );

    \I__2731\ : CascadeMux
    port map (
            O => \N__21891\,
            I => \N__21872\
        );

    \I__2730\ : CascadeMux
    port map (
            O => \N__21890\,
            I => \N__21869\
        );

    \I__2729\ : InMux
    port map (
            O => \N__21887\,
            I => \N__21866\
        );

    \I__2728\ : InMux
    port map (
            O => \N__21884\,
            I => \N__21863\
        );

    \I__2727\ : InMux
    port map (
            O => \N__21881\,
            I => \N__21855\
        );

    \I__2726\ : InMux
    port map (
            O => \N__21878\,
            I => \N__21855\
        );

    \I__2725\ : InMux
    port map (
            O => \N__21875\,
            I => \N__21850\
        );

    \I__2724\ : InMux
    port map (
            O => \N__21872\,
            I => \N__21850\
        );

    \I__2723\ : InMux
    port map (
            O => \N__21869\,
            I => \N__21847\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__21866\,
            I => \N__21844\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__21863\,
            I => \N__21841\
        );

    \I__2720\ : InMux
    port map (
            O => \N__21862\,
            I => \N__21836\
        );

    \I__2719\ : InMux
    port map (
            O => \N__21861\,
            I => \N__21836\
        );

    \I__2718\ : InMux
    port map (
            O => \N__21860\,
            I => \N__21833\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__21855\,
            I => \N__21830\
        );

    \I__2716\ : LocalMux
    port map (
            O => \N__21850\,
            I => \N__21825\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__21847\,
            I => \N__21825\
        );

    \I__2714\ : Span4Mux_v
    port map (
            O => \N__21844\,
            I => \N__21818\
        );

    \I__2713\ : Span4Mux_s2_h
    port map (
            O => \N__21841\,
            I => \N__21818\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__21836\,
            I => \N__21818\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__21833\,
            I => \N__21815\
        );

    \I__2710\ : Span4Mux_h
    port map (
            O => \N__21830\,
            I => \N__21810\
        );

    \I__2709\ : Span4Mux_h
    port map (
            O => \N__21825\,
            I => \N__21810\
        );

    \I__2708\ : Span4Mux_h
    port map (
            O => \N__21818\,
            I => \N__21807\
        );

    \I__2707\ : Span12Mux_s5_h
    port map (
            O => \N__21815\,
            I => \N__21804\
        );

    \I__2706\ : Span4Mux_v
    port map (
            O => \N__21810\,
            I => \N__21801\
        );

    \I__2705\ : Span4Mux_v
    port map (
            O => \N__21807\,
            I => \N__21798\
        );

    \I__2704\ : Odrv12
    port map (
            O => \N__21804\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__2703\ : Odrv4
    port map (
            O => \N__21801\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__2702\ : Odrv4
    port map (
            O => \N__21798\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__2701\ : CascadeMux
    port map (
            O => \N__21791\,
            I => \N__21788\
        );

    \I__2700\ : InMux
    port map (
            O => \N__21788\,
            I => \N__21785\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__21785\,
            I => \N__21782\
        );

    \I__2698\ : Odrv4
    port map (
            O => \N__21782\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_19\
        );

    \I__2697\ : InMux
    port map (
            O => \N__21779\,
            I => \N__21776\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__21776\,
            I => \N__21773\
        );

    \I__2695\ : Odrv4
    port map (
            O => \N__21773\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_6\
        );

    \I__2694\ : InMux
    port map (
            O => \N__21770\,
            I => \N__21767\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__21767\,
            I => \N__21764\
        );

    \I__2692\ : Span4Mux_v
    port map (
            O => \N__21764\,
            I => \N__21761\
        );

    \I__2691\ : Span4Mux_h
    port map (
            O => \N__21761\,
            I => \N__21758\
        );

    \I__2690\ : Odrv4
    port map (
            O => \N__21758\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_2\
        );

    \I__2689\ : InMux
    port map (
            O => \N__21755\,
            I => \N__21752\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__21752\,
            I => \N__21749\
        );

    \I__2687\ : Odrv12
    port map (
            O => \N__21749\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_0\
        );

    \I__2686\ : InMux
    port map (
            O => \N__21746\,
            I => \N__21743\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__21743\,
            I => \N__21740\
        );

    \I__2684\ : Odrv4
    port map (
            O => \N__21740\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_5\
        );

    \I__2683\ : InMux
    port map (
            O => \N__21737\,
            I => \N__21734\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__21734\,
            I => \N__21731\
        );

    \I__2681\ : Span4Mux_h
    port map (
            O => \N__21731\,
            I => \N__21728\
        );

    \I__2680\ : Odrv4
    port map (
            O => \N__21728\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_7\
        );

    \I__2679\ : InMux
    port map (
            O => \N__21725\,
            I => \N__21722\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__21722\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_21\
        );

    \I__2677\ : InMux
    port map (
            O => \N__21719\,
            I => \N__21715\
        );

    \I__2676\ : InMux
    port map (
            O => \N__21718\,
            I => \N__21712\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__21715\,
            I => \N__21709\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__21712\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__2673\ : Odrv4
    port map (
            O => \N__21709\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__2672\ : InMux
    port map (
            O => \N__21704\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\
        );

    \I__2671\ : InMux
    port map (
            O => \N__21701\,
            I => \N__21697\
        );

    \I__2670\ : InMux
    port map (
            O => \N__21700\,
            I => \N__21694\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__21697\,
            I => \N__21691\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__21694\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__2667\ : Odrv4
    port map (
            O => \N__21691\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__2666\ : InMux
    port map (
            O => \N__21686\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\
        );

    \I__2665\ : InMux
    port map (
            O => \N__21683\,
            I => \N__21677\
        );

    \I__2664\ : InMux
    port map (
            O => \N__21682\,
            I => \N__21677\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__21677\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\
        );

    \I__2662\ : InMux
    port map (
            O => \N__21674\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\
        );

    \I__2661\ : InMux
    port map (
            O => \N__21671\,
            I => \N__21668\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__21668\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_24\
        );

    \I__2659\ : InMux
    port map (
            O => \N__21665\,
            I => \N__21661\
        );

    \I__2658\ : InMux
    port map (
            O => \N__21664\,
            I => \N__21658\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__21661\,
            I => \N__21653\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__21658\,
            I => \N__21653\
        );

    \I__2655\ : Span4Mux_h
    port map (
            O => \N__21653\,
            I => \N__21650\
        );

    \I__2654\ : Odrv4
    port map (
            O => \N__21650\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\
        );

    \I__2653\ : InMux
    port map (
            O => \N__21647\,
            I => \bfn_5_12_0_\
        );

    \I__2652\ : InMux
    port map (
            O => \N__21644\,
            I => \N__21638\
        );

    \I__2651\ : InMux
    port map (
            O => \N__21643\,
            I => \N__21638\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__21638\,
            I => \N__21635\
        );

    \I__2649\ : Span4Mux_v
    port map (
            O => \N__21635\,
            I => \N__21632\
        );

    \I__2648\ : Odrv4
    port map (
            O => \N__21632\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\
        );

    \I__2647\ : InMux
    port map (
            O => \N__21629\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\
        );

    \I__2646\ : CascadeMux
    port map (
            O => \N__21626\,
            I => \N__21622\
        );

    \I__2645\ : InMux
    port map (
            O => \N__21625\,
            I => \N__21619\
        );

    \I__2644\ : InMux
    port map (
            O => \N__21622\,
            I => \N__21616\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__21619\,
            I => \N__21613\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__21616\,
            I => \N__21610\
        );

    \I__2641\ : Span4Mux_v
    port map (
            O => \N__21613\,
            I => \N__21607\
        );

    \I__2640\ : Span4Mux_v
    port map (
            O => \N__21610\,
            I => \N__21602\
        );

    \I__2639\ : Span4Mux_v
    port map (
            O => \N__21607\,
            I => \N__21602\
        );

    \I__2638\ : Odrv4
    port map (
            O => \N__21602\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\
        );

    \I__2637\ : InMux
    port map (
            O => \N__21599\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\
        );

    \I__2636\ : CascadeMux
    port map (
            O => \N__21596\,
            I => \N__21592\
        );

    \I__2635\ : InMux
    port map (
            O => \N__21595\,
            I => \N__21587\
        );

    \I__2634\ : InMux
    port map (
            O => \N__21592\,
            I => \N__21587\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__21587\,
            I => \N__21584\
        );

    \I__2632\ : Span4Mux_h
    port map (
            O => \N__21584\,
            I => \N__21581\
        );

    \I__2631\ : Odrv4
    port map (
            O => \N__21581\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__2630\ : InMux
    port map (
            O => \N__21578\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\
        );

    \I__2629\ : InMux
    port map (
            O => \N__21575\,
            I => \N__21569\
        );

    \I__2628\ : InMux
    port map (
            O => \N__21574\,
            I => \N__21569\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__21569\,
            I => \N__21566\
        );

    \I__2626\ : Span4Mux_h
    port map (
            O => \N__21566\,
            I => \N__21563\
        );

    \I__2625\ : Odrv4
    port map (
            O => \N__21563\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__2624\ : InMux
    port map (
            O => \N__21560\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\
        );

    \I__2623\ : InMux
    port map (
            O => \N__21557\,
            I => \N__21551\
        );

    \I__2622\ : InMux
    port map (
            O => \N__21556\,
            I => \N__21551\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__21551\,
            I => \N__21548\
        );

    \I__2620\ : Span4Mux_h
    port map (
            O => \N__21548\,
            I => \N__21545\
        );

    \I__2619\ : Odrv4
    port map (
            O => \N__21545\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__2618\ : InMux
    port map (
            O => \N__21542\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\
        );

    \I__2617\ : CascadeMux
    port map (
            O => \N__21539\,
            I => \N__21535\
        );

    \I__2616\ : InMux
    port map (
            O => \N__21538\,
            I => \N__21532\
        );

    \I__2615\ : InMux
    port map (
            O => \N__21535\,
            I => \N__21529\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__21532\,
            I => \N__21526\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__21529\,
            I => \N__21521\
        );

    \I__2612\ : Span4Mux_v
    port map (
            O => \N__21526\,
            I => \N__21521\
        );

    \I__2611\ : Odrv4
    port map (
            O => \N__21521\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__2610\ : InMux
    port map (
            O => \N__21518\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\
        );

    \I__2609\ : InMux
    port map (
            O => \N__21515\,
            I => \N__21509\
        );

    \I__2608\ : InMux
    port map (
            O => \N__21514\,
            I => \N__21509\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__21509\,
            I => \N__21506\
        );

    \I__2606\ : Odrv4
    port map (
            O => \N__21506\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__2605\ : InMux
    port map (
            O => \N__21503\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\
        );

    \I__2604\ : InMux
    port map (
            O => \N__21500\,
            I => \N__21497\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__21497\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_15\
        );

    \I__2602\ : InMux
    port map (
            O => \N__21494\,
            I => \N__21488\
        );

    \I__2601\ : InMux
    port map (
            O => \N__21493\,
            I => \N__21488\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__21488\,
            I => \N__21485\
        );

    \I__2599\ : Odrv4
    port map (
            O => \N__21485\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__2598\ : InMux
    port map (
            O => \N__21482\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\
        );

    \I__2597\ : InMux
    port map (
            O => \N__21479\,
            I => \N__21476\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__21476\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_16\
        );

    \I__2595\ : InMux
    port map (
            O => \N__21473\,
            I => \N__21470\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__21470\,
            I => \N__21466\
        );

    \I__2593\ : InMux
    port map (
            O => \N__21469\,
            I => \N__21463\
        );

    \I__2592\ : Span4Mux_v
    port map (
            O => \N__21466\,
            I => \N__21460\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__21463\,
            I => \N__21457\
        );

    \I__2590\ : Odrv4
    port map (
            O => \N__21460\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__2589\ : Odrv12
    port map (
            O => \N__21457\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__2588\ : InMux
    port map (
            O => \N__21452\,
            I => \bfn_5_11_0_\
        );

    \I__2587\ : CascadeMux
    port map (
            O => \N__21449\,
            I => \N__21445\
        );

    \I__2586\ : InMux
    port map (
            O => \N__21448\,
            I => \N__21440\
        );

    \I__2585\ : InMux
    port map (
            O => \N__21445\,
            I => \N__21440\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__21440\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__2583\ : InMux
    port map (
            O => \N__21437\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\
        );

    \I__2582\ : CascadeMux
    port map (
            O => \N__21434\,
            I => \N__21431\
        );

    \I__2581\ : InMux
    port map (
            O => \N__21431\,
            I => \N__21428\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__21428\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_18\
        );

    \I__2579\ : InMux
    port map (
            O => \N__21425\,
            I => \N__21421\
        );

    \I__2578\ : InMux
    port map (
            O => \N__21424\,
            I => \N__21418\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__21421\,
            I => \N__21415\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__21418\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__2575\ : Odrv12
    port map (
            O => \N__21415\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__2574\ : InMux
    port map (
            O => \N__21410\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\
        );

    \I__2573\ : InMux
    port map (
            O => \N__21407\,
            I => \N__21401\
        );

    \I__2572\ : InMux
    port map (
            O => \N__21406\,
            I => \N__21401\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__21401\,
            I => \N__21398\
        );

    \I__2570\ : Odrv4
    port map (
            O => \N__21398\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__2569\ : InMux
    port map (
            O => \N__21395\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\
        );

    \I__2568\ : CascadeMux
    port map (
            O => \N__21392\,
            I => \N__21389\
        );

    \I__2567\ : InMux
    port map (
            O => \N__21389\,
            I => \N__21386\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__21386\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_20\
        );

    \I__2565\ : InMux
    port map (
            O => \N__21383\,
            I => \N__21379\
        );

    \I__2564\ : InMux
    port map (
            O => \N__21382\,
            I => \N__21376\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__21379\,
            I => \N__21373\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__21376\,
            I => \N__21370\
        );

    \I__2561\ : Span4Mux_h
    port map (
            O => \N__21373\,
            I => \N__21367\
        );

    \I__2560\ : Odrv4
    port map (
            O => \N__21370\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__2559\ : Odrv4
    port map (
            O => \N__21367\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__2558\ : InMux
    port map (
            O => \N__21362\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\
        );

    \I__2557\ : CascadeMux
    port map (
            O => \N__21359\,
            I => \N__21356\
        );

    \I__2556\ : InMux
    port map (
            O => \N__21356\,
            I => \N__21353\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__21353\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\
        );

    \I__2554\ : InMux
    port map (
            O => \N__21350\,
            I => \N__21344\
        );

    \I__2553\ : InMux
    port map (
            O => \N__21349\,
            I => \N__21344\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__21344\,
            I => \N__21340\
        );

    \I__2551\ : InMux
    port map (
            O => \N__21343\,
            I => \N__21337\
        );

    \I__2550\ : Span4Mux_s3_h
    port map (
            O => \N__21340\,
            I => \N__21332\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__21337\,
            I => \N__21332\
        );

    \I__2548\ : Span4Mux_v
    port map (
            O => \N__21332\,
            I => \N__21329\
        );

    \I__2547\ : Odrv4
    port map (
            O => \N__21329\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__2546\ : InMux
    port map (
            O => \N__21326\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\
        );

    \I__2545\ : InMux
    port map (
            O => \N__21323\,
            I => \N__21319\
        );

    \I__2544\ : InMux
    port map (
            O => \N__21322\,
            I => \N__21316\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__21319\,
            I => \N__21310\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__21316\,
            I => \N__21310\
        );

    \I__2541\ : InMux
    port map (
            O => \N__21315\,
            I => \N__21307\
        );

    \I__2540\ : Span4Mux_v
    port map (
            O => \N__21310\,
            I => \N__21302\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__21307\,
            I => \N__21302\
        );

    \I__2538\ : Span4Mux_h
    port map (
            O => \N__21302\,
            I => \N__21299\
        );

    \I__2537\ : Odrv4
    port map (
            O => \N__21299\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__2536\ : InMux
    port map (
            O => \N__21296\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\
        );

    \I__2535\ : InMux
    port map (
            O => \N__21293\,
            I => \N__21290\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__21290\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\
        );

    \I__2533\ : InMux
    port map (
            O => \N__21287\,
            I => \N__21283\
        );

    \I__2532\ : InMux
    port map (
            O => \N__21286\,
            I => \N__21280\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__21283\,
            I => \N__21274\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__21280\,
            I => \N__21274\
        );

    \I__2529\ : InMux
    port map (
            O => \N__21279\,
            I => \N__21271\
        );

    \I__2528\ : Span4Mux_v
    port map (
            O => \N__21274\,
            I => \N__21266\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__21271\,
            I => \N__21266\
        );

    \I__2526\ : Span4Mux_h
    port map (
            O => \N__21266\,
            I => \N__21263\
        );

    \I__2525\ : Odrv4
    port map (
            O => \N__21263\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__2524\ : InMux
    port map (
            O => \N__21260\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\
        );

    \I__2523\ : CascadeMux
    port map (
            O => \N__21257\,
            I => \N__21254\
        );

    \I__2522\ : InMux
    port map (
            O => \N__21254\,
            I => \N__21251\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__21251\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\
        );

    \I__2520\ : InMux
    port map (
            O => \N__21248\,
            I => \N__21244\
        );

    \I__2519\ : InMux
    port map (
            O => \N__21247\,
            I => \N__21241\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__21244\,
            I => \N__21237\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__21241\,
            I => \N__21234\
        );

    \I__2516\ : InMux
    port map (
            O => \N__21240\,
            I => \N__21231\
        );

    \I__2515\ : Span4Mux_v
    port map (
            O => \N__21237\,
            I => \N__21228\
        );

    \I__2514\ : Span4Mux_v
    port map (
            O => \N__21234\,
            I => \N__21223\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__21231\,
            I => \N__21223\
        );

    \I__2512\ : Span4Mux_h
    port map (
            O => \N__21228\,
            I => \N__21220\
        );

    \I__2511\ : Span4Mux_h
    port map (
            O => \N__21223\,
            I => \N__21217\
        );

    \I__2510\ : Odrv4
    port map (
            O => \N__21220\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__2509\ : Odrv4
    port map (
            O => \N__21217\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__2508\ : InMux
    port map (
            O => \N__21212\,
            I => \bfn_5_10_0_\
        );

    \I__2507\ : InMux
    port map (
            O => \N__21209\,
            I => \N__21205\
        );

    \I__2506\ : InMux
    port map (
            O => \N__21208\,
            I => \N__21202\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__21205\,
            I => \N__21198\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__21202\,
            I => \N__21195\
        );

    \I__2503\ : InMux
    port map (
            O => \N__21201\,
            I => \N__21192\
        );

    \I__2502\ : Span4Mux_v
    port map (
            O => \N__21198\,
            I => \N__21189\
        );

    \I__2501\ : Span4Mux_v
    port map (
            O => \N__21195\,
            I => \N__21184\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__21192\,
            I => \N__21184\
        );

    \I__2499\ : Span4Mux_h
    port map (
            O => \N__21189\,
            I => \N__21181\
        );

    \I__2498\ : Span4Mux_h
    port map (
            O => \N__21184\,
            I => \N__21178\
        );

    \I__2497\ : Odrv4
    port map (
            O => \N__21181\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__2496\ : Odrv4
    port map (
            O => \N__21178\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__2495\ : InMux
    port map (
            O => \N__21173\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\
        );

    \I__2494\ : CascadeMux
    port map (
            O => \N__21170\,
            I => \N__21167\
        );

    \I__2493\ : InMux
    port map (
            O => \N__21167\,
            I => \N__21164\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__21164\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\
        );

    \I__2491\ : InMux
    port map (
            O => \N__21161\,
            I => \N__21155\
        );

    \I__2490\ : InMux
    port map (
            O => \N__21160\,
            I => \N__21155\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__21155\,
            I => \N__21152\
        );

    \I__2488\ : Odrv4
    port map (
            O => \N__21152\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\
        );

    \I__2487\ : InMux
    port map (
            O => \N__21149\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\
        );

    \I__2486\ : CascadeMux
    port map (
            O => \N__21146\,
            I => \N__21143\
        );

    \I__2485\ : InMux
    port map (
            O => \N__21143\,
            I => \N__21140\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__21140\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\
        );

    \I__2483\ : InMux
    port map (
            O => \N__21137\,
            I => \N__21133\
        );

    \I__2482\ : InMux
    port map (
            O => \N__21136\,
            I => \N__21130\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__21133\,
            I => \N__21127\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__21130\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\
        );

    \I__2479\ : Odrv4
    port map (
            O => \N__21127\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\
        );

    \I__2478\ : InMux
    port map (
            O => \N__21122\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\
        );

    \I__2477\ : CascadeMux
    port map (
            O => \N__21119\,
            I => \N__21116\
        );

    \I__2476\ : InMux
    port map (
            O => \N__21116\,
            I => \N__21113\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__21113\,
            I => \N__21110\
        );

    \I__2474\ : Odrv4
    port map (
            O => \N__21110\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\
        );

    \I__2473\ : InMux
    port map (
            O => \N__21107\,
            I => \N__21101\
        );

    \I__2472\ : InMux
    port map (
            O => \N__21106\,
            I => \N__21101\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__21101\,
            I => \N__21098\
        );

    \I__2470\ : Odrv4
    port map (
            O => \N__21098\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__2469\ : InMux
    port map (
            O => \N__21095\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\
        );

    \I__2468\ : CascadeMux
    port map (
            O => \N__21092\,
            I => \N__21086\
        );

    \I__2467\ : InMux
    port map (
            O => \N__21091\,
            I => \N__21077\
        );

    \I__2466\ : InMux
    port map (
            O => \N__21090\,
            I => \N__21077\
        );

    \I__2465\ : InMux
    port map (
            O => \N__21089\,
            I => \N__21077\
        );

    \I__2464\ : InMux
    port map (
            O => \N__21086\,
            I => \N__21074\
        );

    \I__2463\ : InMux
    port map (
            O => \N__21085\,
            I => \N__21071\
        );

    \I__2462\ : InMux
    port map (
            O => \N__21084\,
            I => \N__21068\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__21077\,
            I => un2_counter_8
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__21074\,
            I => un2_counter_8
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__21071\,
            I => un2_counter_8
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__21068\,
            I => un2_counter_8
        );

    \I__2457\ : InMux
    port map (
            O => \N__21059\,
            I => \N__21051\
        );

    \I__2456\ : InMux
    port map (
            O => \N__21058\,
            I => \N__21046\
        );

    \I__2455\ : InMux
    port map (
            O => \N__21057\,
            I => \N__21046\
        );

    \I__2454\ : InMux
    port map (
            O => \N__21056\,
            I => \N__21043\
        );

    \I__2453\ : InMux
    port map (
            O => \N__21055\,
            I => \N__21040\
        );

    \I__2452\ : InMux
    port map (
            O => \N__21054\,
            I => \N__21037\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__21051\,
            I => un2_counter_7
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__21046\,
            I => un2_counter_7
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__21043\,
            I => un2_counter_7
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__21040\,
            I => un2_counter_7
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__21037\,
            I => un2_counter_7
        );

    \I__2446\ : InMux
    port map (
            O => \N__21026\,
            I => \N__21018\
        );

    \I__2445\ : InMux
    port map (
            O => \N__21025\,
            I => \N__21015\
        );

    \I__2444\ : InMux
    port map (
            O => \N__21024\,
            I => \N__21012\
        );

    \I__2443\ : InMux
    port map (
            O => \N__21023\,
            I => \N__21005\
        );

    \I__2442\ : InMux
    port map (
            O => \N__21022\,
            I => \N__21005\
        );

    \I__2441\ : InMux
    port map (
            O => \N__21021\,
            I => \N__21005\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__21018\,
            I => \N__20998\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__21015\,
            I => \N__20998\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__21012\,
            I => \N__20998\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__21005\,
            I => un2_counter_9
        );

    \I__2436\ : Odrv4
    port map (
            O => \N__20998\,
            I => un2_counter_9
        );

    \I__2435\ : CascadeMux
    port map (
            O => \N__20993\,
            I => \clk_10khz_RNIIENAZ0Z2_cascade_\
        );

    \I__2434\ : InMux
    port map (
            O => \N__20990\,
            I => \N__20987\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__20987\,
            I => \N__20984\
        );

    \I__2432\ : Span4Mux_v
    port map (
            O => \N__20984\,
            I => \N__20981\
        );

    \I__2431\ : Odrv4
    port map (
            O => \N__20981\,
            I => \current_shift_inst.PI_CTRL.N_98\
        );

    \I__2430\ : CascadeMux
    port map (
            O => \N__20978\,
            I => \N__20975\
        );

    \I__2429\ : InMux
    port map (
            O => \N__20975\,
            I => \N__20972\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__20972\,
            I => \N__20969\
        );

    \I__2427\ : Span4Mux_h
    port map (
            O => \N__20969\,
            I => \N__20966\
        );

    \I__2426\ : Odrv4
    port map (
            O => \N__20966\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\
        );

    \I__2425\ : CascadeMux
    port map (
            O => \N__20963\,
            I => \N__20960\
        );

    \I__2424\ : InMux
    port map (
            O => \N__20960\,
            I => \N__20957\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__20957\,
            I => \N__20954\
        );

    \I__2422\ : Span4Mux_s2_h
    port map (
            O => \N__20954\,
            I => \N__20951\
        );

    \I__2421\ : Span4Mux_h
    port map (
            O => \N__20951\,
            I => \N__20948\
        );

    \I__2420\ : Odrv4
    port map (
            O => \N__20948\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\
        );

    \I__2419\ : InMux
    port map (
            O => \N__20945\,
            I => \N__20942\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__20942\,
            I => \N__20939\
        );

    \I__2417\ : Span4Mux_h
    port map (
            O => \N__20939\,
            I => \N__20936\
        );

    \I__2416\ : Odrv4
    port map (
            O => \N__20936\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\
        );

    \I__2415\ : InMux
    port map (
            O => \N__20933\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\
        );

    \I__2414\ : CascadeMux
    port map (
            O => \N__20930\,
            I => \N__20927\
        );

    \I__2413\ : InMux
    port map (
            O => \N__20927\,
            I => \N__20924\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__20924\,
            I => \N__20921\
        );

    \I__2411\ : Span4Mux_v
    port map (
            O => \N__20921\,
            I => \N__20918\
        );

    \I__2410\ : Odrv4
    port map (
            O => \N__20918\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\
        );

    \I__2409\ : InMux
    port map (
            O => \N__20915\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\
        );

    \I__2408\ : CascadeMux
    port map (
            O => \N__20912\,
            I => \N__20909\
        );

    \I__2407\ : InMux
    port map (
            O => \N__20909\,
            I => \N__20906\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__20906\,
            I => \N__20903\
        );

    \I__2405\ : Span4Mux_v
    port map (
            O => \N__20903\,
            I => \N__20900\
        );

    \I__2404\ : Odrv4
    port map (
            O => \N__20900\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\
        );

    \I__2403\ : InMux
    port map (
            O => \N__20897\,
            I => \N__20893\
        );

    \I__2402\ : InMux
    port map (
            O => \N__20896\,
            I => \N__20890\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__20893\,
            I => \N__20885\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__20890\,
            I => \N__20885\
        );

    \I__2399\ : Span4Mux_h
    port map (
            O => \N__20885\,
            I => \N__20881\
        );

    \I__2398\ : InMux
    port map (
            O => \N__20884\,
            I => \N__20878\
        );

    \I__2397\ : Odrv4
    port map (
            O => \N__20881\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__20878\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__2395\ : InMux
    port map (
            O => \N__20873\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\
        );

    \I__2394\ : InMux
    port map (
            O => \N__20870\,
            I => \N__20867\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__20867\,
            I => \N__20863\
        );

    \I__2392\ : InMux
    port map (
            O => \N__20866\,
            I => \N__20860\
        );

    \I__2391\ : Span4Mux_s3_h
    port map (
            O => \N__20863\,
            I => \N__20854\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__20860\,
            I => \N__20854\
        );

    \I__2389\ : InMux
    port map (
            O => \N__20859\,
            I => \N__20851\
        );

    \I__2388\ : Span4Mux_h
    port map (
            O => \N__20854\,
            I => \N__20846\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__20851\,
            I => \N__20846\
        );

    \I__2386\ : Span4Mux_v
    port map (
            O => \N__20846\,
            I => \N__20842\
        );

    \I__2385\ : InMux
    port map (
            O => \N__20845\,
            I => \N__20839\
        );

    \I__2384\ : Odrv4
    port map (
            O => \N__20842\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__20839\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__2382\ : InMux
    port map (
            O => \N__20834\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\
        );

    \I__2381\ : InMux
    port map (
            O => \N__20831\,
            I => \N__20828\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__20828\,
            I => \N__20825\
        );

    \I__2379\ : Glb2LocalMux
    port map (
            O => \N__20825\,
            I => \N__20822\
        );

    \I__2378\ : GlobalMux
    port map (
            O => \N__20822\,
            I => clk_12mhz
        );

    \I__2377\ : IoInMux
    port map (
            O => \N__20819\,
            I => \N__20816\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__20816\,
            I => \N__20813\
        );

    \I__2375\ : IoSpan4Mux
    port map (
            O => \N__20813\,
            I => \N__20810\
        );

    \I__2374\ : Span4Mux_s0_v
    port map (
            O => \N__20810\,
            I => \N__20807\
        );

    \I__2373\ : Odrv4
    port map (
            O => \N__20807\,
            I => \GB_BUFFER_clk_12mhz_THRU_CO\
        );

    \I__2372\ : InMux
    port map (
            O => \N__20804\,
            I => \N__20800\
        );

    \I__2371\ : InMux
    port map (
            O => \N__20803\,
            I => \N__20797\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__20800\,
            I => \counterZ0Z_4\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__20797\,
            I => \counterZ0Z_4\
        );

    \I__2368\ : InMux
    port map (
            O => \N__20792\,
            I => \N__20788\
        );

    \I__2367\ : InMux
    port map (
            O => \N__20791\,
            I => \N__20785\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__20788\,
            I => \counterZ0Z_3\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__20785\,
            I => \counterZ0Z_3\
        );

    \I__2364\ : InMux
    port map (
            O => \N__20780\,
            I => \N__20776\
        );

    \I__2363\ : InMux
    port map (
            O => \N__20779\,
            I => \N__20773\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__20776\,
            I => \counterZ0Z_5\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__20773\,
            I => \counterZ0Z_5\
        );

    \I__2360\ : InMux
    port map (
            O => \N__20768\,
            I => \N__20764\
        );

    \I__2359\ : InMux
    port map (
            O => \N__20767\,
            I => \N__20761\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__20764\,
            I => \counterZ0Z_6\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__20761\,
            I => \counterZ0Z_6\
        );

    \I__2356\ : CascadeMux
    port map (
            O => \N__20756\,
            I => \un2_counter_5_cascade_\
        );

    \I__2355\ : CascadeMux
    port map (
            O => \N__20753\,
            I => \N__20750\
        );

    \I__2354\ : InMux
    port map (
            O => \N__20750\,
            I => \N__20747\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__20747\,
            I => \counter_RNO_0Z0Z_12\
        );

    \I__2352\ : CascadeMux
    port map (
            O => \N__20744\,
            I => \N__20740\
        );

    \I__2351\ : InMux
    port map (
            O => \N__20743\,
            I => \N__20737\
        );

    \I__2350\ : InMux
    port map (
            O => \N__20740\,
            I => \N__20734\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__20737\,
            I => \counterZ0Z_12\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__20734\,
            I => \counterZ0Z_12\
        );

    \I__2347\ : CascadeMux
    port map (
            O => \N__20729\,
            I => \N__20726\
        );

    \I__2346\ : InMux
    port map (
            O => \N__20726\,
            I => \N__20723\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__20723\,
            I => \counter_RNO_0Z0Z_10\
        );

    \I__2344\ : CascadeMux
    port map (
            O => \N__20720\,
            I => \N__20716\
        );

    \I__2343\ : InMux
    port map (
            O => \N__20719\,
            I => \N__20713\
        );

    \I__2342\ : InMux
    port map (
            O => \N__20716\,
            I => \N__20710\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__20713\,
            I => \counterZ0Z_10\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__20710\,
            I => \counterZ0Z_10\
        );

    \I__2339\ : InMux
    port map (
            O => \N__20705\,
            I => \N__20700\
        );

    \I__2338\ : InMux
    port map (
            O => \N__20704\,
            I => \N__20697\
        );

    \I__2337\ : InMux
    port map (
            O => \N__20703\,
            I => \N__20694\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__20700\,
            I => \counterZ0Z_1\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__20697\,
            I => \counterZ0Z_1\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__20694\,
            I => \counterZ0Z_1\
        );

    \I__2333\ : CascadeMux
    port map (
            O => \N__20687\,
            I => \N__20682\
        );

    \I__2332\ : CascadeMux
    port map (
            O => \N__20686\,
            I => \N__20679\
        );

    \I__2331\ : InMux
    port map (
            O => \N__20685\,
            I => \N__20673\
        );

    \I__2330\ : InMux
    port map (
            O => \N__20682\,
            I => \N__20673\
        );

    \I__2329\ : InMux
    port map (
            O => \N__20679\,
            I => \N__20670\
        );

    \I__2328\ : InMux
    port map (
            O => \N__20678\,
            I => \N__20667\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__20673\,
            I => \counterZ0Z_0\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__20670\,
            I => \counterZ0Z_0\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__20667\,
            I => \counterZ0Z_0\
        );

    \I__2324\ : InMux
    port map (
            O => \N__20660\,
            I => \N__20657\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__20657\,
            I => \N__20654\
        );

    \I__2322\ : Odrv12
    port map (
            O => \N__20654\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_3\
        );

    \I__2321\ : InMux
    port map (
            O => \N__20651\,
            I => \N__20648\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__20648\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\
        );

    \I__2319\ : InMux
    port map (
            O => \N__20645\,
            I => \N__20642\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__20642\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6\
        );

    \I__2317\ : InMux
    port map (
            O => \N__20639\,
            I => \N__20636\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__20636\,
            I => \N__20633\
        );

    \I__2315\ : Odrv12
    port map (
            O => \N__20633\,
            I => \counter_RNO_0Z0Z_7\
        );

    \I__2314\ : InMux
    port map (
            O => \N__20630\,
            I => \N__20627\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__20627\,
            I => \N__20623\
        );

    \I__2312\ : InMux
    port map (
            O => \N__20626\,
            I => \N__20620\
        );

    \I__2311\ : Odrv4
    port map (
            O => \N__20623\,
            I => \counterZ0Z_7\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__20620\,
            I => \counterZ0Z_7\
        );

    \I__2309\ : InMux
    port map (
            O => \N__20615\,
            I => \N__20594\
        );

    \I__2308\ : InMux
    port map (
            O => \N__20614\,
            I => \N__20591\
        );

    \I__2307\ : InMux
    port map (
            O => \N__20613\,
            I => \N__20574\
        );

    \I__2306\ : InMux
    port map (
            O => \N__20612\,
            I => \N__20574\
        );

    \I__2305\ : InMux
    port map (
            O => \N__20611\,
            I => \N__20574\
        );

    \I__2304\ : InMux
    port map (
            O => \N__20610\,
            I => \N__20574\
        );

    \I__2303\ : InMux
    port map (
            O => \N__20609\,
            I => \N__20574\
        );

    \I__2302\ : InMux
    port map (
            O => \N__20608\,
            I => \N__20574\
        );

    \I__2301\ : InMux
    port map (
            O => \N__20607\,
            I => \N__20574\
        );

    \I__2300\ : InMux
    port map (
            O => \N__20606\,
            I => \N__20574\
        );

    \I__2299\ : InMux
    port map (
            O => \N__20605\,
            I => \N__20559\
        );

    \I__2298\ : InMux
    port map (
            O => \N__20604\,
            I => \N__20559\
        );

    \I__2297\ : InMux
    port map (
            O => \N__20603\,
            I => \N__20559\
        );

    \I__2296\ : InMux
    port map (
            O => \N__20602\,
            I => \N__20559\
        );

    \I__2295\ : InMux
    port map (
            O => \N__20601\,
            I => \N__20559\
        );

    \I__2294\ : InMux
    port map (
            O => \N__20600\,
            I => \N__20559\
        );

    \I__2293\ : InMux
    port map (
            O => \N__20599\,
            I => \N__20559\
        );

    \I__2292\ : InMux
    port map (
            O => \N__20598\,
            I => \N__20548\
        );

    \I__2291\ : InMux
    port map (
            O => \N__20597\,
            I => \N__20548\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__20594\,
            I => \N__20545\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__20591\,
            I => \N__20540\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__20574\,
            I => \N__20540\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__20559\,
            I => \N__20537\
        );

    \I__2286\ : InMux
    port map (
            O => \N__20558\,
            I => \N__20532\
        );

    \I__2285\ : InMux
    port map (
            O => \N__20557\,
            I => \N__20532\
        );

    \I__2284\ : CascadeMux
    port map (
            O => \N__20556\,
            I => \N__20526\
        );

    \I__2283\ : CascadeMux
    port map (
            O => \N__20555\,
            I => \N__20523\
        );

    \I__2282\ : CascadeMux
    port map (
            O => \N__20554\,
            I => \N__20520\
        );

    \I__2281\ : CascadeMux
    port map (
            O => \N__20553\,
            I => \N__20517\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__20548\,
            I => \N__20510\
        );

    \I__2279\ : Span4Mux_v
    port map (
            O => \N__20545\,
            I => \N__20503\
        );

    \I__2278\ : Span4Mux_v
    port map (
            O => \N__20540\,
            I => \N__20503\
        );

    \I__2277\ : Span4Mux_v
    port map (
            O => \N__20537\,
            I => \N__20503\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__20532\,
            I => \N__20500\
        );

    \I__2275\ : InMux
    port map (
            O => \N__20531\,
            I => \N__20493\
        );

    \I__2274\ : InMux
    port map (
            O => \N__20530\,
            I => \N__20493\
        );

    \I__2273\ : InMux
    port map (
            O => \N__20529\,
            I => \N__20493\
        );

    \I__2272\ : InMux
    port map (
            O => \N__20526\,
            I => \N__20488\
        );

    \I__2271\ : InMux
    port map (
            O => \N__20523\,
            I => \N__20488\
        );

    \I__2270\ : InMux
    port map (
            O => \N__20520\,
            I => \N__20483\
        );

    \I__2269\ : InMux
    port map (
            O => \N__20517\,
            I => \N__20483\
        );

    \I__2268\ : InMux
    port map (
            O => \N__20516\,
            I => \N__20474\
        );

    \I__2267\ : InMux
    port map (
            O => \N__20515\,
            I => \N__20474\
        );

    \I__2266\ : InMux
    port map (
            O => \N__20514\,
            I => \N__20474\
        );

    \I__2265\ : InMux
    port map (
            O => \N__20513\,
            I => \N__20474\
        );

    \I__2264\ : Span4Mux_v
    port map (
            O => \N__20510\,
            I => \N__20471\
        );

    \I__2263\ : Span4Mux_v
    port map (
            O => \N__20503\,
            I => \N__20466\
        );

    \I__2262\ : Span4Mux_s1_h
    port map (
            O => \N__20500\,
            I => \N__20466\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__20493\,
            I => \N__20463\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__20488\,
            I => \N_19_1\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__20483\,
            I => \N_19_1\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__20474\,
            I => \N_19_1\
        );

    \I__2257\ : Odrv4
    port map (
            O => \N__20471\,
            I => \N_19_1\
        );

    \I__2256\ : Odrv4
    port map (
            O => \N__20466\,
            I => \N_19_1\
        );

    \I__2255\ : Odrv12
    port map (
            O => \N__20463\,
            I => \N_19_1\
        );

    \I__2254\ : InMux
    port map (
            O => \N__20450\,
            I => \N__20432\
        );

    \I__2253\ : InMux
    port map (
            O => \N__20449\,
            I => \N__20432\
        );

    \I__2252\ : InMux
    port map (
            O => \N__20448\,
            I => \N__20432\
        );

    \I__2251\ : InMux
    port map (
            O => \N__20447\,
            I => \N__20432\
        );

    \I__2250\ : InMux
    port map (
            O => \N__20446\,
            I => \N__20432\
        );

    \I__2249\ : InMux
    port map (
            O => \N__20445\,
            I => \N__20432\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__20432\,
            I => \N__20427\
        );

    \I__2247\ : InMux
    port map (
            O => \N__20431\,
            I => \N__20422\
        );

    \I__2246\ : InMux
    port map (
            O => \N__20430\,
            I => \N__20422\
        );

    \I__2245\ : Span4Mux_v
    port map (
            O => \N__20427\,
            I => \N__20417\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__20422\,
            I => \N__20414\
        );

    \I__2243\ : InMux
    port map (
            O => \N__20421\,
            I => \N__20409\
        );

    \I__2242\ : InMux
    port map (
            O => \N__20420\,
            I => \N__20409\
        );

    \I__2241\ : Odrv4
    port map (
            O => \N__20417\,
            I => \pwm_generator_inst.N_17\
        );

    \I__2240\ : Odrv12
    port map (
            O => \N__20414\,
            I => \pwm_generator_inst.N_17\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__20409\,
            I => \pwm_generator_inst.N_17\
        );

    \I__2238\ : InMux
    port map (
            O => \N__20402\,
            I => \N__20392\
        );

    \I__2237\ : InMux
    port map (
            O => \N__20401\,
            I => \N__20392\
        );

    \I__2236\ : CascadeMux
    port map (
            O => \N__20400\,
            I => \N__20389\
        );

    \I__2235\ : CascadeMux
    port map (
            O => \N__20399\,
            I => \N__20386\
        );

    \I__2234\ : CascadeMux
    port map (
            O => \N__20398\,
            I => \N__20383\
        );

    \I__2233\ : CascadeMux
    port map (
            O => \N__20397\,
            I => \N__20380\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__20392\,
            I => \N__20375\
        );

    \I__2231\ : InMux
    port map (
            O => \N__20389\,
            I => \N__20362\
        );

    \I__2230\ : InMux
    port map (
            O => \N__20386\,
            I => \N__20362\
        );

    \I__2229\ : InMux
    port map (
            O => \N__20383\,
            I => \N__20362\
        );

    \I__2228\ : InMux
    port map (
            O => \N__20380\,
            I => \N__20362\
        );

    \I__2227\ : InMux
    port map (
            O => \N__20379\,
            I => \N__20362\
        );

    \I__2226\ : InMux
    port map (
            O => \N__20378\,
            I => \N__20362\
        );

    \I__2225\ : Span4Mux_v
    port map (
            O => \N__20375\,
            I => \N__20357\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__20362\,
            I => \N__20354\
        );

    \I__2223\ : InMux
    port map (
            O => \N__20361\,
            I => \N__20349\
        );

    \I__2222\ : InMux
    port map (
            O => \N__20360\,
            I => \N__20349\
        );

    \I__2221\ : Odrv4
    port map (
            O => \N__20357\,
            I => \pwm_generator_inst.N_16\
        );

    \I__2220\ : Odrv4
    port map (
            O => \N__20354\,
            I => \pwm_generator_inst.N_16\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__20349\,
            I => \pwm_generator_inst.N_16\
        );

    \I__2218\ : InMux
    port map (
            O => \N__20342\,
            I => \N__20339\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__20339\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7\
        );

    \I__2216\ : CascadeMux
    port map (
            O => \N__20336\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_\
        );

    \I__2215\ : InMux
    port map (
            O => \N__20333\,
            I => \N__20330\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__20330\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\
        );

    \I__2213\ : InMux
    port map (
            O => \N__20327\,
            I => \N__20324\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__20324\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\
        );

    \I__2211\ : InMux
    port map (
            O => \N__20321\,
            I => un5_counter_cry_9
        );

    \I__2210\ : InMux
    port map (
            O => \N__20318\,
            I => un5_counter_cry_10
        );

    \I__2209\ : InMux
    port map (
            O => \N__20315\,
            I => un5_counter_cry_11
        );

    \I__2208\ : InMux
    port map (
            O => \N__20312\,
            I => \N__20308\
        );

    \I__2207\ : InMux
    port map (
            O => \N__20311\,
            I => \N__20305\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__20308\,
            I => \N__20302\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__20305\,
            I => \counterZ0Z_11\
        );

    \I__2204\ : Odrv4
    port map (
            O => \N__20302\,
            I => \counterZ0Z_11\
        );

    \I__2203\ : InMux
    port map (
            O => \N__20297\,
            I => \N__20293\
        );

    \I__2202\ : InMux
    port map (
            O => \N__20296\,
            I => \N__20290\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__20293\,
            I => \counterZ0Z_9\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__20290\,
            I => \counterZ0Z_9\
        );

    \I__2199\ : InMux
    port map (
            O => \N__20285\,
            I => \N__20281\
        );

    \I__2198\ : InMux
    port map (
            O => \N__20284\,
            I => \N__20278\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__20281\,
            I => \N__20275\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__20278\,
            I => \counterZ0Z_8\
        );

    \I__2195\ : Odrv4
    port map (
            O => \N__20275\,
            I => \counterZ0Z_8\
        );

    \I__2194\ : InMux
    port map (
            O => \N__20270\,
            I => \N__20266\
        );

    \I__2193\ : InMux
    port map (
            O => \N__20269\,
            I => \N__20263\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__20266\,
            I => \N__20260\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__20263\,
            I => \counterZ0Z_2\
        );

    \I__2190\ : Odrv4
    port map (
            O => \N__20260\,
            I => \counterZ0Z_2\
        );

    \I__2189\ : InMux
    port map (
            O => \N__20255\,
            I => \N__20252\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__20252\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4\
        );

    \I__2187\ : InMux
    port map (
            O => \N__20249\,
            I => \N__20246\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__20246\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1\
        );

    \I__2185\ : InMux
    port map (
            O => \N__20243\,
            I => \N__20240\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__20240\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5\
        );

    \I__2183\ : InMux
    port map (
            O => \N__20237\,
            I => \N__20234\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__20234\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0\
        );

    \I__2181\ : InMux
    port map (
            O => \N__20231\,
            I => un5_counter_cry_1
        );

    \I__2180\ : InMux
    port map (
            O => \N__20228\,
            I => un5_counter_cry_2
        );

    \I__2179\ : InMux
    port map (
            O => \N__20225\,
            I => un5_counter_cry_3
        );

    \I__2178\ : InMux
    port map (
            O => \N__20222\,
            I => un5_counter_cry_4
        );

    \I__2177\ : InMux
    port map (
            O => \N__20219\,
            I => un5_counter_cry_5
        );

    \I__2176\ : InMux
    port map (
            O => \N__20216\,
            I => un5_counter_cry_6
        );

    \I__2175\ : InMux
    port map (
            O => \N__20213\,
            I => un5_counter_cry_7
        );

    \I__2174\ : InMux
    port map (
            O => \N__20210\,
            I => \bfn_4_6_0_\
        );

    \I__2173\ : CascadeMux
    port map (
            O => \N__20207\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_9_9_cascade_\
        );

    \I__2172\ : InMux
    port map (
            O => \N__20204\,
            I => \N__20201\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__20201\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\
        );

    \I__2170\ : InMux
    port map (
            O => \N__20198\,
            I => \N__20195\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__20195\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\
        );

    \I__2168\ : CascadeMux
    port map (
            O => \N__20192\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_\
        );

    \I__2167\ : InMux
    port map (
            O => \N__20189\,
            I => \N__20186\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__20186\,
            I => \N__20183\
        );

    \I__2165\ : Odrv4
    port map (
            O => \N__20183\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\
        );

    \I__2164\ : CascadeMux
    port map (
            O => \N__20180\,
            I => \N__20177\
        );

    \I__2163\ : InMux
    port map (
            O => \N__20177\,
            I => \N__20174\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__20174\,
            I => \N__20171\
        );

    \I__2161\ : Odrv4
    port map (
            O => \N__20171\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\
        );

    \I__2160\ : InMux
    port map (
            O => \N__20168\,
            I => \N__20164\
        );

    \I__2159\ : InMux
    port map (
            O => \N__20167\,
            I => \N__20160\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__20164\,
            I => \N__20157\
        );

    \I__2157\ : InMux
    port map (
            O => \N__20163\,
            I => \N__20154\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__20160\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_13\
        );

    \I__2155\ : Odrv4
    port map (
            O => \N__20157\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_13\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__20154\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_13\
        );

    \I__2153\ : InMux
    port map (
            O => \N__20147\,
            I => \N__20144\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__20144\,
            I => \N__20141\
        );

    \I__2151\ : Span4Mux_v
    port map (
            O => \N__20141\,
            I => \N__20137\
        );

    \I__2150\ : InMux
    port map (
            O => \N__20140\,
            I => \N__20134\
        );

    \I__2149\ : Odrv4
    port map (
            O => \N__20137\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__20134\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\
        );

    \I__2147\ : CascadeMux
    port map (
            O => \N__20129\,
            I => \N__20126\
        );

    \I__2146\ : InMux
    port map (
            O => \N__20126\,
            I => \N__20123\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__20123\,
            I => \N__20120\
        );

    \I__2144\ : Span4Mux_h
    port map (
            O => \N__20120\,
            I => \N__20117\
        );

    \I__2143\ : Span4Mux_v
    port map (
            O => \N__20117\,
            I => \N__20114\
        );

    \I__2142\ : Odrv4
    port map (
            O => \N__20114\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO\
        );

    \I__2141\ : InMux
    port map (
            O => \N__20111\,
            I => \N__20108\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__20108\,
            I => \N__20105\
        );

    \I__2139\ : Span4Mux_h
    port map (
            O => \N__20105\,
            I => \N__20102\
        );

    \I__2138\ : Odrv4
    port map (
            O => \N__20102\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_3\
        );

    \I__2137\ : InMux
    port map (
            O => \N__20099\,
            I => \N__20094\
        );

    \I__2136\ : InMux
    port map (
            O => \N__20098\,
            I => \N__20091\
        );

    \I__2135\ : InMux
    port map (
            O => \N__20097\,
            I => \N__20088\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__20094\,
            I => \N__20085\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__20091\,
            I => \N__20082\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__20088\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_12\
        );

    \I__2131\ : Odrv4
    port map (
            O => \N__20085\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_12\
        );

    \I__2130\ : Odrv4
    port map (
            O => \N__20082\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_12\
        );

    \I__2129\ : InMux
    port map (
            O => \N__20075\,
            I => \N__20072\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__20072\,
            I => \N__20069\
        );

    \I__2127\ : Span4Mux_h
    port map (
            O => \N__20069\,
            I => \N__20065\
        );

    \I__2126\ : InMux
    port map (
            O => \N__20068\,
            I => \N__20062\
        );

    \I__2125\ : Odrv4
    port map (
            O => \N__20065\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__20062\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\
        );

    \I__2123\ : CascadeMux
    port map (
            O => \N__20057\,
            I => \N__20054\
        );

    \I__2122\ : InMux
    port map (
            O => \N__20054\,
            I => \N__20051\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__20051\,
            I => \N__20048\
        );

    \I__2120\ : Span4Mux_v
    port map (
            O => \N__20048\,
            I => \N__20045\
        );

    \I__2119\ : Odrv4
    port map (
            O => \N__20045\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO\
        );

    \I__2118\ : CascadeMux
    port map (
            O => \N__20042\,
            I => \N__20037\
        );

    \I__2117\ : InMux
    port map (
            O => \N__20041\,
            I => \N__20027\
        );

    \I__2116\ : InMux
    port map (
            O => \N__20040\,
            I => \N__20024\
        );

    \I__2115\ : InMux
    port map (
            O => \N__20037\,
            I => \N__20021\
        );

    \I__2114\ : InMux
    port map (
            O => \N__20036\,
            I => \N__20012\
        );

    \I__2113\ : InMux
    port map (
            O => \N__20035\,
            I => \N__20012\
        );

    \I__2112\ : InMux
    port map (
            O => \N__20034\,
            I => \N__20012\
        );

    \I__2111\ : InMux
    port map (
            O => \N__20033\,
            I => \N__20012\
        );

    \I__2110\ : InMux
    port map (
            O => \N__20032\,
            I => \N__20007\
        );

    \I__2109\ : InMux
    port map (
            O => \N__20031\,
            I => \N__20007\
        );

    \I__2108\ : InMux
    port map (
            O => \N__20030\,
            I => \N__20004\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__20027\,
            I => \N__19997\
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__20024\,
            I => \N__19997\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__20021\,
            I => \N__19997\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__20012\,
            I => \N__19990\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__20007\,
            I => \N__19990\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__20004\,
            I => \N__19987\
        );

    \I__2101\ : Span4Mux_v
    port map (
            O => \N__19997\,
            I => \N__19984\
        );

    \I__2100\ : InMux
    port map (
            O => \N__19996\,
            I => \N__19979\
        );

    \I__2099\ : InMux
    port map (
            O => \N__19995\,
            I => \N__19979\
        );

    \I__2098\ : Span4Mux_v
    port map (
            O => \N__19990\,
            I => \N__19974\
        );

    \I__2097\ : Span4Mux_v
    port map (
            O => \N__19987\,
            I => \N__19974\
        );

    \I__2096\ : Odrv4
    port map (
            O => \N__19984\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__19979\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2094\ : Odrv4
    port map (
            O => \N__19974\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2093\ : InMux
    port map (
            O => \N__19967\,
            I => \N__19964\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__19964\,
            I => \N__19961\
        );

    \I__2091\ : Odrv12
    port map (
            O => \N__19961\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_2\
        );

    \I__2090\ : InMux
    port map (
            O => \N__19958\,
            I => \N__19955\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__19955\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_7\
        );

    \I__2088\ : InMux
    port map (
            O => \N__19952\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_6\
        );

    \I__2087\ : CascadeMux
    port map (
            O => \N__19949\,
            I => \N__19946\
        );

    \I__2086\ : InMux
    port map (
            O => \N__19946\,
            I => \N__19943\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__19943\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_8\
        );

    \I__2084\ : CascadeMux
    port map (
            O => \N__19940\,
            I => \N__19937\
        );

    \I__2083\ : InMux
    port map (
            O => \N__19937\,
            I => \N__19934\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__19934\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8\
        );

    \I__2081\ : InMux
    port map (
            O => \N__19931\,
            I => \bfn_3_9_0_\
        );

    \I__2080\ : InMux
    port map (
            O => \N__19928\,
            I => \N__19925\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__19925\,
            I => \N__19922\
        );

    \I__2078\ : Odrv4
    port map (
            O => \N__19922\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO\
        );

    \I__2077\ : CascadeMux
    port map (
            O => \N__19919\,
            I => \N__19916\
        );

    \I__2076\ : InMux
    port map (
            O => \N__19916\,
            I => \N__19913\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__19913\,
            I => \N__19910\
        );

    \I__2074\ : Span4Mux_h
    port map (
            O => \N__19910\,
            I => \N__19907\
        );

    \I__2073\ : Odrv4
    port map (
            O => \N__19907\,
            I => \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9\
        );

    \I__2072\ : InMux
    port map (
            O => \N__19904\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_8\
        );

    \I__2071\ : CascadeMux
    port map (
            O => \N__19901\,
            I => \N__19898\
        );

    \I__2070\ : InMux
    port map (
            O => \N__19898\,
            I => \N__19895\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__19895\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9\
        );

    \I__2068\ : InMux
    port map (
            O => \N__19892\,
            I => \N__19882\
        );

    \I__2067\ : InMux
    port map (
            O => \N__19891\,
            I => \N__19877\
        );

    \I__2066\ : InMux
    port map (
            O => \N__19890\,
            I => \N__19877\
        );

    \I__2065\ : InMux
    port map (
            O => \N__19889\,
            I => \N__19872\
        );

    \I__2064\ : InMux
    port map (
            O => \N__19888\,
            I => \N__19872\
        );

    \I__2063\ : InMux
    port map (
            O => \N__19887\,
            I => \N__19867\
        );

    \I__2062\ : InMux
    port map (
            O => \N__19886\,
            I => \N__19867\
        );

    \I__2061\ : InMux
    port map (
            O => \N__19885\,
            I => \N__19864\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__19882\,
            I => \N__19858\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__19877\,
            I => \N__19858\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__19872\,
            I => \N__19855\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__19867\,
            I => \N__19850\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__19864\,
            I => \N__19850\
        );

    \I__2055\ : InMux
    port map (
            O => \N__19863\,
            I => \N__19847\
        );

    \I__2054\ : Span12Mux_s8_v
    port map (
            O => \N__19858\,
            I => \N__19844\
        );

    \I__2053\ : Span4Mux_v
    port map (
            O => \N__19855\,
            I => \N__19839\
        );

    \I__2052\ : Span4Mux_s3_h
    port map (
            O => \N__19850\,
            I => \N__19839\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__19847\,
            I => \N__19836\
        );

    \I__2050\ : Odrv12
    port map (
            O => \N__19844\,
            I => \current_shift_inst.PI_CTRL.N_178\
        );

    \I__2049\ : Odrv4
    port map (
            O => \N__19839\,
            I => \current_shift_inst.PI_CTRL.N_178\
        );

    \I__2048\ : Odrv12
    port map (
            O => \N__19836\,
            I => \current_shift_inst.PI_CTRL.N_178\
        );

    \I__2047\ : InMux
    port map (
            O => \N__19829\,
            I => \N__19823\
        );

    \I__2046\ : InMux
    port map (
            O => \N__19828\,
            I => \N__19816\
        );

    \I__2045\ : InMux
    port map (
            O => \N__19827\,
            I => \N__19816\
        );

    \I__2044\ : InMux
    port map (
            O => \N__19826\,
            I => \N__19816\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__19823\,
            I => \N__19810\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__19816\,
            I => \N__19807\
        );

    \I__2041\ : InMux
    port map (
            O => \N__19815\,
            I => \N__19802\
        );

    \I__2040\ : InMux
    port map (
            O => \N__19814\,
            I => \N__19802\
        );

    \I__2039\ : InMux
    port map (
            O => \N__19813\,
            I => \N__19799\
        );

    \I__2038\ : Span4Mux_v
    port map (
            O => \N__19810\,
            I => \N__19794\
        );

    \I__2037\ : Span4Mux_s2_h
    port map (
            O => \N__19807\,
            I => \N__19794\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__19802\,
            I => \N__19791\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__19799\,
            I => \N__19788\
        );

    \I__2034\ : Span4Mux_v
    port map (
            O => \N__19794\,
            I => \N__19785\
        );

    \I__2033\ : Span4Mux_v
    port map (
            O => \N__19791\,
            I => \N__19780\
        );

    \I__2032\ : Span4Mux_s3_h
    port map (
            O => \N__19788\,
            I => \N__19780\
        );

    \I__2031\ : Odrv4
    port map (
            O => \N__19785\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__2030\ : Odrv4
    port map (
            O => \N__19780\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__2029\ : InMux
    port map (
            O => \N__19775\,
            I => \N__19772\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__19772\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\
        );

    \I__2027\ : CascadeMux
    port map (
            O => \N__19769\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\
        );

    \I__2026\ : InMux
    port map (
            O => \N__19766\,
            I => \N__19763\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__19763\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\
        );

    \I__2024\ : CascadeMux
    port map (
            O => \N__19760\,
            I => \N__19757\
        );

    \I__2023\ : InMux
    port map (
            O => \N__19757\,
            I => \N__19754\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__19754\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\
        );

    \I__2021\ : InMux
    port map (
            O => \N__19751\,
            I => \N__19748\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__19748\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_0\
        );

    \I__2019\ : CascadeMux
    port map (
            O => \N__19745\,
            I => \N__19742\
        );

    \I__2018\ : InMux
    port map (
            O => \N__19742\,
            I => \N__19739\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__19739\,
            I => \N__19736\
        );

    \I__2016\ : Odrv4
    port map (
            O => \N__19736\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_1\
        );

    \I__2015\ : InMux
    port map (
            O => \N__19733\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_0\
        );

    \I__2014\ : InMux
    port map (
            O => \N__19730\,
            I => \N__19727\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__19727\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2\
        );

    \I__2012\ : InMux
    port map (
            O => \N__19724\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_1\
        );

    \I__2011\ : InMux
    port map (
            O => \N__19721\,
            I => \N__19718\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__19718\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3\
        );

    \I__2009\ : InMux
    port map (
            O => \N__19715\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_2\
        );

    \I__2008\ : InMux
    port map (
            O => \N__19712\,
            I => \N__19709\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__19709\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_4\
        );

    \I__2006\ : InMux
    port map (
            O => \N__19706\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_3\
        );

    \I__2005\ : InMux
    port map (
            O => \N__19703\,
            I => \N__19700\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__19700\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_5\
        );

    \I__2003\ : InMux
    port map (
            O => \N__19697\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_4\
        );

    \I__2002\ : InMux
    port map (
            O => \N__19694\,
            I => \N__19691\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__19691\,
            I => \N__19688\
        );

    \I__2000\ : Odrv4
    port map (
            O => \N__19688\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_6\
        );

    \I__1999\ : InMux
    port map (
            O => \N__19685\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_5\
        );

    \I__1998\ : InMux
    port map (
            O => \N__19682\,
            I => \N__19679\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__19679\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0\
        );

    \I__1996\ : InMux
    port map (
            O => \N__19676\,
            I => \N__19669\
        );

    \I__1995\ : CascadeMux
    port map (
            O => \N__19675\,
            I => \N__19666\
        );

    \I__1994\ : CascadeMux
    port map (
            O => \N__19674\,
            I => \N__19662\
        );

    \I__1993\ : CascadeMux
    port map (
            O => \N__19673\,
            I => \N__19658\
        );

    \I__1992\ : InMux
    port map (
            O => \N__19672\,
            I => \N__19654\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__19669\,
            I => \N__19651\
        );

    \I__1990\ : InMux
    port map (
            O => \N__19666\,
            I => \N__19638\
        );

    \I__1989\ : InMux
    port map (
            O => \N__19665\,
            I => \N__19638\
        );

    \I__1988\ : InMux
    port map (
            O => \N__19662\,
            I => \N__19638\
        );

    \I__1987\ : InMux
    port map (
            O => \N__19661\,
            I => \N__19638\
        );

    \I__1986\ : InMux
    port map (
            O => \N__19658\,
            I => \N__19638\
        );

    \I__1985\ : InMux
    port map (
            O => \N__19657\,
            I => \N__19638\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__19654\,
            I => \N__19631\
        );

    \I__1983\ : Span4Mux_v
    port map (
            O => \N__19651\,
            I => \N__19631\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__19638\,
            I => \N__19631\
        );

    \I__1981\ : Span4Mux_v
    port map (
            O => \N__19631\,
            I => \N__19628\
        );

    \I__1980\ : Odrv4
    port map (
            O => \N__19628\,
            I => \pwm_generator_inst.un2_threshold_acc_1_25\
        );

    \I__1979\ : InMux
    port map (
            O => \N__19625\,
            I => \N__19622\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__19622\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0\
        );

    \I__1977\ : InMux
    port map (
            O => \N__19619\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\
        );

    \I__1976\ : InMux
    port map (
            O => \N__19616\,
            I => \N__19613\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__19613\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO\
        );

    \I__1974\ : InMux
    port map (
            O => \N__19610\,
            I => \N__19607\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__19607\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16\
        );

    \I__1972\ : InMux
    port map (
            O => \N__19604\,
            I => \bfn_2_13_0_\
        );

    \I__1971\ : InMux
    port map (
            O => \N__19601\,
            I => \N__19598\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__19598\,
            I => \N__19595\
        );

    \I__1969\ : Span4Mux_s1_v
    port map (
            O => \N__19595\,
            I => \N__19592\
        );

    \I__1968\ : Odrv4
    port map (
            O => \N__19592\,
            I => \N_32_i_i\
        );

    \I__1967\ : InMux
    port map (
            O => \N__19589\,
            I => \N__19586\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__19586\,
            I => \N__19583\
        );

    \I__1965\ : Odrv4
    port map (
            O => \N__19583\,
            I => \current_shift_inst.PI_CTRL.N_91\
        );

    \I__1964\ : CascadeMux
    port map (
            O => \N__19580\,
            I => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\
        );

    \I__1963\ : InMux
    port map (
            O => \N__19577\,
            I => \N__19572\
        );

    \I__1962\ : InMux
    port map (
            O => \N__19576\,
            I => \N__19567\
        );

    \I__1961\ : InMux
    port map (
            O => \N__19575\,
            I => \N__19567\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__19572\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__19567\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__1958\ : InMux
    port map (
            O => \N__19562\,
            I => \N__19559\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__19559\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\
        );

    \I__1956\ : InMux
    port map (
            O => \N__19556\,
            I => \N__19552\
        );

    \I__1955\ : InMux
    port map (
            O => \N__19555\,
            I => \N__19548\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__19552\,
            I => \N__19545\
        );

    \I__1953\ : InMux
    port map (
            O => \N__19551\,
            I => \N__19542\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__19548\,
            I => pwm_duty_input_3
        );

    \I__1951\ : Odrv4
    port map (
            O => \N__19545\,
            I => pwm_duty_input_3
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__19542\,
            I => pwm_duty_input_3
        );

    \I__1949\ : CascadeMux
    port map (
            O => \N__19535\,
            I => \N__19532\
        );

    \I__1948\ : InMux
    port map (
            O => \N__19532\,
            I => \N__19529\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__19529\,
            I => \pwm_generator_inst.un1_duty_inputlt3\
        );

    \I__1946\ : InMux
    port map (
            O => \N__19526\,
            I => \N__19522\
        );

    \I__1945\ : InMux
    port map (
            O => \N__19525\,
            I => \N__19519\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__19522\,
            I => \N__19515\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__19519\,
            I => \N__19512\
        );

    \I__1942\ : InMux
    port map (
            O => \N__19518\,
            I => \N__19509\
        );

    \I__1941\ : Span4Mux_v
    port map (
            O => \N__19515\,
            I => \N__19504\
        );

    \I__1940\ : Span4Mux_v
    port map (
            O => \N__19512\,
            I => \N__19504\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__19509\,
            I => pwm_duty_input_4
        );

    \I__1938\ : Odrv4
    port map (
            O => \N__19504\,
            I => pwm_duty_input_4
        );

    \I__1937\ : InMux
    port map (
            O => \N__19499\,
            I => \N__19496\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__19496\,
            I => \N__19493\
        );

    \I__1935\ : Span4Mux_v
    port map (
            O => \N__19493\,
            I => \N__19490\
        );

    \I__1934\ : Odrv4
    port map (
            O => \N__19490\,
            I => \pwm_generator_inst.un2_threshold_acc_1_22\
        );

    \I__1933\ : CascadeMux
    port map (
            O => \N__19487\,
            I => \N__19484\
        );

    \I__1932\ : InMux
    port map (
            O => \N__19484\,
            I => \N__19481\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__19481\,
            I => \N__19478\
        );

    \I__1930\ : Span4Mux_h
    port map (
            O => \N__19478\,
            I => \N__19475\
        );

    \I__1929\ : Odrv4
    port map (
            O => \N__19475\,
            I => \pwm_generator_inst.un2_threshold_acc_2_7\
        );

    \I__1928\ : InMux
    port map (
            O => \N__19472\,
            I => \N__19469\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__19469\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0\
        );

    \I__1926\ : InMux
    port map (
            O => \N__19466\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\
        );

    \I__1925\ : InMux
    port map (
            O => \N__19463\,
            I => \N__19460\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__19460\,
            I => \N__19457\
        );

    \I__1923\ : Span4Mux_h
    port map (
            O => \N__19457\,
            I => \N__19454\
        );

    \I__1922\ : Span4Mux_v
    port map (
            O => \N__19454\,
            I => \N__19451\
        );

    \I__1921\ : Odrv4
    port map (
            O => \N__19451\,
            I => \pwm_generator_inst.un2_threshold_acc_1_23\
        );

    \I__1920\ : CascadeMux
    port map (
            O => \N__19448\,
            I => \N__19445\
        );

    \I__1919\ : InMux
    port map (
            O => \N__19445\,
            I => \N__19442\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__19442\,
            I => \N__19439\
        );

    \I__1917\ : Span4Mux_h
    port map (
            O => \N__19439\,
            I => \N__19436\
        );

    \I__1916\ : Odrv4
    port map (
            O => \N__19436\,
            I => \pwm_generator_inst.un2_threshold_acc_2_8\
        );

    \I__1915\ : InMux
    port map (
            O => \N__19433\,
            I => \N__19430\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__19430\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0\
        );

    \I__1913\ : InMux
    port map (
            O => \N__19427\,
            I => \bfn_2_12_0_\
        );

    \I__1912\ : InMux
    port map (
            O => \N__19424\,
            I => \N__19421\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__19421\,
            I => \N__19418\
        );

    \I__1910\ : Span4Mux_v
    port map (
            O => \N__19418\,
            I => \N__19415\
        );

    \I__1909\ : Odrv4
    port map (
            O => \N__19415\,
            I => \pwm_generator_inst.un2_threshold_acc_1_24\
        );

    \I__1908\ : CascadeMux
    port map (
            O => \N__19412\,
            I => \N__19409\
        );

    \I__1907\ : InMux
    port map (
            O => \N__19409\,
            I => \N__19406\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__19406\,
            I => \N__19403\
        );

    \I__1905\ : Span4Mux_h
    port map (
            O => \N__19403\,
            I => \N__19400\
        );

    \I__1904\ : Odrv4
    port map (
            O => \N__19400\,
            I => \pwm_generator_inst.un2_threshold_acc_2_9\
        );

    \I__1903\ : InMux
    port map (
            O => \N__19397\,
            I => \N__19394\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__19394\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0\
        );

    \I__1901\ : InMux
    port map (
            O => \N__19391\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\
        );

    \I__1900\ : CascadeMux
    port map (
            O => \N__19388\,
            I => \N__19385\
        );

    \I__1899\ : InMux
    port map (
            O => \N__19385\,
            I => \N__19382\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__19382\,
            I => \N__19379\
        );

    \I__1897\ : Span4Mux_h
    port map (
            O => \N__19379\,
            I => \N__19376\
        );

    \I__1896\ : Odrv4
    port map (
            O => \N__19376\,
            I => \pwm_generator_inst.un2_threshold_acc_2_10\
        );

    \I__1895\ : InMux
    port map (
            O => \N__19373\,
            I => \N__19370\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__19370\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0\
        );

    \I__1893\ : InMux
    port map (
            O => \N__19367\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\
        );

    \I__1892\ : InMux
    port map (
            O => \N__19364\,
            I => \N__19361\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__19361\,
            I => \N__19358\
        );

    \I__1890\ : Span4Mux_h
    port map (
            O => \N__19358\,
            I => \N__19355\
        );

    \I__1889\ : Odrv4
    port map (
            O => \N__19355\,
            I => \pwm_generator_inst.un2_threshold_acc_2_11\
        );

    \I__1888\ : InMux
    port map (
            O => \N__19352\,
            I => \N__19349\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__19349\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0\
        );

    \I__1886\ : InMux
    port map (
            O => \N__19346\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\
        );

    \I__1885\ : CascadeMux
    port map (
            O => \N__19343\,
            I => \N__19340\
        );

    \I__1884\ : InMux
    port map (
            O => \N__19340\,
            I => \N__19337\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__19337\,
            I => \N__19334\
        );

    \I__1882\ : Span4Mux_v
    port map (
            O => \N__19334\,
            I => \N__19331\
        );

    \I__1881\ : Odrv4
    port map (
            O => \N__19331\,
            I => \pwm_generator_inst.un2_threshold_acc_2_12\
        );

    \I__1880\ : InMux
    port map (
            O => \N__19328\,
            I => \N__19325\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__19325\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0\
        );

    \I__1878\ : InMux
    port map (
            O => \N__19322\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\
        );

    \I__1877\ : InMux
    port map (
            O => \N__19319\,
            I => \N__19316\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__19316\,
            I => \N__19313\
        );

    \I__1875\ : Span4Mux_v
    port map (
            O => \N__19313\,
            I => \N__19310\
        );

    \I__1874\ : Odrv4
    port map (
            O => \N__19310\,
            I => \pwm_generator_inst.un2_threshold_acc_2_13\
        );

    \I__1873\ : InMux
    port map (
            O => \N__19307\,
            I => \N__19304\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__19304\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0\
        );

    \I__1871\ : InMux
    port map (
            O => \N__19301\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\
        );

    \I__1870\ : CascadeMux
    port map (
            O => \N__19298\,
            I => \N__19295\
        );

    \I__1869\ : InMux
    port map (
            O => \N__19295\,
            I => \N__19292\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__19292\,
            I => \N__19289\
        );

    \I__1867\ : Span4Mux_h
    port map (
            O => \N__19289\,
            I => \N__19286\
        );

    \I__1866\ : Odrv4
    port map (
            O => \N__19286\,
            I => \pwm_generator_inst.un2_threshold_acc_2_14\
        );

    \I__1865\ : InMux
    port map (
            O => \N__19283\,
            I => \N__19280\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__19280\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0\
        );

    \I__1863\ : InMux
    port map (
            O => \N__19277\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\
        );

    \I__1862\ : InMux
    port map (
            O => \N__19274\,
            I => \N__19271\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__19271\,
            I => \N__19268\
        );

    \I__1860\ : Span4Mux_h
    port map (
            O => \N__19268\,
            I => \N__19265\
        );

    \I__1859\ : Odrv4
    port map (
            O => \N__19265\,
            I => \pwm_generator_inst.un2_threshold_acc_2_0\
        );

    \I__1858\ : CascadeMux
    port map (
            O => \N__19262\,
            I => \N__19259\
        );

    \I__1857\ : InMux
    port map (
            O => \N__19259\,
            I => \N__19256\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__19256\,
            I => \N__19253\
        );

    \I__1855\ : Span4Mux_h
    port map (
            O => \N__19253\,
            I => \N__19250\
        );

    \I__1854\ : Span4Mux_v
    port map (
            O => \N__19250\,
            I => \N__19247\
        );

    \I__1853\ : Odrv4
    port map (
            O => \N__19247\,
            I => \pwm_generator_inst.un2_threshold_acc_1_15\
        );

    \I__1852\ : InMux
    port map (
            O => \N__19244\,
            I => \N__19241\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__19241\,
            I => \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4\
        );

    \I__1850\ : InMux
    port map (
            O => \N__19238\,
            I => \N__19235\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__19235\,
            I => \N__19232\
        );

    \I__1848\ : Span4Mux_v
    port map (
            O => \N__19232\,
            I => \N__19229\
        );

    \I__1847\ : Odrv4
    port map (
            O => \N__19229\,
            I => \pwm_generator_inst.un2_threshold_acc_1_16\
        );

    \I__1846\ : CascadeMux
    port map (
            O => \N__19226\,
            I => \N__19223\
        );

    \I__1845\ : InMux
    port map (
            O => \N__19223\,
            I => \N__19220\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__19220\,
            I => \N__19217\
        );

    \I__1843\ : Span4Mux_h
    port map (
            O => \N__19217\,
            I => \N__19214\
        );

    \I__1842\ : Odrv4
    port map (
            O => \N__19214\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1\
        );

    \I__1841\ : CascadeMux
    port map (
            O => \N__19211\,
            I => \N__19208\
        );

    \I__1840\ : InMux
    port map (
            O => \N__19208\,
            I => \N__19205\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__19205\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0\
        );

    \I__1838\ : InMux
    port map (
            O => \N__19202\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\
        );

    \I__1837\ : InMux
    port map (
            O => \N__19199\,
            I => \N__19196\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__19196\,
            I => \N__19193\
        );

    \I__1835\ : Span4Mux_v
    port map (
            O => \N__19193\,
            I => \N__19190\
        );

    \I__1834\ : Odrv4
    port map (
            O => \N__19190\,
            I => \pwm_generator_inst.un2_threshold_acc_1_17\
        );

    \I__1833\ : CascadeMux
    port map (
            O => \N__19187\,
            I => \N__19184\
        );

    \I__1832\ : InMux
    port map (
            O => \N__19184\,
            I => \N__19181\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__19181\,
            I => \N__19178\
        );

    \I__1830\ : Span4Mux_h
    port map (
            O => \N__19178\,
            I => \N__19175\
        );

    \I__1829\ : Odrv4
    port map (
            O => \N__19175\,
            I => \pwm_generator_inst.un2_threshold_acc_2_2\
        );

    \I__1828\ : InMux
    port map (
            O => \N__19172\,
            I => \N__19169\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__19169\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0\
        );

    \I__1826\ : InMux
    port map (
            O => \N__19166\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\
        );

    \I__1825\ : InMux
    port map (
            O => \N__19163\,
            I => \N__19160\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__19160\,
            I => \N__19157\
        );

    \I__1823\ : Span4Mux_s3_h
    port map (
            O => \N__19157\,
            I => \N__19154\
        );

    \I__1822\ : Span4Mux_v
    port map (
            O => \N__19154\,
            I => \N__19151\
        );

    \I__1821\ : Odrv4
    port map (
            O => \N__19151\,
            I => \pwm_generator_inst.un2_threshold_acc_1_18\
        );

    \I__1820\ : CascadeMux
    port map (
            O => \N__19148\,
            I => \N__19145\
        );

    \I__1819\ : InMux
    port map (
            O => \N__19145\,
            I => \N__19142\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__19142\,
            I => \N__19139\
        );

    \I__1817\ : Span4Mux_h
    port map (
            O => \N__19139\,
            I => \N__19136\
        );

    \I__1816\ : Odrv4
    port map (
            O => \N__19136\,
            I => \pwm_generator_inst.un2_threshold_acc_2_3\
        );

    \I__1815\ : InMux
    port map (
            O => \N__19133\,
            I => \N__19130\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__19130\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0\
        );

    \I__1813\ : InMux
    port map (
            O => \N__19127\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\
        );

    \I__1812\ : InMux
    port map (
            O => \N__19124\,
            I => \N__19121\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__19121\,
            I => \N__19118\
        );

    \I__1810\ : Span4Mux_v
    port map (
            O => \N__19118\,
            I => \N__19115\
        );

    \I__1809\ : Odrv4
    port map (
            O => \N__19115\,
            I => \pwm_generator_inst.un2_threshold_acc_1_19\
        );

    \I__1808\ : CascadeMux
    port map (
            O => \N__19112\,
            I => \N__19109\
        );

    \I__1807\ : InMux
    port map (
            O => \N__19109\,
            I => \N__19106\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__19106\,
            I => \N__19103\
        );

    \I__1805\ : Span4Mux_v
    port map (
            O => \N__19103\,
            I => \N__19100\
        );

    \I__1804\ : Odrv4
    port map (
            O => \N__19100\,
            I => \pwm_generator_inst.un2_threshold_acc_2_4\
        );

    \I__1803\ : InMux
    port map (
            O => \N__19097\,
            I => \N__19094\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__19094\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0\
        );

    \I__1801\ : InMux
    port map (
            O => \N__19091\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\
        );

    \I__1800\ : InMux
    port map (
            O => \N__19088\,
            I => \N__19085\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__19085\,
            I => \N__19082\
        );

    \I__1798\ : Span4Mux_v
    port map (
            O => \N__19082\,
            I => \N__19079\
        );

    \I__1797\ : Odrv4
    port map (
            O => \N__19079\,
            I => \pwm_generator_inst.un2_threshold_acc_1_20\
        );

    \I__1796\ : CascadeMux
    port map (
            O => \N__19076\,
            I => \N__19073\
        );

    \I__1795\ : InMux
    port map (
            O => \N__19073\,
            I => \N__19070\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__19070\,
            I => \N__19067\
        );

    \I__1793\ : Span4Mux_v
    port map (
            O => \N__19067\,
            I => \N__19064\
        );

    \I__1792\ : Odrv4
    port map (
            O => \N__19064\,
            I => \pwm_generator_inst.un2_threshold_acc_2_5\
        );

    \I__1791\ : InMux
    port map (
            O => \N__19061\,
            I => \N__19058\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__19058\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0\
        );

    \I__1789\ : InMux
    port map (
            O => \N__19055\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\
        );

    \I__1788\ : InMux
    port map (
            O => \N__19052\,
            I => \N__19049\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__19049\,
            I => \N__19046\
        );

    \I__1786\ : Span4Mux_v
    port map (
            O => \N__19046\,
            I => \N__19043\
        );

    \I__1785\ : Odrv4
    port map (
            O => \N__19043\,
            I => \pwm_generator_inst.un2_threshold_acc_1_21\
        );

    \I__1784\ : CascadeMux
    port map (
            O => \N__19040\,
            I => \N__19037\
        );

    \I__1783\ : InMux
    port map (
            O => \N__19037\,
            I => \N__19034\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__19034\,
            I => \N__19031\
        );

    \I__1781\ : Span4Mux_h
    port map (
            O => \N__19031\,
            I => \N__19028\
        );

    \I__1780\ : Odrv4
    port map (
            O => \N__19028\,
            I => \pwm_generator_inst.un2_threshold_acc_2_6\
        );

    \I__1779\ : InMux
    port map (
            O => \N__19025\,
            I => \N__19022\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__19022\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0\
        );

    \I__1777\ : InMux
    port map (
            O => \N__19019\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\
        );

    \I__1776\ : InMux
    port map (
            O => \N__19016\,
            I => \N__19010\
        );

    \I__1775\ : InMux
    port map (
            O => \N__19015\,
            I => \N__19010\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__19010\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\
        );

    \I__1773\ : InMux
    port map (
            O => \N__19007\,
            I => \N__19004\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__19004\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO\
        );

    \I__1771\ : CascadeMux
    port map (
            O => \N__19001\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_15_cascade_\
        );

    \I__1770\ : InMux
    port map (
            O => \N__18998\,
            I => \N__18994\
        );

    \I__1769\ : InMux
    port map (
            O => \N__18997\,
            I => \N__18991\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__18994\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_16\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__18991\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_16\
        );

    \I__1766\ : InMux
    port map (
            O => \N__18986\,
            I => \N__18980\
        );

    \I__1765\ : InMux
    port map (
            O => \N__18985\,
            I => \N__18980\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__18980\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\
        );

    \I__1763\ : InMux
    port map (
            O => \N__18977\,
            I => \N__18974\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__18974\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO\
        );

    \I__1761\ : CascadeMux
    port map (
            O => \N__18971\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_16_cascade_\
        );

    \I__1760\ : CascadeMux
    port map (
            O => \N__18968\,
            I => \N__18964\
        );

    \I__1759\ : InMux
    port map (
            O => \N__18967\,
            I => \N__18961\
        );

    \I__1758\ : InMux
    port map (
            O => \N__18964\,
            I => \N__18958\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__18961\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_17\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__18958\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_17\
        );

    \I__1755\ : InMux
    port map (
            O => \N__18953\,
            I => \N__18947\
        );

    \I__1754\ : InMux
    port map (
            O => \N__18952\,
            I => \N__18947\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__18947\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\
        );

    \I__1752\ : InMux
    port map (
            O => \N__18944\,
            I => \N__18941\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__18941\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO\
        );

    \I__1750\ : CascadeMux
    port map (
            O => \N__18938\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_\
        );

    \I__1749\ : InMux
    port map (
            O => \N__18935\,
            I => \N__18932\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__18932\,
            I => \N__18928\
        );

    \I__1747\ : InMux
    port map (
            O => \N__18931\,
            I => \N__18925\
        );

    \I__1746\ : Odrv4
    port map (
            O => \N__18928\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__18925\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\
        );

    \I__1744\ : CascadeMux
    port map (
            O => \N__18920\,
            I => \N__18917\
        );

    \I__1743\ : InMux
    port map (
            O => \N__18917\,
            I => \N__18914\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__18914\,
            I => \N__18911\
        );

    \I__1741\ : Span4Mux_h
    port map (
            O => \N__18911\,
            I => \N__18906\
        );

    \I__1740\ : InMux
    port map (
            O => \N__18910\,
            I => \N__18901\
        );

    \I__1739\ : InMux
    port map (
            O => \N__18909\,
            I => \N__18901\
        );

    \I__1738\ : Odrv4
    port map (
            O => \N__18906\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_18\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__18901\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_18\
        );

    \I__1736\ : InMux
    port map (
            O => \N__18896\,
            I => \N__18893\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__18893\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO\
        );

    \I__1734\ : CascadeMux
    port map (
            O => \N__18890\,
            I => \N__18886\
        );

    \I__1733\ : InMux
    port map (
            O => \N__18889\,
            I => \N__18883\
        );

    \I__1732\ : InMux
    port map (
            O => \N__18886\,
            I => \N__18880\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__18883\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_10\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__18880\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_10\
        );

    \I__1729\ : InMux
    port map (
            O => \N__18875\,
            I => \N__18872\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__18872\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO\
        );

    \I__1727\ : InMux
    port map (
            O => \N__18869\,
            I => \N__18863\
        );

    \I__1726\ : InMux
    port map (
            O => \N__18868\,
            I => \N__18863\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__18863\,
            I => \N__18860\
        );

    \I__1724\ : Span4Mux_v
    port map (
            O => \N__18860\,
            I => \N__18857\
        );

    \I__1723\ : Odrv4
    port map (
            O => \N__18857\,
            I => \pwm_generator_inst.O_10\
        );

    \I__1722\ : CascadeMux
    port map (
            O => \N__18854\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_10_cascade_\
        );

    \I__1721\ : InMux
    port map (
            O => \N__18851\,
            I => \N__18847\
        );

    \I__1720\ : InMux
    port map (
            O => \N__18850\,
            I => \N__18844\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__18847\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__18844\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\
        );

    \I__1717\ : InMux
    port map (
            O => \N__18839\,
            I => \N__18834\
        );

    \I__1716\ : InMux
    port map (
            O => \N__18838\,
            I => \N__18831\
        );

    \I__1715\ : InMux
    port map (
            O => \N__18837\,
            I => \N__18828\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__18834\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_14\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__18831\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_14\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__18828\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_14\
        );

    \I__1711\ : CascadeMux
    port map (
            O => \N__18821\,
            I => \N__18818\
        );

    \I__1710\ : InMux
    port map (
            O => \N__18818\,
            I => \N__18815\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__18815\,
            I => \N__18812\
        );

    \I__1708\ : Odrv4
    port map (
            O => \N__18812\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO\
        );

    \I__1707\ : CascadeMux
    port map (
            O => \N__18809\,
            I => \N__18805\
        );

    \I__1706\ : InMux
    port map (
            O => \N__18808\,
            I => \N__18802\
        );

    \I__1705\ : InMux
    port map (
            O => \N__18805\,
            I => \N__18799\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__18802\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_15\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__18799\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_15\
        );

    \I__1702\ : CascadeMux
    port map (
            O => \N__18794\,
            I => \N__18791\
        );

    \I__1701\ : InMux
    port map (
            O => \N__18791\,
            I => \N__18785\
        );

    \I__1700\ : InMux
    port map (
            O => \N__18790\,
            I => \N__18785\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__18785\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\
        );

    \I__1698\ : CascadeMux
    port map (
            O => \N__18782\,
            I => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_\
        );

    \I__1697\ : InMux
    port map (
            O => \N__18779\,
            I => \N__18776\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__18776\,
            I => \N__18771\
        );

    \I__1695\ : InMux
    port map (
            O => \N__18775\,
            I => \N__18766\
        );

    \I__1694\ : InMux
    port map (
            O => \N__18774\,
            I => \N__18766\
        );

    \I__1693\ : Span4Mux_s1_h
    port map (
            O => \N__18771\,
            I => \N__18763\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__18766\,
            I => pwm_duty_input_7
        );

    \I__1691\ : Odrv4
    port map (
            O => \N__18763\,
            I => pwm_duty_input_7
        );

    \I__1690\ : InMux
    port map (
            O => \N__18758\,
            I => \N__18753\
        );

    \I__1689\ : InMux
    port map (
            O => \N__18757\,
            I => \N__18748\
        );

    \I__1688\ : InMux
    port map (
            O => \N__18756\,
            I => \N__18748\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__18753\,
            I => \N__18745\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__18748\,
            I => pwm_duty_input_5
        );

    \I__1685\ : Odrv4
    port map (
            O => \N__18745\,
            I => pwm_duty_input_5
        );

    \I__1684\ : InMux
    port map (
            O => \N__18740\,
            I => \N__18736\
        );

    \I__1683\ : CascadeMux
    port map (
            O => \N__18739\,
            I => \N__18733\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__18736\,
            I => \N__18729\
        );

    \I__1681\ : InMux
    port map (
            O => \N__18733\,
            I => \N__18724\
        );

    \I__1680\ : InMux
    port map (
            O => \N__18732\,
            I => \N__18724\
        );

    \I__1679\ : Span4Mux_s2_h
    port map (
            O => \N__18729\,
            I => \N__18721\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__18724\,
            I => pwm_duty_input_8
        );

    \I__1677\ : Odrv4
    port map (
            O => \N__18721\,
            I => pwm_duty_input_8
        );

    \I__1676\ : InMux
    port map (
            O => \N__18716\,
            I => \N__18713\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__18713\,
            I => \N__18708\
        );

    \I__1674\ : InMux
    port map (
            O => \N__18712\,
            I => \N__18703\
        );

    \I__1673\ : InMux
    port map (
            O => \N__18711\,
            I => \N__18703\
        );

    \I__1672\ : Span4Mux_s2_h
    port map (
            O => \N__18708\,
            I => \N__18700\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__18703\,
            I => pwm_duty_input_9
        );

    \I__1670\ : Odrv4
    port map (
            O => \N__18700\,
            I => pwm_duty_input_9
        );

    \I__1669\ : CascadeMux
    port map (
            O => \N__18695\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\
        );

    \I__1668\ : InMux
    port map (
            O => \N__18692\,
            I => \N__18687\
        );

    \I__1667\ : InMux
    port map (
            O => \N__18691\,
            I => \N__18682\
        );

    \I__1666\ : InMux
    port map (
            O => \N__18690\,
            I => \N__18682\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__18687\,
            I => \N__18679\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__18682\,
            I => \N__18676\
        );

    \I__1663\ : Span4Mux_s1_h
    port map (
            O => \N__18679\,
            I => \N__18673\
        );

    \I__1662\ : Odrv4
    port map (
            O => \N__18676\,
            I => pwm_duty_input_6
        );

    \I__1661\ : Odrv4
    port map (
            O => \N__18673\,
            I => pwm_duty_input_6
        );

    \I__1660\ : InMux
    port map (
            O => \N__18668\,
            I => \N__18659\
        );

    \I__1659\ : InMux
    port map (
            O => \N__18667\,
            I => \N__18659\
        );

    \I__1658\ : InMux
    port map (
            O => \N__18666\,
            I => \N__18659\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__18659\,
            I => \current_shift_inst.PI_CTRL.N_97\
        );

    \I__1656\ : InMux
    port map (
            O => \N__18656\,
            I => \N__18652\
        );

    \I__1655\ : InMux
    port map (
            O => \N__18655\,
            I => \N__18649\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__18652\,
            I => pwm_duty_input_0
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__18649\,
            I => pwm_duty_input_0
        );

    \I__1652\ : InMux
    port map (
            O => \N__18644\,
            I => \N__18640\
        );

    \I__1651\ : InMux
    port map (
            O => \N__18643\,
            I => \N__18637\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__18640\,
            I => pwm_duty_input_2
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__18637\,
            I => pwm_duty_input_2
        );

    \I__1648\ : InMux
    port map (
            O => \N__18632\,
            I => \N__18628\
        );

    \I__1647\ : InMux
    port map (
            O => \N__18631\,
            I => \N__18625\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__18628\,
            I => pwm_duty_input_1
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__18625\,
            I => pwm_duty_input_1
        );

    \I__1644\ : InMux
    port map (
            O => \N__18620\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_19\
        );

    \I__1643\ : InMux
    port map (
            O => \N__18617\,
            I => \N__18614\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__18614\,
            I => \N__18610\
        );

    \I__1641\ : InMux
    port map (
            O => \N__18613\,
            I => \N__18607\
        );

    \I__1640\ : Odrv4
    port map (
            O => \N__18610\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1_15\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__18607\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1_15\
        );

    \I__1638\ : CascadeMux
    port map (
            O => \N__18602\,
            I => \N__18599\
        );

    \I__1637\ : InMux
    port map (
            O => \N__18599\,
            I => \N__18596\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__18596\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1_16\
        );

    \I__1635\ : InMux
    port map (
            O => \N__18593\,
            I => \N__18590\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__18590\,
            I => un7_start_stop_0_a3
        );

    \I__1633\ : InMux
    port map (
            O => \N__18587\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_6\
        );

    \I__1632\ : InMux
    port map (
            O => \N__18584\,
            I => \bfn_1_11_0_\
        );

    \I__1631\ : InMux
    port map (
            O => \N__18581\,
            I => \N__18577\
        );

    \I__1630\ : InMux
    port map (
            O => \N__18580\,
            I => \N__18574\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__18577\,
            I => \N__18569\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__18574\,
            I => \N__18569\
        );

    \I__1627\ : Span4Mux_v
    port map (
            O => \N__18569\,
            I => \N__18566\
        );

    \I__1626\ : Odrv4
    port map (
            O => \N__18566\,
            I => \pwm_generator_inst.un3_threshold_acc\
        );

    \I__1625\ : InMux
    port map (
            O => \N__18563\,
            I => \N__18560\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__18560\,
            I => \N__18557\
        );

    \I__1623\ : Span4Mux_v
    port map (
            O => \N__18557\,
            I => \N__18554\
        );

    \I__1622\ : Odrv4
    port map (
            O => \N__18554\,
            I => \pwm_generator_inst.O_12\
        );

    \I__1621\ : InMux
    port map (
            O => \N__18551\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_0\
        );

    \I__1620\ : InMux
    port map (
            O => \N__18548\,
            I => \N__18545\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__18545\,
            I => \N__18542\
        );

    \I__1618\ : Span4Mux_v
    port map (
            O => \N__18542\,
            I => \N__18539\
        );

    \I__1617\ : Odrv4
    port map (
            O => \N__18539\,
            I => \pwm_generator_inst.O_13\
        );

    \I__1616\ : InMux
    port map (
            O => \N__18536\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_1\
        );

    \I__1615\ : InMux
    port map (
            O => \N__18533\,
            I => \N__18530\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__18530\,
            I => \N__18527\
        );

    \I__1613\ : Span4Mux_v
    port map (
            O => \N__18527\,
            I => \N__18524\
        );

    \I__1612\ : Odrv4
    port map (
            O => \N__18524\,
            I => \pwm_generator_inst.O_14\
        );

    \I__1611\ : InMux
    port map (
            O => \N__18521\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_2\
        );

    \I__1610\ : InMux
    port map (
            O => \N__18518\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_3\
        );

    \I__1609\ : InMux
    port map (
            O => \N__18515\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_4\
        );

    \I__1608\ : InMux
    port map (
            O => \N__18512\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_5\
        );

    \I__1607\ : InMux
    port map (
            O => \N__18509\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_10\
        );

    \I__1606\ : InMux
    port map (
            O => \N__18506\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_11\
        );

    \I__1605\ : InMux
    port map (
            O => \N__18503\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_12\
        );

    \I__1604\ : InMux
    port map (
            O => \N__18500\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_13\
        );

    \I__1603\ : InMux
    port map (
            O => \N__18497\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_14\
        );

    \I__1602\ : InMux
    port map (
            O => \N__18494\,
            I => \bfn_1_9_0_\
        );

    \I__1601\ : InMux
    port map (
            O => \N__18491\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_16\
        );

    \I__1600\ : InMux
    port map (
            O => \N__18488\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_17\
        );

    \I__1599\ : InMux
    port map (
            O => \N__18485\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_18\
        );

    \I__1598\ : InMux
    port map (
            O => \N__18482\,
            I => \N__18479\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__18479\,
            I => \N__18476\
        );

    \I__1596\ : Odrv4
    port map (
            O => \N__18476\,
            I => \pwm_generator_inst.O_3\
        );

    \I__1595\ : InMux
    port map (
            O => \N__18473\,
            I => \N__18470\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__18470\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_3\
        );

    \I__1593\ : InMux
    port map (
            O => \N__18467\,
            I => \N__18464\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__18464\,
            I => \N__18461\
        );

    \I__1591\ : Span4Mux_h
    port map (
            O => \N__18461\,
            I => \N__18458\
        );

    \I__1590\ : Odrv4
    port map (
            O => \N__18458\,
            I => \pwm_generator_inst.O_4\
        );

    \I__1589\ : InMux
    port map (
            O => \N__18455\,
            I => \N__18452\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__18452\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_4\
        );

    \I__1587\ : InMux
    port map (
            O => \N__18449\,
            I => \N__18446\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__18446\,
            I => \N__18443\
        );

    \I__1585\ : Odrv4
    port map (
            O => \N__18443\,
            I => \pwm_generator_inst.O_5\
        );

    \I__1584\ : InMux
    port map (
            O => \N__18440\,
            I => \N__18437\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__18437\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_5\
        );

    \I__1582\ : InMux
    port map (
            O => \N__18434\,
            I => \N__18431\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__18431\,
            I => \N__18428\
        );

    \I__1580\ : Span4Mux_h
    port map (
            O => \N__18428\,
            I => \N__18425\
        );

    \I__1579\ : Odrv4
    port map (
            O => \N__18425\,
            I => \pwm_generator_inst.O_6\
        );

    \I__1578\ : InMux
    port map (
            O => \N__18422\,
            I => \N__18419\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__18419\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_6\
        );

    \I__1576\ : InMux
    port map (
            O => \N__18416\,
            I => \N__18413\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__18413\,
            I => \N__18410\
        );

    \I__1574\ : Span4Mux_v
    port map (
            O => \N__18410\,
            I => \N__18407\
        );

    \I__1573\ : Odrv4
    port map (
            O => \N__18407\,
            I => \pwm_generator_inst.O_7\
        );

    \I__1572\ : InMux
    port map (
            O => \N__18404\,
            I => \N__18401\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__18401\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_7\
        );

    \I__1570\ : InMux
    port map (
            O => \N__18398\,
            I => \N__18395\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__18395\,
            I => \N__18392\
        );

    \I__1568\ : Odrv4
    port map (
            O => \N__18392\,
            I => \pwm_generator_inst.O_8\
        );

    \I__1567\ : InMux
    port map (
            O => \N__18389\,
            I => \N__18386\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__18386\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_8\
        );

    \I__1565\ : InMux
    port map (
            O => \N__18383\,
            I => \N__18380\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__18380\,
            I => \N__18377\
        );

    \I__1563\ : Odrv4
    port map (
            O => \N__18377\,
            I => \pwm_generator_inst.O_9\
        );

    \I__1562\ : CascadeMux
    port map (
            O => \N__18374\,
            I => \N__18371\
        );

    \I__1561\ : InMux
    port map (
            O => \N__18371\,
            I => \N__18368\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__18368\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_9\
        );

    \I__1559\ : InMux
    port map (
            O => \N__18365\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_9\
        );

    \I__1558\ : InMux
    port map (
            O => \N__18362\,
            I => \N__18359\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__18359\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__1556\ : CascadeMux
    port map (
            O => \N__18356\,
            I => \current_shift_inst.PI_CTRL.N_96_cascade_\
        );

    \I__1555\ : CascadeMux
    port map (
            O => \N__18353\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_3_cascade_\
        );

    \I__1554\ : InMux
    port map (
            O => \N__18350\,
            I => \N__18344\
        );

    \I__1553\ : InMux
    port map (
            O => \N__18349\,
            I => \N__18344\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__18344\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_3\
        );

    \I__1551\ : InMux
    port map (
            O => \N__18341\,
            I => \N__18329\
        );

    \I__1550\ : InMux
    port map (
            O => \N__18340\,
            I => \N__18329\
        );

    \I__1549\ : InMux
    port map (
            O => \N__18339\,
            I => \N__18329\
        );

    \I__1548\ : InMux
    port map (
            O => \N__18338\,
            I => \N__18329\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__18329\,
            I => \current_shift_inst.PI_CTRL.N_96\
        );

    \I__1546\ : InMux
    port map (
            O => \N__18326\,
            I => \N__18323\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__18323\,
            I => \N__18320\
        );

    \I__1544\ : Odrv4
    port map (
            O => \N__18320\,
            I => \pwm_generator_inst.O_0\
        );

    \I__1543\ : InMux
    port map (
            O => \N__18317\,
            I => \N__18314\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__18314\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_0\
        );

    \I__1541\ : InMux
    port map (
            O => \N__18311\,
            I => \N__18308\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__18308\,
            I => \N__18305\
        );

    \I__1539\ : Span4Mux_v
    port map (
            O => \N__18305\,
            I => \N__18302\
        );

    \I__1538\ : Odrv4
    port map (
            O => \N__18302\,
            I => \pwm_generator_inst.O_1\
        );

    \I__1537\ : InMux
    port map (
            O => \N__18299\,
            I => \N__18296\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__18296\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_1\
        );

    \I__1535\ : InMux
    port map (
            O => \N__18293\,
            I => \N__18290\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__18290\,
            I => \N__18287\
        );

    \I__1533\ : Odrv4
    port map (
            O => \N__18287\,
            I => \pwm_generator_inst.O_2\
        );

    \I__1532\ : InMux
    port map (
            O => \N__18284\,
            I => \N__18281\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__18281\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_2\
        );

    \I__1530\ : CascadeMux
    port map (
            O => \N__18278\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_\
        );

    \I__1529\ : CascadeMux
    port map (
            O => \N__18275\,
            I => \current_shift_inst.PI_CTRL.N_27_cascade_\
        );

    \IN_MUX_bfv_9_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_13_0_\
        );

    \IN_MUX_bfv_9_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_0_cry_6\,
            carryinitout => \bfn_9_14_0_\
        );

    \IN_MUX_bfv_9_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_0_cry_14\,
            carryinitout => \bfn_9_15_0_\
        );

    \IN_MUX_bfv_9_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_0_cry_22\,
            carryinitout => \bfn_9_16_0_\
        );

    \IN_MUX_bfv_9_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_0_cry_30\,
            carryinitout => \bfn_9_17_0_\
        );

    \IN_MUX_bfv_4_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_5_0_\
        );

    \IN_MUX_bfv_4_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un5_counter_cry_8,
            carryinitout => \bfn_4_6_0_\
        );

    \IN_MUX_bfv_1_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_10_0_\
        );

    \IN_MUX_bfv_1_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_acc_cry_7\,
            carryinitout => \bfn_1_11_0_\
        );

    \IN_MUX_bfv_1_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_acc_cry_15\,
            carryinitout => \bfn_1_12_0_\
        );

    \IN_MUX_bfv_14_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_18_0_\
        );

    \IN_MUX_bfv_14_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_14_19_0_\
        );

    \IN_MUX_bfv_14_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_14_20_0_\
        );

    \IN_MUX_bfv_15_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_16_0_\
        );

    \IN_MUX_bfv_15_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_15_17_0_\
        );

    \IN_MUX_bfv_15_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_15_18_0_\
        );

    \IN_MUX_bfv_18_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_19_0_\
        );

    \IN_MUX_bfv_18_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_18_20_0_\
        );

    \IN_MUX_bfv_18_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_18_21_0_\
        );

    \IN_MUX_bfv_13_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_24_0_\
        );

    \IN_MUX_bfv_13_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_13_25_0_\
        );

    \IN_MUX_bfv_13_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_13_26_0_\
        );

    \IN_MUX_bfv_13_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_13_0_\
        );

    \IN_MUX_bfv_13_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_13_14_0_\
        );

    \IN_MUX_bfv_13_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_13_15_0_\
        );

    \IN_MUX_bfv_15_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_13_0_\
        );

    \IN_MUX_bfv_15_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_15_14_0_\
        );

    \IN_MUX_bfv_15_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_15_15_0_\
        );

    \IN_MUX_bfv_8_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_17_0_\
        );

    \IN_MUX_bfv_8_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.z_5_cry_8\,
            carryinitout => \bfn_8_18_0_\
        );

    \IN_MUX_bfv_8_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.z_5_cry_16\,
            carryinitout => \bfn_8_19_0_\
        );

    \IN_MUX_bfv_8_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.z_5_cry_24\,
            carryinitout => \bfn_8_20_0_\
        );

    \IN_MUX_bfv_2_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_11_0_\
        );

    \IN_MUX_bfv_2_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7\,
            carryinitout => \bfn_2_12_0_\
        );

    \IN_MUX_bfv_2_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15\,
            carryinitout => \bfn_2_13_0_\
        );

    \IN_MUX_bfv_1_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_7_0_\
        );

    \IN_MUX_bfv_1_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_acc_1_cry_7\,
            carryinitout => \bfn_1_8_0_\
        );

    \IN_MUX_bfv_1_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_acc_1_cry_15\,
            carryinitout => \bfn_1_9_0_\
        );

    \IN_MUX_bfv_8_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_8_0_\
        );

    \IN_MUX_bfv_8_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un14_counter_cry_7\,
            carryinitout => \bfn_8_9_0_\
        );

    \IN_MUX_bfv_3_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_8_0_\
        );

    \IN_MUX_bfv_3_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un19_threshold_acc_cry_7\,
            carryinitout => \bfn_3_9_0_\
        );

    \IN_MUX_bfv_9_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_7_0_\
        );

    \IN_MUX_bfv_9_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.counter_cry_7\,
            carryinitout => \bfn_9_8_0_\
        );

    \IN_MUX_bfv_15_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_21_0_\
        );

    \IN_MUX_bfv_15_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8\,
            carryinitout => \bfn_15_22_0_\
        );

    \IN_MUX_bfv_15_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16\,
            carryinitout => \bfn_15_23_0_\
        );

    \IN_MUX_bfv_15_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_24_0_\
        );

    \IN_MUX_bfv_15_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            carryinitout => \bfn_15_25_0_\
        );

    \IN_MUX_bfv_15_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            carryinitout => \bfn_15_26_0_\
        );

    \IN_MUX_bfv_18_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_15_0_\
        );

    \IN_MUX_bfv_18_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_18_16_0_\
        );

    \IN_MUX_bfv_18_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_18_17_0_\
        );

    \IN_MUX_bfv_18_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_18_18_0_\
        );

    \IN_MUX_bfv_17_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_13_0_\
        );

    \IN_MUX_bfv_17_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            carryinitout => \bfn_17_14_0_\
        );

    \IN_MUX_bfv_17_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            carryinitout => \bfn_17_15_0_\
        );

    \IN_MUX_bfv_17_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            carryinitout => \bfn_17_16_0_\
        );

    \IN_MUX_bfv_17_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_8_0_\
        );

    \IN_MUX_bfv_17_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_17_9_0_\
        );

    \IN_MUX_bfv_17_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_17_10_0_\
        );

    \IN_MUX_bfv_17_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_17_11_0_\
        );

    \IN_MUX_bfv_16_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_7_0_\
        );

    \IN_MUX_bfv_16_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            carryinitout => \bfn_16_8_0_\
        );

    \IN_MUX_bfv_16_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            carryinitout => \bfn_16_9_0_\
        );

    \IN_MUX_bfv_16_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            carryinitout => \bfn_16_10_0_\
        );

    \IN_MUX_bfv_9_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_18_0_\
        );

    \IN_MUX_bfv_9_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.z_cry_7\,
            carryinitout => \bfn_9_19_0_\
        );

    \IN_MUX_bfv_9_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.z_cry_15\,
            carryinitout => \bfn_9_20_0_\
        );

    \IN_MUX_bfv_9_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.z_cry_23\,
            carryinitout => \bfn_9_21_0_\
        );

    \IN_MUX_bfv_10_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_17_0_\
        );

    \IN_MUX_bfv_10_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_cry_8\,
            carryinitout => \bfn_10_18_0_\
        );

    \IN_MUX_bfv_10_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_cry_16\,
            carryinitout => \bfn_10_19_0_\
        );

    \IN_MUX_bfv_10_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_cry_24\,
            carryinitout => \bfn_10_20_0_\
        );

    \IN_MUX_bfv_12_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_19_0_\
        );

    \IN_MUX_bfv_12_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_12_20_0_\
        );

    \IN_MUX_bfv_12_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_12_21_0_\
        );

    \IN_MUX_bfv_12_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_12_22_0_\
        );

    \IN_MUX_bfv_10_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_21_0_\
        );

    \IN_MUX_bfv_10_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_7\,
            carryinitout => \bfn_10_22_0_\
        );

    \IN_MUX_bfv_10_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_15\,
            carryinitout => \bfn_10_23_0_\
        );

    \IN_MUX_bfv_10_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_23\,
            carryinitout => \bfn_10_24_0_\
        );

    \IN_MUX_bfv_7_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_19_0_\
        );

    \IN_MUX_bfv_7_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_7_20_0_\
        );

    \IN_MUX_bfv_7_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_7_21_0_\
        );

    \IN_MUX_bfv_7_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_7_22_0_\
        );

    \IN_MUX_bfv_8_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_21_0_\
        );

    \IN_MUX_bfv_8_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_phase.counter_cry_7\,
            carryinitout => \bfn_8_22_0_\
        );

    \IN_MUX_bfv_8_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_phase.counter_cry_15\,
            carryinitout => \bfn_8_23_0_\
        );

    \IN_MUX_bfv_8_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_phase.counter_cry_23\,
            carryinitout => \bfn_8_24_0_\
        );

    \IN_MUX_bfv_8_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_13_0_\
        );

    \IN_MUX_bfv_8_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_1_cry_7\,
            carryinitout => \bfn_8_14_0_\
        );

    \IN_MUX_bfv_8_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_1_cry_15\,
            carryinitout => \bfn_8_15_0_\
        );

    \IN_MUX_bfv_8_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_1_cry_23\,
            carryinitout => \bfn_8_16_0_\
        );

    \IN_MUX_bfv_5_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_9_0_\
        );

    \IN_MUX_bfv_5_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            carryinitout => \bfn_5_10_0_\
        );

    \IN_MUX_bfv_5_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            carryinitout => \bfn_5_11_0_\
        );

    \IN_MUX_bfv_5_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            carryinitout => \bfn_5_12_0_\
        );

    \IN_MUX_bfv_11_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_10_0_\
        );

    \IN_MUX_bfv_11_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\,
            carryinitout => \bfn_11_11_0_\
        );

    \IN_MUX_bfv_11_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\,
            carryinitout => \bfn_11_12_0_\
        );

    \IN_MUX_bfv_11_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\,
            carryinitout => \bfn_11_13_0_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__34067\,
            GLOBALBUFFEROUTPUT => \delay_measurement_inst.delay_hc_timer.N_335_i_g\
        );

    \current_shift_inst.timer_s1.running_RNII51H_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__24020\,
            GLOBALBUFFEROUTPUT => \current_shift_inst.timer_s1.N_187_i_g\
        );

    \current_shift_inst.timer_phase.running_RNIC90O_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__27425\,
            GLOBALBUFFEROUTPUT => \current_shift_inst.timer_phase.N_188_i_g\
        );

    \osc\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b10"
        )
    port map (
            CLKHFPU => \N__22857\,
            CLKHFEN => \N__22859\,
            CLKHF => clk_12mhz
        );

    \rgb_drv\ : SB_RGBA_DRV
    generic map (
            RGB2_CURRENT => "0b111111",
            CURRENT_MODE => "0b0",
            RGB0_CURRENT => "0b111111",
            RGB1_CURRENT => "0b111111"
        )
    port map (
            RGBLEDEN => \N__22858\,
            RGB2PWM => \N__19601\,
            RGB1 => rgb_g_wire,
            CURREN => \N__22993\,
            RGB2 => rgb_b_wire,
            RGB1PWM => \N__18593\,
            RGB0PWM => \N__47463\,
            RGB0 => rgb_r_wire
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_6_LC_1_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000001110"
        )
    port map (
            in0 => \N__21323\,
            in1 => \N__19892\,
            in2 => \N__21896\,
            in3 => \N__19829\,
            lcout => pwm_duty_input_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48008\,
            ce => \N__32559\,
            sr => \N__47350\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21208\,
            in2 => \_gnd_net_\,
            in3 => \N__21349\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21247\,
            in1 => \N__21286\,
            in2 => \N__18278\,
            in3 => \N__21322\,
            lcout => \current_shift_inst.PI_CTRL.N_27\,
            ltout => \current_shift_inst.PI_CTRL.N_27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_4_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011011111"
        )
    port map (
            in0 => \N__19828\,
            in1 => \N__20870\,
            in2 => \N__18275\,
            in3 => \N__19589\,
            lcout => pwm_duty_input_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48007\,
            ce => \N__32560\,
            sr => \N__47357\
        );

    \current_shift_inst.PI_CTRL.control_out_5_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000001110"
        )
    port map (
            in0 => \N__21350\,
            in1 => \N__19890\,
            in2 => \N__21893\,
            in3 => \N__19826\,
            lcout => pwm_duty_input_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48007\,
            ce => \N__32560\,
            sr => \N__47357\
        );

    \current_shift_inst.PI_CTRL.control_out_7_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000001110"
        )
    port map (
            in0 => \N__21287\,
            in1 => \N__19891\,
            in2 => \N__21894\,
            in3 => \N__19827\,
            lcout => pwm_duty_input_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48007\,
            ce => \N__32560\,
            sr => \N__47357\
        );

    \current_shift_inst.PI_CTRL.control_out_2_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__18668\,
            in1 => \N__18340\,
            in2 => \N__20930\,
            in3 => \N__18350\,
            lcout => pwm_duty_input_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48005\,
            ce => \N__32540\,
            sr => \N__47367\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__20990\,
            in1 => \N__18362\,
            in2 => \N__21895\,
            in3 => \N__19813\,
            lcout => \current_shift_inst.PI_CTRL.N_96\,
            ltout => \current_shift_inst.PI_CTRL.N_96_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100110000"
        )
    port map (
            in0 => \N__19886\,
            in1 => \N__20896\,
            in2 => \N__18356\,
            in3 => \N__18790\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_0_3\,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_1_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__18339\,
            in1 => \N__20945\,
            in2 => \N__18353\,
            in3 => \N__18667\,
            lcout => pwm_duty_input_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48005\,
            ce => \N__32540\,
            sr => \N__47367\
        );

    \current_shift_inst.PI_CTRL.control_out_0_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__18666\,
            in1 => \N__18338\,
            in2 => \N__20963\,
            in3 => \N__18349\,
            lcout => pwm_duty_input_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48005\,
            ce => \N__32540\,
            sr => \N__47367\
        );

    \current_shift_inst.PI_CTRL.control_out_3_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110111001101"
        )
    port map (
            in0 => \N__18341\,
            in1 => \N__20897\,
            in2 => \N__18794\,
            in3 => \N__19887\,
            lcout => pwm_duty_input_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48005\,
            ce => \N__32540\,
            sr => \N__47367\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__18326\,
            in1 => \N__18317\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_1_7_0_\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18299\,
            in2 => \_gnd_net_\,
            in3 => \N__18311\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_0\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18284\,
            in2 => \_gnd_net_\,
            in3 => \N__18293\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_1\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18473\,
            in2 => \_gnd_net_\,
            in3 => \N__18482\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_2\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18455\,
            in2 => \_gnd_net_\,
            in3 => \N__18467\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_3\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18440\,
            in2 => \_gnd_net_\,
            in3 => \N__18449\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_4\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18422\,
            in2 => \_gnd_net_\,
            in3 => \N__18434\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_5\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18404\,
            in2 => \_gnd_net_\,
            in3 => \N__18416\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_6\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__18398\,
            in1 => \N__18389\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_8\,
            ltout => OPEN,
            carryin => \bfn_1_8_0_\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18374\,
            in3 => \N__18383\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_8\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18890\,
            in3 => \N__18365\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_9\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__20030\,
            in1 => \N__18581\,
            in2 => \_gnd_net_\,
            in3 => \N__18509\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_10\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20098\,
            in2 => \_gnd_net_\,
            in3 => \N__18506\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_11\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20163\,
            in2 => \_gnd_net_\,
            in3 => \N__18503\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_12\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18837\,
            in2 => \_gnd_net_\,
            in3 => \N__18500\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_13\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18809\,
            in3 => \N__18497\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_14\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18997\,
            in2 => \_gnd_net_\,
            in3 => \N__18494\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_1_9_0_\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18968\,
            in3 => \N__18491\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_16\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18909\,
            in2 => \_gnd_net_\,
            in3 => \N__18488\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_17\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18485\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18839\,
            in2 => \_gnd_net_\,
            in3 => \N__18850\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__18910\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18931\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18580\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_10_0_\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18563\,
            in2 => \_gnd_net_\,
            in3 => \N__18551\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_0\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18548\,
            in2 => \_gnd_net_\,
            in3 => \N__18536\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_1\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18533\,
            in2 => \_gnd_net_\,
            in3 => \N__18521\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_2\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19244\,
            in2 => \_gnd_net_\,
            in3 => \N__18518\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_3\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22994\,
            in2 => \N__19211\,
            in3 => \N__18515\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_4\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19172\,
            in2 => \N__23055\,
            in3 => \N__18512\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_5\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19133\,
            in2 => \N__23056\,
            in3 => \N__18587\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_6\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19097\,
            in2 => \_gnd_net_\,
            in3 => \N__18584\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_1_11_0_\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19061\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_8\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19025\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_9\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19472\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_10\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19433\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_11\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19397\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_12\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19373\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_13\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19352\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_14\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19328\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_12_0_\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19307\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_16\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19283\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_17\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19625\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_18\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18620\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__18613\,
            in1 => \N__19672\,
            in2 => \_gnd_net_\,
            in3 => \N__20615\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001011010"
        )
    port map (
            in0 => \N__19676\,
            in1 => \N__18617\,
            in2 => \N__18602\,
            in3 => \N__20614\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un7_start_stop_0_a3_LC_1_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__47462\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33731\,
            lcout => un7_start_stop_0_a3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_8_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000001110"
        )
    port map (
            in0 => \N__21248\,
            in1 => \N__19888\,
            in2 => \N__21891\,
            in3 => \N__19814\,
            lcout => pwm_duty_input_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48006\,
            ce => \N__32548\,
            sr => \N__47351\
        );

    \current_shift_inst.PI_CTRL.control_out_9_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000001110"
        )
    port map (
            in0 => \N__21209\,
            in1 => \N__19889\,
            in2 => \N__21892\,
            in3 => \N__19815\,
            lcout => pwm_duty_input_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48006\,
            ce => \N__32548\,
            sr => \N__47351\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110011"
        )
    port map (
            in0 => \N__19575\,
            in1 => \N__21861\,
            in2 => \_gnd_net_\,
            in3 => \N__20859\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18775\,
            in1 => \N__18712\,
            in2 => \N__18739\,
            in3 => \N__18691\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__19555\,
            in1 => \N__19518\,
            in2 => \N__18782\,
            in3 => \N__18757\,
            lcout => \pwm_generator_inst.N_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18774\,
            in2 => \_gnd_net_\,
            in3 => \N__18756\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__18732\,
            in1 => \N__18711\,
            in2 => \N__18695\,
            in3 => \N__18690\,
            lcout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__19576\,
            in1 => \N__21862\,
            in2 => \_gnd_net_\,
            in3 => \N__19885\,
            lcout => \current_shift_inst.PI_CTRL.N_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un1_duty_inputlto2_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__18656\,
            in1 => \N__18644\,
            in2 => \_gnd_net_\,
            in3 => \N__18632\,
            lcout => \pwm_generator_inst.un1_duty_inputlt3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_2_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__20420\,
            in1 => \N__20360\,
            in2 => \N__20553\,
            in3 => \N__19730\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48003\,
            ce => 'H',
            sr => \N__47368\
        );

    \pwm_generator_inst.threshold_ACC_3_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__20421\,
            in1 => \N__20361\,
            in2 => \N__20554\,
            in3 => \N__19721\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48003\,
            ce => 'H',
            sr => \N__47368\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__18935\,
            in1 => \N__20032\,
            in2 => \N__18920\,
            in3 => \N__18896\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__18868\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18889\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_10\,
            ltout => \pwm_generator_inst.un15_threshold_acc_1_axb_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010111001100"
        )
    port map (
            in0 => \N__18875\,
            in1 => \N__18869\,
            in2 => \N__18854\,
            in3 => \N__20031\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_0_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__34990\,
            in1 => \N__35617\,
            in2 => \N__40553\,
            in3 => \N__39596\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48000\,
            ce => \N__33569\,
            sr => \N__47375\
        );

    \phase_controller_inst1.stoper_hc.target_time_9_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010000000101"
        )
    port map (
            in0 => \N__35616\,
            in1 => \N__36418\,
            in2 => \N__40559\,
            in3 => \N__34989\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48000\,
            ce => \N__33569\,
            sr => \N__47375\
        );

    \phase_controller_inst1.stoper_hc.target_time_10_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__34991\,
            in1 => \_gnd_net_\,
            in2 => \N__34691\,
            in3 => \N__40554\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48000\,
            ce => \N__33569\,
            sr => \N__47375\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__18851\,
            in1 => \N__18838\,
            in2 => \N__18821\,
            in3 => \N__20034\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__18808\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19015\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_15\,
            ltout => \pwm_generator_inst.un15_threshold_acc_1_axb_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__19016\,
            in1 => \N__19007\,
            in2 => \N__19001\,
            in3 => \N__20035\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18985\,
            in2 => \_gnd_net_\,
            in3 => \N__18998\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_16\,
            ltout => \pwm_generator_inst.un15_threshold_acc_1_axb_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__18986\,
            in1 => \N__18977\,
            in2 => \N__18971\,
            in3 => \N__20033\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18952\,
            in2 => \_gnd_net_\,
            in3 => \N__18967\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_17\,
            ltout => \pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__18953\,
            in1 => \N__18944\,
            in2 => \N__18938\,
            in3 => \N__20036\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20167\,
            in2 => \_gnd_net_\,
            in3 => \N__20140\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_8_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111010111110011"
        )
    port map (
            in0 => \N__20430\,
            in1 => \N__20401\,
            in2 => \N__19940\,
            in3 => \N__20597\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47996\,
            ce => 'H',
            sr => \N__47388\
        );

    \pwm_generator_inst.threshold_ACC_9_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011000000"
        )
    port map (
            in0 => \N__20431\,
            in1 => \N__20402\,
            in2 => \N__19901\,
            in3 => \N__20598\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47996\,
            ce => 'H',
            sr => \N__47388\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20068\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20097\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_axb_4_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19274\,
            in2 => \N__19262\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \bfn_2_11_0_\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19238\,
            in2 => \N__19226\,
            in3 => \N__19202\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19199\,
            in2 => \N__19187\,
            in3 => \N__19166\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19163\,
            in2 => \N__19148\,
            in3 => \N__19127\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19124\,
            in2 => \N__19112\,
            in3 => \N__19091\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19088\,
            in2 => \N__19076\,
            in3 => \N__19055\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19052\,
            in2 => \N__19040\,
            in3 => \N__19019\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19499\,
            in2 => \N__19487\,
            in3 => \N__19466\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19463\,
            in2 => \N__19448\,
            in3 => \N__19427\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0\,
            ltout => OPEN,
            carryin => \bfn_2_12_0_\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19424\,
            in2 => \N__19412\,
            in3 => \N__19391\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19657\,
            in2 => \N__19388\,
            in3 => \N__19367\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19364\,
            in2 => \N__19673\,
            in3 => \N__19346\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19661\,
            in2 => \N__19343\,
            in3 => \N__19322\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19319\,
            in2 => \N__19674\,
            in3 => \N__19301\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19665\,
            in2 => \N__19298\,
            in3 => \N__19277\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19682\,
            in2 => \N__19675\,
            in3 => \N__19619\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__19616\,
            in1 => \N__19610\,
            in2 => \_gnd_net_\,
            in3 => \N__19604\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.N_32_i_i_LC_2_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33730\,
            in2 => \_gnd_net_\,
            in3 => \N__47461\,
            lcout => \N_32_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_3_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000111"
        )
    port map (
            in0 => \N__20866\,
            in1 => \N__19577\,
            in2 => \N__21890\,
            in3 => \N__19863\,
            lcout => \current_shift_inst.PI_CTRL.N_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_0_5_LC_3_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21201\,
            in2 => \_gnd_net_\,
            in3 => \N__21343\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_3_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__21240\,
            in1 => \N__21279\,
            in2 => \N__19580\,
            in3 => \N__21315\,
            lcout => \current_shift_inst.PI_CTRL.N_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_LC_3_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111011"
        )
    port map (
            in0 => \N__19562\,
            in1 => \N__19556\,
            in2 => \N__19535\,
            in3 => \N__19526\,
            lcout => \pwm_generator_inst.N_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_10_LC_3_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21860\,
            lcout => \N_19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48001\,
            ce => \N__32547\,
            sr => \N__47358\
        );

    \current_shift_inst.PI_CTRL.prop_term_3_LC_3_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27836\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48001\,
            ce => \N__32547\,
            sr => \N__47358\
        );

    \current_shift_inst.PI_CTRL.prop_term_0_LC_3_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27965\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48001\,
            ce => \N__32547\,
            sr => \N__47358\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_3_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19751\,
            in2 => \N__20042\,
            in3 => \N__20041\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_3_8_0_\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_3_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19745\,
            in3 => \N__19733\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_0\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_3_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19967\,
            in2 => \_gnd_net_\,
            in3 => \N__19724\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_1\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_3_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20111\,
            in2 => \_gnd_net_\,
            in3 => \N__19715\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_2\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_3_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19712\,
            in2 => \_gnd_net_\,
            in3 => \N__19706\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_3\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_3_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19703\,
            in2 => \_gnd_net_\,
            in3 => \N__19697\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_4\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_3_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19694\,
            in2 => \_gnd_net_\,
            in3 => \N__19685\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_5\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_3_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19958\,
            in2 => \_gnd_net_\,
            in3 => \N__19952\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_6\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_3_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19949\,
            in3 => \N__19931\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \bfn_3_9_0_\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_3_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011101111000"
        )
    port map (
            in0 => \N__19928\,
            in1 => \N__20040\,
            in2 => \N__19919\,
            in3 => \N__19904\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_10_LC_3_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19775\,
            in1 => \N__20189\,
            in2 => \N__19760\,
            in3 => \N__20333\,
            lcout => \current_shift_inst.PI_CTRL.N_178\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_3_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20651\,
            in1 => \N__20204\,
            in2 => \N__20180\,
            in3 => \N__19766\,
            lcout => \current_shift_inst.PI_CTRL.N_118\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNINKF4_12_LC_3_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21557\,
            in1 => \N__21107\,
            in2 => \N__21932\,
            in3 => \N__21575\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIRO62_11_LC_3_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21556\,
            in2 => \_gnd_net_\,
            in3 => \N__21137\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI4TS8_10_LC_3_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21160\,
            in1 => \N__20198\,
            in2 => \N__19769\,
            in3 => \N__21574\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNID6B4_10_LC_3_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21515\,
            in1 => \N__21473\,
            in2 => \N__21539\,
            in3 => \N__21161\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMK72_20_LC_3_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21664\,
            in2 => \_gnd_net_\,
            in3 => \N__21383\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_9_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIR5H5_12_LC_3_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21625\,
            in1 => \N__21514\,
            in2 => \N__20207\,
            in3 => \N__21106\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIGDF4_19_LC_3_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21701\,
            in1 => \N__21719\,
            in2 => \N__21931\,
            in3 => \N__21406\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI1U52_18_LC_3_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__21407\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21425\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI8JH5_20_LC_3_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21644\,
            in1 => \N__21382\,
            in2 => \N__20192\,
            in3 => \N__21595\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNINID4_13_LC_3_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21469\,
            in1 => \N__21643\,
            in2 => \N__21596\,
            in3 => \N__21538\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_3_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010111001100"
        )
    port map (
            in0 => \N__20168\,
            in1 => \N__20147\,
            in2 => \N__20129\,
            in3 => \N__19996\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_3_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010111001100"
        )
    port map (
            in0 => \N__20099\,
            in1 => \N__20075\,
            in2 => \N__20057\,
            in3 => \N__19995\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_counter_cry_1_c_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20704\,
            in2 => \N__20686\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_5_0_\,
            carryout => un5_counter_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_2_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20269\,
            in2 => \_gnd_net_\,
            in3 => \N__20231\,
            lcout => \counterZ0Z_2\,
            ltout => OPEN,
            carryin => un5_counter_cry_1,
            carryout => un5_counter_cry_2,
            clk => \N__48004\,
            ce => 'H',
            sr => \N__47328\
        );

    \counter_3_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20792\,
            in2 => \_gnd_net_\,
            in3 => \N__20228\,
            lcout => \counterZ0Z_3\,
            ltout => OPEN,
            carryin => un5_counter_cry_2,
            carryout => un5_counter_cry_3,
            clk => \N__48004\,
            ce => 'H',
            sr => \N__47328\
        );

    \counter_4_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20804\,
            in2 => \_gnd_net_\,
            in3 => \N__20225\,
            lcout => \counterZ0Z_4\,
            ltout => OPEN,
            carryin => un5_counter_cry_3,
            carryout => un5_counter_cry_4,
            clk => \N__48004\,
            ce => 'H',
            sr => \N__47328\
        );

    \counter_5_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20780\,
            in2 => \_gnd_net_\,
            in3 => \N__20222\,
            lcout => \counterZ0Z_5\,
            ltout => OPEN,
            carryin => un5_counter_cry_4,
            carryout => un5_counter_cry_5,
            clk => \N__48004\,
            ce => 'H',
            sr => \N__47328\
        );

    \counter_6_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20768\,
            in2 => \_gnd_net_\,
            in3 => \N__20219\,
            lcout => \counterZ0Z_6\,
            ltout => OPEN,
            carryin => un5_counter_cry_5,
            carryout => un5_counter_cry_6,
            clk => \N__48004\,
            ce => 'H',
            sr => \N__47328\
        );

    \counter_RNO_0_7_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20630\,
            in2 => \_gnd_net_\,
            in3 => \N__20216\,
            lcout => \counter_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => un5_counter_cry_6,
            carryout => un5_counter_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_8_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20284\,
            in2 => \_gnd_net_\,
            in3 => \N__20213\,
            lcout => \counterZ0Z_8\,
            ltout => OPEN,
            carryin => un5_counter_cry_7,
            carryout => un5_counter_cry_8,
            clk => \N__48004\,
            ce => 'H',
            sr => \N__47328\
        );

    \counter_9_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20297\,
            in2 => \_gnd_net_\,
            in3 => \N__20210\,
            lcout => \counterZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_4_6_0_\,
            carryout => un5_counter_cry_9,
            clk => \N__48002\,
            ce => 'H',
            sr => \N__47341\
        );

    \counter_RNO_0_10_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20719\,
            in2 => \_gnd_net_\,
            in3 => \N__20321\,
            lcout => \counter_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => un5_counter_cry_9,
            carryout => un5_counter_cry_10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_11_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20311\,
            in2 => \_gnd_net_\,
            in3 => \N__20318\,
            lcout => \counterZ0Z_11\,
            ltout => OPEN,
            carryin => un5_counter_cry_10,
            carryout => un5_counter_cry_11,
            clk => \N__48002\,
            ce => 'H',
            sr => \N__47341\
        );

    \counter_RNO_0_12_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20743\,
            in2 => \_gnd_net_\,
            in3 => \N__20315\,
            lcout => \counter_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIM6001_12_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__20312\,
            in1 => \N__20296\,
            in2 => \N__20744\,
            in3 => \N__20285\,
            lcout => un2_counter_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIRTIM_1_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__20270\,
            in1 => \N__20626\,
            in2 => \N__20720\,
            in3 => \N__20703\,
            lcout => un2_counter_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_4_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__20513\,
            in1 => \N__20447\,
            in2 => \N__20397\,
            in3 => \N__20255\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47997\,
            ce => 'H',
            sr => \N__47359\
        );

    \pwm_generator_inst.threshold_ACC_1_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101010011"
        )
    port map (
            in0 => \N__20446\,
            in1 => \N__20379\,
            in2 => \N__20556\,
            in3 => \N__20249\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47997\,
            ce => 'H',
            sr => \N__47359\
        );

    \pwm_generator_inst.threshold_ACC_5_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__20514\,
            in1 => \N__20448\,
            in2 => \N__20398\,
            in3 => \N__20243\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47997\,
            ce => 'H',
            sr => \N__47359\
        );

    \pwm_generator_inst.threshold_ACC_0_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__20445\,
            in1 => \N__20237\,
            in2 => \N__20555\,
            in3 => \N__20378\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47997\,
            ce => 'H',
            sr => \N__47359\
        );

    \pwm_generator_inst.threshold_ACC_6_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100100111"
        )
    port map (
            in0 => \N__20515\,
            in1 => \N__20449\,
            in2 => \N__20399\,
            in3 => \N__20645\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47997\,
            ce => 'H',
            sr => \N__47359\
        );

    \counter_7_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__21056\,
            in1 => \N__20639\,
            in2 => \N__21092\,
            in3 => \N__21026\,
            lcout => \counterZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47997\,
            ce => 'H',
            sr => \N__47359\
        );

    \pwm_generator_inst.threshold_ACC_7_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100100111"
        )
    port map (
            in0 => \N__20516\,
            in1 => \N__20450\,
            in2 => \N__20400\,
            in3 => \N__20342\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47997\,
            ce => 'H',
            sr => \N__47359\
        );

    \current_shift_inst.PI_CTRL.prop_term_7_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28412\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47994\,
            ce => \N__32485\,
            sr => \N__47369\
        );

    \current_shift_inst.PI_CTRL.prop_term_5_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27656\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47994\,
            ce => \N__32485\,
            sr => \N__47369\
        );

    \current_shift_inst.PI_CTRL.prop_term_10_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28184\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47994\,
            ce => \N__32485\,
            sr => \N__47369\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMIE4_17_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21448\,
            in1 => \N__21700\,
            in2 => \N__21626\,
            in3 => \N__21665\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI2QR8_11_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21494\,
            in1 => \N__20327\,
            in2 => \N__20336\,
            in3 => \N__21136\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMK72_21_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__21682\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21718\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIOIC4_15_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21683\,
            in1 => \N__21493\,
            in2 => \N__21449\,
            in3 => \N__21424\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_8_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28339\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47987\,
            ce => \N__32490\,
            sr => \N__47381\
        );

    \current_shift_inst.PI_CTRL.prop_term_15_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28876\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47987\,
            ce => \N__32490\,
            sr => \N__47381\
        );

    \current_shift_inst.PI_CTRL.prop_term_16_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28792\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47987\,
            ce => \N__32490\,
            sr => \N__47381\
        );

    \current_shift_inst.PI_CTRL.prop_term_11_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28108\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47987\,
            ce => \N__32490\,
            sr => \N__47381\
        );

    \current_shift_inst.PI_CTRL.prop_term_20_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29447\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47987\,
            ce => \N__32490\,
            sr => \N__47381\
        );

    \current_shift_inst.PI_CTRL.prop_term_12_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28030\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47978\,
            ce => \N__32497\,
            sr => \N__47389\
        );

    \current_shift_inst.PI_CTRL.prop_term_21_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29335\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47978\,
            ce => \N__32497\,
            sr => \N__47389\
        );

    \current_shift_inst.PI_CTRL.prop_term_24_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29146\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47978\,
            ce => \N__32497\,
            sr => \N__47389\
        );

    \current_shift_inst.PI_CTRL.prop_term_18_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28633\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47978\,
            ce => \N__32497\,
            sr => \N__47389\
        );

    \GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_4_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20831\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_clk_12mhz_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIN1J6_3_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20803\,
            in2 => \_gnd_net_\,
            in3 => \N__20791\,
            lcout => OPEN,
            ltout => \un2_counter_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIQKFG_5_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__20779\,
            in1 => \N__20767\,
            in2 => \N__20756\,
            in3 => \N__20678\,
            lcout => un2_counter_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_12_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__21091\,
            in1 => \N__21058\,
            in2 => \N__20753\,
            in3 => \N__21023\,
            lcout => \counterZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47999\,
            ce => 'H',
            sr => \N__47329\
        );

    \counter_10_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__21022\,
            in1 => \N__21090\,
            in2 => \N__20729\,
            in3 => \N__21059\,
            lcout => \counterZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47999\,
            ce => 'H',
            sr => \N__47329\
        );

    \counter_1_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__20685\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20705\,
            lcout => \counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47999\,
            ce => 'H',
            sr => \N__47329\
        );

    \counter_0_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__21089\,
            in1 => \N__21057\,
            in2 => \N__20687\,
            in3 => \N__21021\,
            lcout => \counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47999\,
            ce => 'H',
            sr => \N__47329\
        );

    \pwm_generator_inst.threshold_3_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20660\,
            lcout => \pwm_generator_inst.thresholdZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47998\,
            ce => 'H',
            sr => \N__47342\
        );

    \clk_10khz_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__21085\,
            in1 => \N__21055\,
            in2 => \N__22096\,
            in3 => \N__21025\,
            lcout => clk_10khz_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47998\,
            ce => 'H',
            sr => \N__47342\
        );

    \clk_10khz_RNIIENA2_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__21084\,
            in1 => \N__21054\,
            in2 => \N__22092\,
            in3 => \N__21024\,
            lcout => \clk_10khz_RNIIENAZ0Z2\,
            ltout => \clk_10khz_RNIIENAZ0Z2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_cnv_0_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33693\,
            in2 => \N__20993\,
            in3 => \N__22085\,
            lcout => \N_605_g\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__20884\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20845\,
            lcout => \current_shift_inst.PI_CTRL.N_98\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27991\,
            in2 => \N__20978\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_5_9_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\,
            clk => \N__47992\,
            ce => \N__32484\,
            sr => \N__47360\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27929\,
            in2 => \N__21947\,
            in3 => \N__20933\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            clk => \N__47992\,
            ce => \N__32484\,
            sr => \N__47360\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22001\,
            in2 => \N__30040\,
            in3 => \N__20915\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            clk => \N__47992\,
            ce => \N__32484\,
            sr => \N__47360\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27809\,
            in2 => \N__20912\,
            in3 => \N__20873\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            clk => \N__47992\,
            ce => \N__32484\,
            sr => \N__47360\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27754\,
            in2 => \N__21977\,
            in3 => \N__20834\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            clk => \N__47992\,
            ce => \N__32484\,
            sr => \N__47360\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27692\,
            in2 => \N__21359\,
            in3 => \N__21326\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            clk => \N__47992\,
            ce => \N__32484\,
            sr => \N__47360\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28517\,
            in2 => \N__25349\,
            in3 => \N__21296\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            clk => \N__47992\,
            ce => \N__32484\,
            sr => \N__47360\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21293\,
            in2 => \N__28448\,
            in3 => \N__21260\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            clk => \N__47992\,
            ce => \N__32484\,
            sr => \N__47360\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28373\,
            in2 => \N__21257\,
            in3 => \N__21212\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_5_10_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            clk => \N__47988\,
            ce => \N__32432\,
            sr => \N__47370\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28303\,
            in2 => \N__25334\,
            in3 => \N__21173\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            clk => \N__47988\,
            ce => \N__32432\,
            sr => \N__47370\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28220\,
            in2 => \N__21170\,
            in3 => \N__21149\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            clk => \N__47988\,
            ce => \N__32432\,
            sr => \N__47370\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28145\,
            in2 => \N__21146\,
            in3 => \N__21122\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            clk => \N__47988\,
            ce => \N__32432\,
            sr => \N__47370\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28070\,
            in2 => \N__21119\,
            in3 => \N__21095\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            clk => \N__47988\,
            ce => \N__32432\,
            sr => \N__47370\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29056\,
            in2 => \N__21989\,
            in3 => \N__21518\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            clk => \N__47988\,
            ce => \N__32432\,
            sr => \N__47370\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28985\,
            in2 => \N__21959\,
            in3 => \N__21503\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            clk => \N__47988\,
            ce => \N__32432\,
            sr => \N__47370\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21500\,
            in2 => \N__28910\,
            in3 => \N__21482\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            clk => \N__47988\,
            ce => \N__32432\,
            sr => \N__47370\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21479\,
            in2 => \N__28841\,
            in3 => \N__21452\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_5_11_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            clk => \N__47979\,
            ce => \N__32489\,
            sr => \N__47376\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28751\,
            in2 => \N__22166\,
            in3 => \N__21437\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            clk => \N__47979\,
            ce => \N__32489\,
            sr => \N__47376\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28670\,
            in2 => \N__21434\,
            in3 => \N__21410\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            clk => \N__47979\,
            ce => \N__32489\,
            sr => \N__47376\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28592\,
            in2 => \N__21791\,
            in3 => \N__21395\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            clk => \N__47979\,
            ce => \N__32489\,
            sr => \N__47376\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29423\,
            in2 => \N__21392\,
            in3 => \N__21362\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            clk => \N__47979\,
            ce => \N__32489\,
            sr => \N__47376\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21725\,
            in2 => \N__29366\,
            in3 => \N__21704\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            clk => \N__47979\,
            ce => \N__32489\,
            sr => \N__47376\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29296\,
            in2 => \N__22181\,
            in3 => \N__21686\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            clk => \N__47979\,
            ce => \N__32489\,
            sr => \N__47376\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29222\,
            in2 => \N__22115\,
            in3 => \N__21674\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            clk => \N__47979\,
            ce => \N__32489\,
            sr => \N__47376\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21671\,
            in2 => \N__30407\,
            in3 => \N__21647\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_5_12_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            clk => \N__47969\,
            ce => \N__32480\,
            sr => \N__47382\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30356\,
            in2 => \N__22149\,
            in3 => \N__21629\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            clk => \N__47969\,
            ce => \N__32480\,
            sr => \N__47382\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22139\,
            in2 => \N__29114\,
            in3 => \N__21599\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            clk => \N__47969\,
            ce => \N__32480\,
            sr => \N__47382\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32596\,
            in2 => \N__22150\,
            in3 => \N__21578\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            clk => \N__47969\,
            ce => \N__32480\,
            sr => \N__47382\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22143\,
            in2 => \N__29705\,
            in3 => \N__21560\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            clk => \N__47969\,
            ce => \N__32480\,
            sr => \N__47382\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29636\,
            in2 => \N__22151\,
            in3 => \N__21542\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            clk => \N__47969\,
            ce => \N__32480\,
            sr => \N__47382\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22147\,
            in2 => \N__29576\,
            in3 => \N__21902\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\,
            clk => \N__47969\,
            ce => \N__32480\,
            sr => \N__47382\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__22148\,
            in1 => \N__33083\,
            in2 => \_gnd_net_\,
            in3 => \N__21899\,
            lcout => \current_shift_inst.PI_CTRL.un8_enablelto31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47969\,
            ce => \N__32480\,
            sr => \N__47382\
        );

    \current_shift_inst.PI_CTRL.prop_term_19_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28555\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47961\,
            ce => \N__32491\,
            sr => \N__47390\
        );

    \CONSTANT_ONE_LUT4_LC_5_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_6_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21779\,
            lcout => \pwm_generator_inst.thresholdZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47989\,
            ce => 'H',
            sr => \N__47330\
        );

    \pwm_generator_inst.threshold_2_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21770\,
            lcout => \pwm_generator_inst.thresholdZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47989\,
            ce => 'H',
            sr => \N__47330\
        );

    \pwm_generator_inst.threshold_0_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21755\,
            lcout => \pwm_generator_inst.thresholdZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47989\,
            ce => 'H',
            sr => \N__47330\
        );

    \pwm_generator_inst.threshold_5_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21746\,
            lcout => \pwm_generator_inst.thresholdZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47989\,
            ce => 'H',
            sr => \N__47330\
        );

    \pwm_generator_inst.threshold_7_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21737\,
            lcout => \pwm_generator_inst.thresholdZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47989\,
            ce => 'H',
            sr => \N__47330\
        );

    \pwm_generator_inst.threshold_1_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22049\,
            lcout => \pwm_generator_inst.thresholdZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47989\,
            ce => 'H',
            sr => \N__47330\
        );

    \pwm_generator_inst.threshold_4_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22040\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.thresholdZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47989\,
            ce => 'H',
            sr => \N__47330\
        );

    \pwm_generator_inst.threshold_9_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22031\,
            lcout => \pwm_generator_inst.thresholdZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47980\,
            ce => 'H',
            sr => \N__47343\
        );

    \pwm_generator_inst.threshold_8_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22016\,
            lcout => \pwm_generator_inst.thresholdZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47980\,
            ce => 'H',
            sr => \N__47343\
        );

    \current_shift_inst.PI_CTRL.prop_term_2_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27859\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47970\,
            ce => \N__32513\,
            sr => \N__47352\
        );

    \current_shift_inst.PI_CTRL.prop_term_13_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29023\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47970\,
            ce => \N__32513\,
            sr => \N__47352\
        );

    \current_shift_inst.PI_CTRL.prop_term_4_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27721\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47970\,
            ce => \N__32513\,
            sr => \N__47352\
        );

    \current_shift_inst.PI_CTRL.prop_term_14_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28951\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47970\,
            ce => \N__32513\,
            sr => \N__47352\
        );

    \current_shift_inst.PI_CTRL.prop_term_1_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27895\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47970\,
            ce => \N__32513\,
            sr => \N__47352\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__29417\,
            in1 => \N__28591\,
            in2 => \N__29297\,
            in3 => \N__28747\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27690\,
            in2 => \_gnd_net_\,
            in3 => \N__28441\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_22_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29257\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47956\,
            ce => \N__32514\,
            sr => \N__47371\
        );

    \current_shift_inst.PI_CTRL.prop_term_17_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28708\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47956\,
            ce => \N__32514\,
            sr => \N__47371\
        );

    \current_shift_inst.PI_CTRL.prop_term_25_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29510\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47956\,
            ce => \N__32514\,
            sr => \N__47371\
        );

    \current_shift_inst.PI_CTRL.prop_term_23_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29185\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47956\,
            ce => \N__32514\,
            sr => \N__47371\
        );

    \current_shift_inst.phase_valid_RNISLOR2_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__30203\,
            in1 => \N__22100\,
            in2 => \N__33722\,
            in3 => \N__22064\,
            lcout => \current_shift_inst.phase_valid_RNISLORZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_RNO_0_21_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011111100"
        )
    port map (
            in0 => \N__22193\,
            in1 => \N__44200\,
            in2 => \N__39353\,
            in3 => \N__43963\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto31_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_1_c_RNO_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__26489\,
            in1 => \N__27133\,
            in2 => \_gnd_net_\,
            in3 => \N__24913\,
            lcout => \current_shift_inst.un38_control_input_0_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4G5K_25_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31231\,
            in2 => \_gnd_net_\,
            in3 => \N__31140\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI4G5K_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU73K_23_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30596\,
            in2 => \_gnd_net_\,
            in3 => \N__30562\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIU73K_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIB4C81_25_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__31366\,
            in1 => \N__31141\,
            in2 => \N__31235\,
            in3 => \N__31336\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIB4C81_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAO7K_27_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30696\,
            in2 => \_gnd_net_\,
            in3 => \N__30656\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIAO7K_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIKKJ81_29_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__27043\,
            in1 => \N__23122\,
            in2 => \N__27011\,
            in3 => \N__27169\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIKKJ81_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDS8K_28_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27042\,
            in2 => \_gnd_net_\,
            in3 => \N__27007\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIDS8K_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVJ781_23_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__30597\,
            in1 => \N__31271\,
            in2 => \N__30566\,
            in3 => \N__31189\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIVJ781_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7OAK_29_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__27170\,
            in1 => \_gnd_net_\,
            in2 => \N__23126\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI7OAK_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJTQ51_12_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001111000011"
        )
    port map (
            in0 => \N__30845\,
            in1 => \N__25681\,
            in2 => \N__26648\,
            in3 => \N__30762\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJTQ51_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR0UI_13_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__25680\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26643\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIR0UI_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_2_c_RNO_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001100110"
        )
    port map (
            in0 => \N__22639\,
            in1 => \N__27119\,
            in2 => \N__26456\,
            in3 => \N__24909\,
            lcout => \current_shift_inst.un38_control_input_0_cry_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_2_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23339\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47919\,
            ce => \N__22388\,
            sr => \N__47398\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8SSQ5_15_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010001"
        )
    port map (
            in0 => \N__42026\,
            in1 => \N__44156\,
            in2 => \N__42380\,
            in3 => \N__36845\,
            lcout => \delay_measurement_inst.delay_hc_reg3lt19_0\,
            ltout => \delay_measurement_inst.delay_hc_reg3lt19_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_31_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011101110"
        )
    port map (
            in0 => \N__39352\,
            in1 => \N__44204\,
            in2 => \N__22184\,
            in3 => \N__43967\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto31_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_1_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23366\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47919\,
            ce => \N__22388\,
            sr => \N__47398\
        );

    \current_shift_inst.control_input_RNO_0_25_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110010110"
        )
    port map (
            in0 => \N__27065\,
            in1 => \N__25297\,
            in2 => \N__27132\,
            in3 => \N__22741\,
            lcout => \current_shift_inst.un38_control_input_0_axb_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQF91_30_LC_7_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__25027\,
            in1 => \N__22740\,
            in2 => \_gnd_net_\,
            in3 => \N__27064\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIVQF91_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31931\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47913\,
            ce => \N__31953\,
            sr => \N__47402\
        );

    \current_shift_inst.un38_control_input_0_cry_3_c_inv_RNO_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101100101"
        )
    port map (
            in0 => \N__22611\,
            in1 => \N__22635\,
            in2 => \N__27131\,
            in3 => \N__24907\,
            lcout => \current_shift_inst.N_1620_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5LGN1_3_LC_7_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__24908\,
            in1 => \N__22612\,
            in2 => \N__22640\,
            in3 => \N__27112\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_3_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23362\,
            in2 => \N__23312\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_3\,
            ltout => OPEN,
            carryin => \bfn_7_19_0_\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_2\,
            clk => \N__47907\,
            ce => \N__22387\,
            sr => \N__47405\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_4_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23335\,
            in2 => \N__23281\,
            in3 => \N__22217\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_2\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_3\,
            clk => \N__47907\,
            ce => \N__22387\,
            sr => \N__47405\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_5_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23311\,
            in2 => \N__23254\,
            in3 => \N__22214\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_3\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_4\,
            clk => \N__47907\,
            ce => \N__22387\,
            sr => \N__47405\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_6_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23224\,
            in2 => \N__23282\,
            in3 => \N__22211\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_4\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_5\,
            clk => \N__47907\,
            ce => \N__22387\,
            sr => \N__47405\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_7_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23200\,
            in2 => \N__23255\,
            in3 => \N__22208\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_5\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_6\,
            clk => \N__47907\,
            ce => \N__22387\,
            sr => \N__47405\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_8_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23225\,
            in2 => \N__23177\,
            in3 => \N__22205\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_6\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_7\,
            clk => \N__47907\,
            ce => \N__22387\,
            sr => \N__47405\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_9_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23201\,
            in2 => \N__23612\,
            in3 => \N__22202\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_7\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_8\,
            clk => \N__47907\,
            ce => \N__22387\,
            sr => \N__47405\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_10_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23176\,
            in2 => \N__23576\,
            in3 => \N__22199\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_8\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_9\,
            clk => \N__47907\,
            ce => \N__22387\,
            sr => \N__47405\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_11_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23548\,
            in2 => \N__23611\,
            in3 => \N__22196\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_11\,
            ltout => OPEN,
            carryin => \bfn_7_20_0_\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_10\,
            clk => \N__47902\,
            ce => \N__22386\,
            sr => \N__47408\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_12_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23575\,
            in2 => \N__23527\,
            in3 => \N__22244\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_10\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_11\,
            clk => \N__47902\,
            ce => \N__22386\,
            sr => \N__47408\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_13_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23549\,
            in2 => \N__23500\,
            in3 => \N__22241\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_11\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_12\,
            clk => \N__47902\,
            ce => \N__22386\,
            sr => \N__47408\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_14_LC_7_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23467\,
            in2 => \N__23528\,
            in3 => \N__22238\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_12\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_13\,
            clk => \N__47902\,
            ce => \N__22386\,
            sr => \N__47408\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_15_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23440\,
            in2 => \N__23501\,
            in3 => \N__22235\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_13\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_14\,
            clk => \N__47902\,
            ce => \N__22386\,
            sr => \N__47408\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_16_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23416\,
            in2 => \N__23471\,
            in3 => \N__22232\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_14\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_15\,
            clk => \N__47902\,
            ce => \N__22386\,
            sr => \N__47408\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_17_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23441\,
            in2 => \N__23396\,
            in3 => \N__22229\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_15\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_16\,
            clk => \N__47902\,
            ce => \N__22386\,
            sr => \N__47408\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_18_LC_7_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23417\,
            in2 => \N__23837\,
            in3 => \N__22226\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_16\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_17\,
            clk => \N__47902\,
            ce => \N__22386\,
            sr => \N__47408\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_19_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23392\,
            in2 => \N__23804\,
            in3 => \N__22223\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_19\,
            ltout => OPEN,
            carryin => \bfn_7_21_0_\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_18\,
            clk => \N__47895\,
            ce => \N__22385\,
            sr => \N__47412\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_20_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23770\,
            in2 => \N__23836\,
            in3 => \N__22220\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_18\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_19\,
            clk => \N__47895\,
            ce => \N__22385\,
            sr => \N__47412\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_21_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23800\,
            in2 => \N__23746\,
            in3 => \N__22271\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_19\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_20\,
            clk => \N__47895\,
            ce => \N__22385\,
            sr => \N__47412\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_22_LC_7_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23771\,
            in2 => \N__23716\,
            in3 => \N__22268\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_20\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_21\,
            clk => \N__47895\,
            ce => \N__22385\,
            sr => \N__47412\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_23_LC_7_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23686\,
            in2 => \N__23747\,
            in3 => \N__22265\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_21\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_22\,
            clk => \N__47895\,
            ce => \N__22385\,
            sr => \N__47412\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_24_LC_7_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23662\,
            in2 => \N__23717\,
            in3 => \N__22262\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_22\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_23\,
            clk => \N__47895\,
            ce => \N__22385\,
            sr => \N__47412\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_25_LC_7_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23687\,
            in2 => \N__23642\,
            in3 => \N__22259\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_23\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_24\,
            clk => \N__47895\,
            ce => \N__22385\,
            sr => \N__47412\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_26_LC_7_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23663\,
            in2 => \N__24149\,
            in3 => \N__22256\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_24\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_25\,
            clk => \N__47895\,
            ce => \N__22385\,
            sr => \N__47412\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_27_LC_7_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23638\,
            in2 => \N__24113\,
            in3 => \N__22253\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_27\,
            ltout => OPEN,
            carryin => \bfn_7_22_0_\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_26\,
            clk => \N__47889\,
            ce => \N__22384\,
            sr => \N__47414\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_28_LC_7_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24082\,
            in2 => \N__24148\,
            in3 => \N__22250\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_26\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_27\,
            clk => \N__47889\,
            ce => \N__22384\,
            sr => \N__47414\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_29_LC_7_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24112\,
            in2 => \N__24062\,
            in3 => \N__22247\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_27\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_28\,
            clk => \N__47889\,
            ce => \N__22384\,
            sr => \N__47414\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_30_LC_7_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24083\,
            in2 => \N__24038\,
            in3 => \N__22394\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_28\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_29\,
            clk => \N__47889\,
            ce => \N__22384\,
            sr => \N__47414\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_31_LC_7_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22391\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47889\,
            ce => \N__22384\,
            sr => \N__47414\
        );

    \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22367\,
            in2 => \N__22361\,
            in3 => \N__24468\,
            lcout => \pwm_generator_inst.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_8_8_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22352\,
            in2 => \N__22346\,
            in3 => \N__24384\,
            lcout => \pwm_generator_inst.counter_i_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_0\,
            carryout => \pwm_generator_inst.un14_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22328\,
            in2 => \N__22337\,
            in3 => \N__24489\,
            lcout => \pwm_generator_inst.counter_i_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_1\,
            carryout => \pwm_generator_inst.un14_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22307\,
            in2 => \N__22322\,
            in3 => \N__24405\,
            lcout => \pwm_generator_inst.counter_i_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_2\,
            carryout => \pwm_generator_inst.un14_counter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22301\,
            in2 => \N__22295\,
            in3 => \N__24360\,
            lcout => \pwm_generator_inst.counter_i_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_3\,
            carryout => \pwm_generator_inst.un14_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22286\,
            in2 => \N__22280\,
            in3 => \N__24315\,
            lcout => \pwm_generator_inst.counter_i_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_4\,
            carryout => \pwm_generator_inst.un14_counter_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22481\,
            in2 => \N__22475\,
            in3 => \N__24339\,
            lcout => \pwm_generator_inst.counter_i_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_5\,
            carryout => \pwm_generator_inst.un14_counter_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22457\,
            in2 => \N__22466\,
            in3 => \N__24213\,
            lcout => \pwm_generator_inst.counter_i_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_6\,
            carryout => \pwm_generator_inst.un14_counter_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22442\,
            in2 => \N__22451\,
            in3 => \N__24235\,
            lcout => \pwm_generator_inst.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_8_9_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22427\,
            in2 => \N__22436\,
            in3 => \N__24255\,
            lcout => \pwm_generator_inst.counter_i_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_8\,
            carryout => \pwm_generator_inst.un14_counter_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.pwm_out_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22421\,
            lcout => pwm_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47971\,
            ce => 'H',
            sr => \N__47331\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__30041\,
            in1 => \N__27922\,
            in2 => \_gnd_net_\,
            in3 => \N__27992\,
            lcout => \current_shift_inst.PI_CTRL.un1_enablelt3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__28984\,
            in1 => \N__28833\,
            in2 => \N__29057\,
            in3 => \N__28144\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__29216\,
            in1 => \N__28906\,
            in2 => \N__29631\,
            in3 => \N__28212\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__29694\,
            in1 => \N__32588\,
            in2 => \N__28069\,
            in3 => \N__29561\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIA31P2_10_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22535\,
            in1 => \N__22529\,
            in2 => \N__22523\,
            in3 => \N__22520\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28365\,
            in1 => \N__28509\,
            in2 => \N__28296\,
            in3 => \N__28440\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__27760\,
            in1 => \N__27804\,
            in2 => \N__22514\,
            in3 => \N__27691\,
            lcout => \current_shift_inst.PI_CTRL.N_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__28510\,
            in1 => \N__28366\,
            in2 => \N__28304\,
            in3 => \N__22511\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110011"
        )
    port map (
            in0 => \N__22505\,
            in1 => \N__27761\,
            in2 => \N__22499\,
            in3 => \N__27805\,
            lcout => \current_shift_inst.PI_CTRL.N_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_21_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__36819\,
            in1 => \N__40724\,
            in2 => \_gnd_net_\,
            in3 => \N__22496\,
            lcout => measured_delay_hc_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47953\,
            ce => 'H',
            sr => \N__47361\
        );

    \current_shift_inst.control_input_0_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24608\,
            in2 => \N__29948\,
            in3 => \N__29947\,
            lcout => \current_shift_inst.control_inputZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_13_0_\,
            carryout => \current_shift_inst.control_input_1_cry_0\,
            clk => \N__47944\,
            ce => \N__24952\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_1_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24599\,
            in2 => \_gnd_net_\,
            in3 => \N__22487\,
            lcout => \current_shift_inst.control_inputZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_0\,
            carryout => \current_shift_inst.control_input_1_cry_1\,
            clk => \N__47944\,
            ce => \N__24952\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_2_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24590\,
            in2 => \_gnd_net_\,
            in3 => \N__22484\,
            lcout => \current_shift_inst.control_inputZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_1\,
            carryout => \current_shift_inst.control_input_1_cry_2\,
            clk => \N__47944\,
            ce => \N__24952\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_3_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24581\,
            in2 => \_gnd_net_\,
            in3 => \N__22562\,
            lcout => \current_shift_inst.control_inputZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_2\,
            carryout => \current_shift_inst.control_input_1_cry_3\,
            clk => \N__47944\,
            ce => \N__24952\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_4_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24572\,
            in2 => \_gnd_net_\,
            in3 => \N__22559\,
            lcout => \current_shift_inst.control_inputZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_3\,
            carryout => \current_shift_inst.control_input_1_cry_4\,
            clk => \N__47944\,
            ce => \N__24952\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_5_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24563\,
            in2 => \_gnd_net_\,
            in3 => \N__22556\,
            lcout => \current_shift_inst.control_inputZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_4\,
            carryout => \current_shift_inst.control_input_1_cry_5\,
            clk => \N__47944\,
            ce => \N__24952\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_6_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24713\,
            in2 => \_gnd_net_\,
            in3 => \N__22553\,
            lcout => \current_shift_inst.control_inputZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_5\,
            carryout => \current_shift_inst.control_input_1_cry_6\,
            clk => \N__47944\,
            ce => \N__24952\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_7_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24692\,
            in2 => \_gnd_net_\,
            in3 => \N__22550\,
            lcout => \current_shift_inst.control_inputZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_6\,
            carryout => \current_shift_inst.control_input_1_cry_7\,
            clk => \N__47944\,
            ce => \N__24952\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_8_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24671\,
            in2 => \_gnd_net_\,
            in3 => \N__22547\,
            lcout => \current_shift_inst.control_inputZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_14_0_\,
            carryout => \current_shift_inst.control_input_1_cry_8\,
            clk => \N__47935\,
            ce => \N__24968\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_9_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24662\,
            in2 => \_gnd_net_\,
            in3 => \N__22544\,
            lcout => \current_shift_inst.control_inputZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_8\,
            carryout => \current_shift_inst.control_input_1_cry_9\,
            clk => \N__47935\,
            ce => \N__24968\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_10_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24653\,
            in2 => \_gnd_net_\,
            in3 => \N__22541\,
            lcout => \current_shift_inst.control_inputZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_9\,
            carryout => \current_shift_inst.control_input_1_cry_10\,
            clk => \N__47935\,
            ce => \N__24968\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_11_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24644\,
            in2 => \_gnd_net_\,
            in3 => \N__22538\,
            lcout => \current_shift_inst.control_inputZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_10\,
            carryout => \current_shift_inst.control_input_1_cry_11\,
            clk => \N__47935\,
            ce => \N__24968\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_12_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24635\,
            in2 => \_gnd_net_\,
            in3 => \N__22589\,
            lcout => \current_shift_inst.control_inputZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_11\,
            carryout => \current_shift_inst.control_input_1_cry_12\,
            clk => \N__47935\,
            ce => \N__24968\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_13_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24626\,
            in2 => \_gnd_net_\,
            in3 => \N__22586\,
            lcout => \current_shift_inst.control_inputZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_12\,
            carryout => \current_shift_inst.control_input_1_cry_13\,
            clk => \N__47935\,
            ce => \N__24968\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_14_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24617\,
            in2 => \_gnd_net_\,
            in3 => \N__22583\,
            lcout => \current_shift_inst.control_inputZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_13\,
            carryout => \current_shift_inst.control_input_1_cry_14\,
            clk => \N__47935\,
            ce => \N__24968\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_15_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24839\,
            in2 => \_gnd_net_\,
            in3 => \N__22580\,
            lcout => \current_shift_inst.control_inputZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_14\,
            carryout => \current_shift_inst.control_input_1_cry_15\,
            clk => \N__47935\,
            ce => \N__24968\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_16_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24830\,
            in2 => \_gnd_net_\,
            in3 => \N__22577\,
            lcout => \current_shift_inst.control_inputZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_8_15_0_\,
            carryout => \current_shift_inst.control_input_1_cry_16\,
            clk => \N__47926\,
            ce => \N__24959\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_17_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24821\,
            in2 => \_gnd_net_\,
            in3 => \N__22574\,
            lcout => \current_shift_inst.control_inputZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_16\,
            carryout => \current_shift_inst.control_input_1_cry_17\,
            clk => \N__47926\,
            ce => \N__24959\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_18_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24791\,
            in2 => \_gnd_net_\,
            in3 => \N__22571\,
            lcout => \current_shift_inst.control_inputZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_17\,
            carryout => \current_shift_inst.control_input_1_cry_18\,
            clk => \N__47926\,
            ce => \N__24959\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_19_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24782\,
            in2 => \_gnd_net_\,
            in3 => \N__22568\,
            lcout => \current_shift_inst.control_inputZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_18\,
            carryout => \current_shift_inst.control_input_1_cry_19\,
            clk => \N__47926\,
            ce => \N__24959\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_20_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24752\,
            in2 => \_gnd_net_\,
            in3 => \N__22565\,
            lcout => \current_shift_inst.control_inputZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_19\,
            carryout => \current_shift_inst.control_input_1_cry_20\,
            clk => \N__47926\,
            ce => \N__24959\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_21_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24743\,
            in2 => \_gnd_net_\,
            in3 => \N__22655\,
            lcout => \current_shift_inst.control_inputZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_20\,
            carryout => \current_shift_inst.control_input_1_cry_21\,
            clk => \N__47926\,
            ce => \N__24959\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_22_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24722\,
            in2 => \_gnd_net_\,
            in3 => \N__22652\,
            lcout => \current_shift_inst.control_inputZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_21\,
            carryout => \current_shift_inst.control_input_1_cry_22\,
            clk => \N__47926\,
            ce => \N__24959\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_23_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25049\,
            in2 => \_gnd_net_\,
            in3 => \N__22649\,
            lcout => \current_shift_inst.control_inputZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_22\,
            carryout => \current_shift_inst.control_input_1_cry_23\,
            clk => \N__47926\,
            ce => \N__24959\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_24_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25001\,
            in2 => \_gnd_net_\,
            in3 => \N__22646\,
            lcout => \current_shift_inst.control_inputZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_8_16_0_\,
            carryout => \current_shift_inst.control_input_1_cry_24\,
            clk => \N__47920\,
            ce => \N__24966\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_1_cry_24_THRU_LUT4_0_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22643\,
            lcout => \current_shift_inst.control_input_1_cry_24_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_1_c_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24900\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_17_0_\,
            carryout => \current_shift_inst.z_5_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_2_s_LC_8_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22634\,
            in2 => \N__23032\,
            in3 => \N__22616\,
            lcout => \current_shift_inst.z_5_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_1\,
            carryout => \current_shift_inst.z_5_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_3_s_LC_8_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22613\,
            in2 => \N__23035\,
            in3 => \N__22595\,
            lcout => \current_shift_inst.z_5_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_2\,
            carryout => \current_shift_inst.z_5_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_4_s_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25590\,
            in2 => \N__23033\,
            in3 => \N__22592\,
            lcout => \current_shift_inst.z_5_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_3\,
            carryout => \current_shift_inst.z_5_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_5_s_LC_8_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25630\,
            in2 => \N__23036\,
            in3 => \N__22682\,
            lcout => \current_shift_inst.z_5_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_4\,
            carryout => \current_shift_inst.z_5_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_6_s_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25488\,
            in2 => \N__23034\,
            in3 => \N__22679\,
            lcout => \current_shift_inst.z_5_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_5\,
            carryout => \current_shift_inst.z_5_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_7_s_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22967\,
            in2 => \N__25880\,
            in3 => \N__22676\,
            lcout => \current_shift_inst.z_5_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_6\,
            carryout => \current_shift_inst.z_5_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_8_s_LC_8_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22974\,
            in2 => \N__25739\,
            in3 => \N__22673\,
            lcout => \current_shift_inst.z_5_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_7\,
            carryout => \current_shift_inst.z_5_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_9_s_LC_8_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25753\,
            in2 => \N__23088\,
            in3 => \N__22670\,
            lcout => \current_shift_inst.z_5_9\,
            ltout => OPEN,
            carryin => \bfn_8_18_0_\,
            carryout => \current_shift_inst.z_5_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_10_s_LC_8_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25909\,
            in2 => \N__23084\,
            in3 => \N__22667\,
            lcout => \current_shift_inst.z_5_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_9\,
            carryout => \current_shift_inst.z_5_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_11_s_LC_8_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30867\,
            in2 => \N__23086\,
            in3 => \N__22664\,
            lcout => \current_shift_inst.z_5_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_10\,
            carryout => \current_shift_inst.z_5_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_12_s_LC_8_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30746\,
            in2 => \N__23085\,
            in3 => \N__22661\,
            lcout => \current_shift_inst.z_5_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_11\,
            carryout => \current_shift_inst.z_5_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_13_s_LC_8_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25676\,
            in2 => \N__23087\,
            in3 => \N__22658\,
            lcout => \current_shift_inst.z_5_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_12\,
            carryout => \current_shift_inst.z_5_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_14_s_LC_8_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23050\,
            in2 => \N__25826\,
            in3 => \N__22709\,
            lcout => \current_shift_inst.z_5_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_13\,
            carryout => \current_shift_inst.z_5_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_15_s_LC_8_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23043\,
            in2 => \N__26139\,
            in3 => \N__22706\,
            lcout => \current_shift_inst.z_5_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_14\,
            carryout => \current_shift_inst.z_5_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_16_s_LC_8_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23051\,
            in2 => \N__26187\,
            in3 => \N__22703\,
            lcout => \current_shift_inst.z_5_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_15\,
            carryout => \current_shift_inst.z_5_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_17_s_LC_8_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26005\,
            in2 => \N__23027\,
            in3 => \N__22700\,
            lcout => \current_shift_inst.z_5_17\,
            ltout => OPEN,
            carryin => \bfn_8_19_0_\,
            carryout => \current_shift_inst.z_5_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_18_s_LC_8_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25971\,
            in2 => \N__23030\,
            in3 => \N__22697\,
            lcout => \current_shift_inst.z_5_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_17\,
            carryout => \current_shift_inst.z_5_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_19_s_LC_8_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26218\,
            in2 => \N__23028\,
            in3 => \N__22694\,
            lcout => \current_shift_inst.z_5_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_18\,
            carryout => \current_shift_inst.z_5_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_20_s_LC_8_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26086\,
            in2 => \N__23031\,
            in3 => \N__22691\,
            lcout => \current_shift_inst.z_5_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_19\,
            carryout => \current_shift_inst.z_5_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_21_s_LC_8_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26049\,
            in2 => \N__23029\,
            in3 => \N__22688\,
            lcout => \current_shift_inst.z_5_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_20\,
            carryout => \current_shift_inst.z_5_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_22_s_LC_8_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22949\,
            in2 => \N__30506\,
            in3 => \N__22685\,
            lcout => \current_shift_inst.z_5_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_21\,
            carryout => \current_shift_inst.z_5_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_23_s_LC_8_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22957\,
            in2 => \N__30598\,
            in3 => \N__23144\,
            lcout => \current_shift_inst.z_5_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_22\,
            carryout => \current_shift_inst.z_5_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_24_s_LC_8_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22950\,
            in2 => \N__31275\,
            in3 => \N__23141\,
            lcout => \current_shift_inst.z_5_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_23\,
            carryout => \current_shift_inst.z_5_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_25_s_LC_8_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31128\,
            in2 => \N__22874\,
            in3 => \N__23138\,
            lcout => \current_shift_inst.z_5_25\,
            ltout => OPEN,
            carryin => \bfn_8_20_0_\,
            carryout => \current_shift_inst.z_5_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_26_s_LC_8_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31353\,
            in2 => \N__22877\,
            in3 => \N__23135\,
            lcout => \current_shift_inst.z_5_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_25\,
            carryout => \current_shift_inst.z_5_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_27_s_LC_8_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30683\,
            in2 => \N__22875\,
            in3 => \N__23132\,
            lcout => \current_shift_inst.z_5_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_26\,
            carryout => \current_shift_inst.z_5_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_28_s_LC_8_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27038\,
            in2 => \N__22878\,
            in3 => \N__23129\,
            lcout => \current_shift_inst.z_5_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_27\,
            carryout => \current_shift_inst.z_5_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_29_s_LC_8_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23121\,
            in2 => \N__22876\,
            in3 => \N__23102\,
            lcout => \current_shift_inst.z_5_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_28\,
            carryout => \current_shift_inst.z_5_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_30_s_LC_8_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22838\,
            in2 => \N__22742\,
            in3 => \N__22715\,
            lcout => \current_shift_inst.z_5_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_29\,
            carryout => \current_shift_inst.z_5_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.z_5_cry_30_THRU_LUT4_0_LC_8_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22712\,
            lcout => \current_shift_inst.z_5_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.counter_0_LC_8_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23955\,
            in1 => \N__23355\,
            in2 => \_gnd_net_\,
            in3 => \N__23342\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_21_0_\,
            carryout => \current_shift_inst.timer_phase.counter_cry_0\,
            clk => \N__47890\,
            ce => \N__24005\,
            sr => \N__47409\
        );

    \current_shift_inst.timer_phase.counter_1_LC_8_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23950\,
            in1 => \N__23328\,
            in2 => \_gnd_net_\,
            in3 => \N__23315\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_0\,
            carryout => \current_shift_inst.timer_phase.counter_cry_1\,
            clk => \N__47890\,
            ce => \N__24005\,
            sr => \N__47409\
        );

    \current_shift_inst.timer_phase.counter_2_LC_8_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23956\,
            in1 => \N__23307\,
            in2 => \_gnd_net_\,
            in3 => \N__23285\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_1\,
            carryout => \current_shift_inst.timer_phase.counter_cry_2\,
            clk => \N__47890\,
            ce => \N__24005\,
            sr => \N__47409\
        );

    \current_shift_inst.timer_phase.counter_3_LC_8_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23951\,
            in1 => \N__23274\,
            in2 => \_gnd_net_\,
            in3 => \N__23258\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_2\,
            carryout => \current_shift_inst.timer_phase.counter_cry_3\,
            clk => \N__47890\,
            ce => \N__24005\,
            sr => \N__47409\
        );

    \current_shift_inst.timer_phase.counter_4_LC_8_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23957\,
            in1 => \N__23242\,
            in2 => \_gnd_net_\,
            in3 => \N__23228\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_3\,
            carryout => \current_shift_inst.timer_phase.counter_cry_4\,
            clk => \N__47890\,
            ce => \N__24005\,
            sr => \N__47409\
        );

    \current_shift_inst.timer_phase.counter_5_LC_8_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23952\,
            in1 => \N__23218\,
            in2 => \_gnd_net_\,
            in3 => \N__23204\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_4\,
            carryout => \current_shift_inst.timer_phase.counter_cry_5\,
            clk => \N__47890\,
            ce => \N__24005\,
            sr => \N__47409\
        );

    \current_shift_inst.timer_phase.counter_6_LC_8_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23954\,
            in1 => \N__23194\,
            in2 => \_gnd_net_\,
            in3 => \N__23180\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_5\,
            carryout => \current_shift_inst.timer_phase.counter_cry_6\,
            clk => \N__47890\,
            ce => \N__24005\,
            sr => \N__47409\
        );

    \current_shift_inst.timer_phase.counter_7_LC_8_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23953\,
            in1 => \N__23161\,
            in2 => \_gnd_net_\,
            in3 => \N__23147\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_6\,
            carryout => \current_shift_inst.timer_phase.counter_cry_7\,
            clk => \N__47890\,
            ce => \N__24005\,
            sr => \N__47409\
        );

    \current_shift_inst.timer_phase.counter_8_LC_8_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23949\,
            in1 => \N__23601\,
            in2 => \_gnd_net_\,
            in3 => \N__23579\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_22_0_\,
            carryout => \current_shift_inst.timer_phase.counter_cry_8\,
            clk => \N__47884\,
            ce => \N__24000\,
            sr => \N__47413\
        );

    \current_shift_inst.timer_phase.counter_9_LC_8_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23961\,
            in1 => \N__23571\,
            in2 => \_gnd_net_\,
            in3 => \N__23552\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_8\,
            carryout => \current_shift_inst.timer_phase.counter_cry_9\,
            clk => \N__47884\,
            ce => \N__24000\,
            sr => \N__47413\
        );

    \current_shift_inst.timer_phase.counter_10_LC_8_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23946\,
            in1 => \N__23547\,
            in2 => \_gnd_net_\,
            in3 => \N__23531\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_9\,
            carryout => \current_shift_inst.timer_phase.counter_cry_10\,
            clk => \N__47884\,
            ce => \N__24000\,
            sr => \N__47413\
        );

    \current_shift_inst.timer_phase.counter_11_LC_8_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23958\,
            in1 => \N__23520\,
            in2 => \_gnd_net_\,
            in3 => \N__23504\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_10\,
            carryout => \current_shift_inst.timer_phase.counter_cry_11\,
            clk => \N__47884\,
            ce => \N__24000\,
            sr => \N__47413\
        );

    \current_shift_inst.timer_phase.counter_12_LC_8_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23947\,
            in1 => \N__23488\,
            in2 => \_gnd_net_\,
            in3 => \N__23474\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_11\,
            carryout => \current_shift_inst.timer_phase.counter_cry_12\,
            clk => \N__47884\,
            ce => \N__24000\,
            sr => \N__47413\
        );

    \current_shift_inst.timer_phase.counter_13_LC_8_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23959\,
            in1 => \N__23460\,
            in2 => \_gnd_net_\,
            in3 => \N__23444\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_12\,
            carryout => \current_shift_inst.timer_phase.counter_cry_13\,
            clk => \N__47884\,
            ce => \N__24000\,
            sr => \N__47413\
        );

    \current_shift_inst.timer_phase.counter_14_LC_8_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23948\,
            in1 => \N__23434\,
            in2 => \_gnd_net_\,
            in3 => \N__23420\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_13\,
            carryout => \current_shift_inst.timer_phase.counter_cry_14\,
            clk => \N__47884\,
            ce => \N__24000\,
            sr => \N__47413\
        );

    \current_shift_inst.timer_phase.counter_15_LC_8_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23960\,
            in1 => \N__23415\,
            in2 => \_gnd_net_\,
            in3 => \N__23399\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_14\,
            carryout => \current_shift_inst.timer_phase.counter_cry_15\,
            clk => \N__47884\,
            ce => \N__24000\,
            sr => \N__47413\
        );

    \current_shift_inst.timer_phase.counter_16_LC_8_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23962\,
            in1 => \N__23388\,
            in2 => \_gnd_net_\,
            in3 => \N__23369\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_8_23_0_\,
            carryout => \current_shift_inst.timer_phase.counter_cry_16\,
            clk => \N__47881\,
            ce => \N__24001\,
            sr => \N__47415\
        );

    \current_shift_inst.timer_phase.counter_17_LC_8_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23966\,
            in1 => \N__23826\,
            in2 => \_gnd_net_\,
            in3 => \N__23807\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_16\,
            carryout => \current_shift_inst.timer_phase.counter_cry_17\,
            clk => \N__47881\,
            ce => \N__24001\,
            sr => \N__47415\
        );

    \current_shift_inst.timer_phase.counter_18_LC_8_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23963\,
            in1 => \N__23799\,
            in2 => \_gnd_net_\,
            in3 => \N__23774\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_17\,
            carryout => \current_shift_inst.timer_phase.counter_cry_18\,
            clk => \N__47881\,
            ce => \N__24001\,
            sr => \N__47415\
        );

    \current_shift_inst.timer_phase.counter_19_LC_8_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23967\,
            in1 => \N__23769\,
            in2 => \_gnd_net_\,
            in3 => \N__23750\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_18\,
            carryout => \current_shift_inst.timer_phase.counter_cry_19\,
            clk => \N__47881\,
            ce => \N__24001\,
            sr => \N__47415\
        );

    \current_shift_inst.timer_phase.counter_20_LC_8_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23964\,
            in1 => \N__23734\,
            in2 => \_gnd_net_\,
            in3 => \N__23720\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_19\,
            carryout => \current_shift_inst.timer_phase.counter_cry_20\,
            clk => \N__47881\,
            ce => \N__24001\,
            sr => \N__47415\
        );

    \current_shift_inst.timer_phase.counter_21_LC_8_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23968\,
            in1 => \N__23704\,
            in2 => \_gnd_net_\,
            in3 => \N__23690\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_20\,
            carryout => \current_shift_inst.timer_phase.counter_cry_21\,
            clk => \N__47881\,
            ce => \N__24001\,
            sr => \N__47415\
        );

    \current_shift_inst.timer_phase.counter_22_LC_8_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23965\,
            in1 => \N__23680\,
            in2 => \_gnd_net_\,
            in3 => \N__23666\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_21\,
            carryout => \current_shift_inst.timer_phase.counter_cry_22\,
            clk => \N__47881\,
            ce => \N__24001\,
            sr => \N__47415\
        );

    \current_shift_inst.timer_phase.counter_23_LC_8_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23969\,
            in1 => \N__23661\,
            in2 => \_gnd_net_\,
            in3 => \N__23645\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_22\,
            carryout => \current_shift_inst.timer_phase.counter_cry_23\,
            clk => \N__47881\,
            ce => \N__24001\,
            sr => \N__47415\
        );

    \current_shift_inst.timer_phase.counter_24_LC_8_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23940\,
            in1 => \N__23634\,
            in2 => \_gnd_net_\,
            in3 => \N__23615\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_8_24_0_\,
            carryout => \current_shift_inst.timer_phase.counter_cry_24\,
            clk => \N__47875\,
            ce => \N__23985\,
            sr => \N__47417\
        );

    \current_shift_inst.timer_phase.counter_25_LC_8_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23944\,
            in1 => \N__24135\,
            in2 => \_gnd_net_\,
            in3 => \N__24116\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_24\,
            carryout => \current_shift_inst.timer_phase.counter_cry_25\,
            clk => \N__47875\,
            ce => \N__23985\,
            sr => \N__47417\
        );

    \current_shift_inst.timer_phase.counter_26_LC_8_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23941\,
            in1 => \N__24108\,
            in2 => \_gnd_net_\,
            in3 => \N__24086\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_25\,
            carryout => \current_shift_inst.timer_phase.counter_cry_26\,
            clk => \N__47875\,
            ce => \N__23985\,
            sr => \N__47417\
        );

    \current_shift_inst.timer_phase.counter_27_LC_8_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23945\,
            in1 => \N__24081\,
            in2 => \_gnd_net_\,
            in3 => \N__24065\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_26\,
            carryout => \current_shift_inst.timer_phase.counter_cry_27\,
            clk => \N__47875\,
            ce => \N__23985\,
            sr => \N__47417\
        );

    \current_shift_inst.timer_phase.counter_28_LC_8_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23942\,
            in1 => \N__24058\,
            in2 => \_gnd_net_\,
            in3 => \N__24044\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_27\,
            carryout => \current_shift_inst.timer_phase.counter_cry_28\,
            clk => \N__47875\,
            ce => \N__23985\,
            sr => \N__47417\
        );

    \current_shift_inst.timer_phase.counter_29_LC_8_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__24034\,
            in1 => \N__23943\,
            in2 => \_gnd_net_\,
            in3 => \N__24041\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47875\,
            ce => \N__23985\,
            sr => \N__47417\
        );

    \current_shift_inst.timer_s1.running_RNII51H_LC_8_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27563\,
            in2 => \_gnd_net_\,
            in3 => \N__27539\,
            lcout => \current_shift_inst.timer_s1.N_187_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.running_RNIL91O_LC_8_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__27472\,
            in1 => \N__25263\,
            in2 => \_gnd_net_\,
            in3 => \N__27452\,
            lcout => \current_shift_inst.timer_phase.N_193_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.running_RNIB31B_LC_8_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27471\,
            lcout => \current_shift_inst.timer_phase.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MAX_D1_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23849\,
            lcout => \il_max_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47995\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_0_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24296\,
            in1 => \N__24469\,
            in2 => \_gnd_net_\,
            in3 => \N__24176\,
            lcout => \pwm_generator_inst.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_9_7_0_\,
            carryout => \pwm_generator_inst.counter_cry_0\,
            clk => \N__47981\,
            ce => 'H',
            sr => \N__47310\
        );

    \pwm_generator_inst.counter_1_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24292\,
            in1 => \N__24388\,
            in2 => \_gnd_net_\,
            in3 => \N__24173\,
            lcout => \pwm_generator_inst.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_0\,
            carryout => \pwm_generator_inst.counter_cry_1\,
            clk => \N__47981\,
            ce => 'H',
            sr => \N__47310\
        );

    \pwm_generator_inst.counter_2_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24297\,
            in1 => \N__24490\,
            in2 => \_gnd_net_\,
            in3 => \N__24170\,
            lcout => \pwm_generator_inst.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_1\,
            carryout => \pwm_generator_inst.counter_cry_2\,
            clk => \N__47981\,
            ce => 'H',
            sr => \N__47310\
        );

    \pwm_generator_inst.counter_3_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24293\,
            in1 => \N__24409\,
            in2 => \_gnd_net_\,
            in3 => \N__24167\,
            lcout => \pwm_generator_inst.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_2\,
            carryout => \pwm_generator_inst.counter_cry_3\,
            clk => \N__47981\,
            ce => 'H',
            sr => \N__47310\
        );

    \pwm_generator_inst.counter_4_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24298\,
            in1 => \N__24364\,
            in2 => \_gnd_net_\,
            in3 => \N__24164\,
            lcout => \pwm_generator_inst.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_3\,
            carryout => \pwm_generator_inst.counter_cry_4\,
            clk => \N__47981\,
            ce => 'H',
            sr => \N__47310\
        );

    \pwm_generator_inst.counter_5_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24294\,
            in1 => \N__24316\,
            in2 => \_gnd_net_\,
            in3 => \N__24161\,
            lcout => \pwm_generator_inst.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_4\,
            carryout => \pwm_generator_inst.counter_cry_5\,
            clk => \N__47981\,
            ce => 'H',
            sr => \N__47310\
        );

    \pwm_generator_inst.counter_6_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24299\,
            in1 => \N__24340\,
            in2 => \_gnd_net_\,
            in3 => \N__24158\,
            lcout => \pwm_generator_inst.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_5\,
            carryout => \pwm_generator_inst.counter_cry_6\,
            clk => \N__47981\,
            ce => 'H',
            sr => \N__47310\
        );

    \pwm_generator_inst.counter_7_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24295\,
            in1 => \N__24217\,
            in2 => \_gnd_net_\,
            in3 => \N__24155\,
            lcout => \pwm_generator_inst.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_6\,
            carryout => \pwm_generator_inst.counter_cry_7\,
            clk => \N__47981\,
            ce => 'H',
            sr => \N__47310\
        );

    \pwm_generator_inst.counter_8_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24291\,
            in1 => \N__24236\,
            in2 => \_gnd_net_\,
            in3 => \N__24152\,
            lcout => \pwm_generator_inst.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_9_8_0_\,
            carryout => \pwm_generator_inst.counter_cry_8\,
            clk => \N__47972\,
            ce => 'H',
            sr => \N__47316\
        );

    \pwm_generator_inst.counter_9_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__24256\,
            in1 => \N__24290\,
            in2 => \_gnd_net_\,
            in3 => \N__24413\,
            lcout => \pwm_generator_inst.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47972\,
            ce => 'H',
            sr => \N__47316\
        );

    \pwm_generator_inst.counter_RNIBO26_1_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000101"
        )
    port map (
            in0 => \N__24410\,
            in1 => \N__24389\,
            in2 => \N__24368\,
            in3 => \N__24449\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlt9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIFA6C_5_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__24197\,
            in1 => \N__24344\,
            in2 => \N__24323\,
            in3 => \N__24320\,
            lcout => \pwm_generator_inst.un1_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIVDL3_9_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__24257\,
            in1 => \N__24234\,
            in2 => \_gnd_net_\,
            in3 => \N__24218\,
            lcout => \pwm_generator_inst.un1_counterlto9_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI3MVS6_31_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101010101"
        )
    port map (
            in0 => \N__33069\,
            in1 => \N__30104\,
            in2 => \_gnd_net_\,
            in3 => \N__30075\,
            lcout => \current_shift_inst.PI_CTRL.N_79\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIB98M_0_10_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29615\,
            in1 => \N__28901\,
            in2 => \N__28219\,
            in3 => \N__29217\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI775B_18_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33011\,
            in2 => \_gnd_net_\,
            in3 => \N__28655\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29693\,
            in1 => \N__32589\,
            in2 => \N__29568\,
            in3 => \N__28056\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI50UD2_10_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24497\,
            in1 => \N__24191\,
            in2 => \N__24185\,
            in3 => \N__24182\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28979\,
            in1 => \N__29046\,
            in2 => \N__28837\,
            in3 => \N__28133\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNISQD2_0_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24491\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24470\,
            lcout => \pwm_generator_inst.un1_counterlto2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30347\,
            in1 => \N__30392\,
            in2 => \N__29100\,
            in3 => \N__29354\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIO0BU3_18_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__33062\,
            in1 => \N__28659\,
            in2 => \N__24443\,
            in3 => \N__24440\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29355\,
            in1 => \N__30348\,
            in2 => \N__30402\,
            in3 => \N__29093\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29418\,
            in1 => \N__28736\,
            in2 => \N__29292\,
            in3 => \N__28583\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIC35V7_17_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24434\,
            in1 => \N__24428\,
            in2 => \N__24422\,
            in3 => \N__24419\,
            lcout => \current_shift_inst.PI_CTRL.N_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_17_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011111111"
        )
    port map (
            in0 => \N__33063\,
            in1 => \N__32826\,
            in2 => \N__28688\,
            in3 => \N__32703\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47945\,
            ce => \N__32549\,
            sr => \N__47353\
        );

    \current_shift_inst.PI_CTRL.integrator_30_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011111111"
        )
    port map (
            in0 => \N__33066\,
            in1 => \N__32835\,
            in2 => \N__29528\,
            in3 => \N__32708\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47945\,
            ce => \N__32549\,
            sr => \N__47353\
        );

    \current_shift_inst.PI_CTRL.integrator_20_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011111111"
        )
    port map (
            in0 => \N__33064\,
            in1 => \N__32830\,
            in2 => \N__29384\,
            in3 => \N__32705\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47945\,
            ce => \N__32549\,
            sr => \N__47353\
        );

    \current_shift_inst.PI_CTRL.integrator_22_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110111010101"
        )
    port map (
            in0 => \N__32706\,
            in1 => \N__29234\,
            in2 => \N__32864\,
            in3 => \N__33068\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47945\,
            ce => \N__32549\,
            sr => \N__47353\
        );

    \current_shift_inst.PI_CTRL.integrator_23_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011111111"
        )
    port map (
            in0 => \N__33065\,
            in1 => \N__32834\,
            in2 => \N__29162\,
            in3 => \N__32707\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47945\,
            ce => \N__32549\,
            sr => \N__47353\
        );

    \current_shift_inst.PI_CTRL.integrator_19_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110111010101"
        )
    port map (
            in0 => \N__32704\,
            in1 => \N__28529\,
            in2 => \N__32863\,
            in3 => \N__33067\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47945\,
            ce => \N__32549\,
            sr => \N__47353\
        );

    \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CRY_0_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27142\,
            in2 => \N__27146\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_13_0_\,
            carryout => \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_0_c_inv_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24554\,
            in2 => \N__26510\,
            in3 => \N__29972\,
            lcout => \current_shift_inst.z_i_0_31\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CO\,
            carryout => \current_shift_inst.un38_control_input_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_1_c_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26488\,
            in2 => \N__24548\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_0\,
            carryout => \current_shift_inst.un38_control_input_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_2_c_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26455\,
            in2 => \N__24533\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_1\,
            carryout => \current_shift_inst.un38_control_input_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_3_c_inv_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24518\,
            in1 => \N__26420\,
            in2 => \N__24506\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un38_control_input_0_cry_3_c_invZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_2\,
            carryout => \current_shift_inst.un38_control_input_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_4_c_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25433\,
            in2 => \N__25459\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_3\,
            carryout => \current_shift_inst.un38_control_input_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_5_c_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25568\,
            in2 => \N__25427\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_4\,
            carryout => \current_shift_inst.un38_control_input_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_5_c_RNI7HN13_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25415\,
            in2 => \N__25370\,
            in3 => \N__24602\,
            lcout => \current_shift_inst.control_input_1_axb_0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_5\,
            carryout => \current_shift_inst.un38_control_input_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_6_c_RNIHVR13_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25511\,
            in2 => \N__25469\,
            in3 => \N__24593\,
            lcout => \current_shift_inst.control_input_1_axb_1\,
            ltout => OPEN,
            carryin => \bfn_9_14_0_\,
            carryout => \current_shift_inst.un38_control_input_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_7_c_RNIRD023_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25847\,
            in2 => \N__25523\,
            in3 => \N__24584\,
            lcout => \current_shift_inst.control_input_1_axb_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_7\,
            carryout => \current_shift_inst.un38_control_input_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_8_c_RNIC9753_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25706\,
            in2 => \N__25397\,
            in3 => \N__24575\,
            lcout => \current_shift_inst.control_input_1_axb_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_8\,
            carryout => \current_shift_inst.un38_control_input_0_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_9_c_RNII9PR2_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25898\,
            in2 => \N__25379\,
            in3 => \N__24566\,
            lcout => \current_shift_inst.control_input_1_axb_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_9\,
            carryout => \current_shift_inst.un38_control_input_0_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_10_c_RNIV96V1_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25949\,
            in2 => \N__25550\,
            in3 => \N__24557\,
            lcout => \current_shift_inst.control_input_1_axb_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_10\,
            carryout => \current_shift_inst.un38_control_input_0_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_11_c_RNI9OAV1_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30725\,
            in2 => \N__25406\,
            in3 => \N__24707\,
            lcout => \current_shift_inst.control_input_1_axb_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_11\,
            carryout => \current_shift_inst.un38_control_input_0_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_12_c_RNIJ6FV1_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24704\,
            in2 => \N__25388\,
            in3 => \N__24686\,
            lcout => \current_shift_inst.control_input_1_axb_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_12\,
            carryout => \current_shift_inst.un38_control_input_0_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_13_c_RNITKJV1_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24683\,
            in2 => \N__25652\,
            in3 => \N__24665\,
            lcout => \current_shift_inst.control_input_1_axb_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_13\,
            carryout => \current_shift_inst.un38_control_input_0_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_14_c_RNI73OV1_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25529\,
            in2 => \N__25793\,
            in3 => \N__24656\,
            lcout => \current_shift_inst.control_input_1_axb_9\,
            ltout => OPEN,
            carryin => \bfn_9_15_0_\,
            carryout => \current_shift_inst.un38_control_input_0_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_15_c_RNIHHSV1_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26108\,
            in2 => \N__25559\,
            in3 => \N__24647\,
            lcout => \current_shift_inst.control_input_1_axb_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_15\,
            carryout => \current_shift_inst.un38_control_input_0_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_16_c_RNIRV002_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26156\,
            in2 => \N__25538\,
            in3 => \N__24638\,
            lcout => \current_shift_inst.control_input_1_axb_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_16\,
            carryout => \current_shift_inst.un38_control_input_0_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_17_c_RNI5E502_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25955\,
            in2 => \N__26258\,
            in3 => \N__24629\,
            lcout => \current_shift_inst.control_input_1_axb_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_17\,
            carryout => \current_shift_inst.un38_control_input_0_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_18_c_RNI6KA02_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25700\,
            in2 => \N__26267\,
            in3 => \N__24620\,
            lcout => \current_shift_inst.control_input_1_axb_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_18\,
            carryout => \current_shift_inst.un38_control_input_0_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_19_c_RNICO912_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26201\,
            in2 => \N__25943\,
            in3 => \N__24611\,
            lcout => \current_shift_inst.control_input_1_axb_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_19\,
            carryout => \current_shift_inst.un38_control_input_0_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_20_c_RNI92P32_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26030\,
            in2 => \N__26249\,
            in3 => \N__24833\,
            lcout => \current_shift_inst.control_input_1_axb_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_20\,
            carryout => \current_shift_inst.un38_control_input_0_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_21_c_RNIJGT32_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25694\,
            in2 => \N__26276\,
            in3 => \N__24824\,
            lcout => \current_shift_inst.control_input_1_axb_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_21\,
            carryout => \current_shift_inst.un38_control_input_0_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_22_c_RNITU142_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30527\,
            in2 => \N__30434\,
            in3 => \N__24815\,
            lcout => \current_shift_inst.control_input_1_axb_17\,
            ltout => OPEN,
            carryin => \bfn_9_16_0_\,
            carryout => \current_shift_inst.un38_control_input_0_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_23_c_RNI7D642_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24812\,
            in2 => \N__24803\,
            in3 => \N__24785\,
            lcout => \current_shift_inst.control_input_1_axb_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_23\,
            carryout => \current_shift_inst.un38_control_input_0_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_24_c_RNIHRA42_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31112\,
            in2 => \N__30713\,
            in3 => \N__24776\,
            lcout => \current_shift_inst.control_input_1_axb_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_24\,
            carryout => \current_shift_inst.un38_control_input_0_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_25_c_RNIR9F42_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24773\,
            in2 => \N__24764\,
            in3 => \N__24746\,
            lcout => \current_shift_inst.control_input_1_axb_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_25\,
            carryout => \current_shift_inst.un38_control_input_0_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_26_c_RNI5OJ42_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30614\,
            in2 => \N__31298\,
            in3 => \N__24737\,
            lcout => \current_shift_inst.control_input_1_axb_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_26\,
            carryout => \current_shift_inst.un38_control_input_0_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_27_c_RNIF6O42_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26978\,
            in2 => \N__24734\,
            in3 => \N__24716\,
            lcout => \current_shift_inst.control_input_1_axb_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_27\,
            carryout => \current_shift_inst.un38_control_input_0_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_28_c_RNIGCT42_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25070\,
            in2 => \N__25061\,
            in3 => \N__25043\,
            lcout => \current_shift_inst.control_input_1_axb_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_28\,
            carryout => \current_shift_inst.un38_control_input_0_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_29_c_RNIMGS52_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25040\,
            in2 => \N__25028\,
            in3 => \N__24995\,
            lcout => \current_shift_inst.control_input_1_axb_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_29\,
            carryout => \current_shift_inst.un38_control_input_0_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_25_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24992\,
            in2 => \N__24980\,
            in3 => \N__24971\,
            lcout => \current_shift_inst.control_inputZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47908\,
            ce => \N__24967\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_0_c_inv_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26500\,
            in2 => \N__24923\,
            in3 => \N__29768\,
            lcout => \G_406\,
            ltout => OPEN,
            carryin => \bfn_9_18_0_\,
            carryout => \current_shift_inst.z_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_1_c_inv_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26475\,
            in2 => \N__24875\,
            in3 => \N__24914\,
            lcout => \G_405\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_0\,
            carryout => \current_shift_inst.z_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_2_c_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24866\,
            in2 => \N__26448\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_1\,
            carryout => \current_shift_inst.z_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_3_c_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26413\,
            in2 => \N__24857\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_2\,
            carryout => \current_shift_inst.z_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_4_c_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26388\,
            in2 => \N__24848\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_3\,
            carryout => \current_shift_inst.z_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_5_c_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25124\,
            in2 => \N__26366\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_4\,
            carryout => \current_shift_inst.z_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_6_c_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25118\,
            in2 => \N__26336\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_5\,
            carryout => \current_shift_inst.z_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_7_c_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25112\,
            in2 => \N__26303\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_6\,
            carryout => \current_shift_inst.z_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_8_c_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25106\,
            in2 => \N__26765\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_19_0_\,
            carryout => \current_shift_inst.z_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_9_c_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25097\,
            in2 => \N__26720\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_8\,
            carryout => \current_shift_inst.z_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_10_c_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25091\,
            in2 => \N__26681\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_9\,
            carryout => \current_shift_inst.z_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_11_c_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25085\,
            in2 => \N__30797\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_10\,
            carryout => \current_shift_inst.z_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_12_c_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30827\,
            in2 => \N__25079\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_11\,
            carryout => \current_shift_inst.z_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_13_c_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25184\,
            in2 => \N__26634\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_12\,
            carryout => \current_shift_inst.z_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_14_c_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25178\,
            in2 => \N__26597\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_13\,
            carryout => \current_shift_inst.z_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_15_c_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26556\,
            in2 => \N__25172\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_14\,
            carryout => \current_shift_inst.z_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_16_c_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26524\,
            in2 => \N__25163\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_20_0_\,
            carryout => \current_shift_inst.z_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_17_c_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25148\,
            in2 => \N__26951\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_16\,
            carryout => \current_shift_inst.z_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_18_c_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25142\,
            in2 => \N__26912\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_17\,
            carryout => \current_shift_inst.z_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_19_c_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25136\,
            in2 => \N__26868\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_18\,
            carryout => \current_shift_inst.z_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_20_c_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25130\,
            in2 => \N__26840\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_19\,
            carryout => \current_shift_inst.z_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_21_c_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26799\,
            in2 => \N__25247\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_20\,
            carryout => \current_shift_inst.z_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_22_c_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25238\,
            in2 => \N__30459\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_21\,
            carryout => \current_shift_inst.z_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_23_c_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25232\,
            in2 => \N__30552\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_22\,
            carryout => \current_shift_inst.z_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_24_c_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25226\,
            in2 => \N__31178\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_21_0_\,
            carryout => \current_shift_inst.z_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_25_c_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25217\,
            in2 => \N__31220\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_24\,
            carryout => \current_shift_inst.z_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_26_c_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25211\,
            in2 => \N__31323\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_25\,
            carryout => \current_shift_inst.z_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_27_c_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25205\,
            in2 => \N__30644\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_26\,
            carryout => \current_shift_inst.z_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_28_c_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25199\,
            in2 => \N__27001\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_27\,
            carryout => \current_shift_inst.z_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_29_c_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27160\,
            in2 => \N__25193\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_28\,
            carryout => \current_shift_inst.z_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_30_c_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27055\,
            in2 => \N__25316\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_29\,
            carryout => \current_shift_inst.z_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_s_31_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__27135\,
            in1 => \N__25307\,
            in2 => \N__25301\,
            in3 => \N__25277\,
            lcout => \current_shift_inst.z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.stop_timer_s1_RNO_0_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30198\,
            in1 => \N__30278\,
            in2 => \N__27614\,
            in3 => \N__30245\,
            lcout => \current_shift_inst.stop_timer_s1_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_LC_9_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__27602\,
            in1 => \N__27568\,
            in2 => \_gnd_net_\,
            in3 => \N__27541\,
            lcout => \current_shift_inst.timer_s1.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47868\,
            ce => 'H',
            sr => \N__47416\
        );

    \current_shift_inst.meas_state_0_LC_9_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111111001100"
        )
    port map (
            in0 => \N__30202\,
            in1 => \N__30279\,
            in2 => \N__27612\,
            in3 => \N__30244\,
            lcout => \current_shift_inst.meas_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47868\,
            ce => 'H',
            sr => \N__47416\
        );

    \current_shift_inst.start_timer_phase_LC_9_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100101010"
        )
    port map (
            in0 => \N__25265\,
            in1 => \N__30281\,
            in2 => \N__32306\,
            in3 => \N__30246\,
            lcout => \current_shift_inst.start_timer_phaseZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47862\,
            ce => \N__35837\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.start_timer_s1_LC_9_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001111110000"
        )
    port map (
            in0 => \N__30194\,
            in1 => \N__30280\,
            in2 => \N__27613\,
            in3 => \N__30247\,
            lcout => \current_shift_inst.start_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47862\,
            ce => \N__35837\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.stop_timer_s1_LC_9_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111001100"
        )
    port map (
            in0 => \N__30248\,
            in1 => \N__25274\,
            in2 => \N__30289\,
            in3 => \N__27542\,
            lcout => \current_shift_inst.stop_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47862\,
            ce => \N__35837\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.running_LC_9_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__25264\,
            in1 => \N__27473\,
            in2 => \_gnd_net_\,
            in3 => \N__27450\,
            lcout => \current_shift_inst.timer_phase.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47857\,
            ce => 'H',
            sr => \N__47422\
        );

    \SB_DFF_inst_PH1_MAX_D2_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25358\,
            lcout => \il_max_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47963\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_6_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28483\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47955\,
            ce => \N__32550\,
            sr => \N__47311\
        );

    \current_shift_inst.PI_CTRL.integrator_7_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000100000000"
        )
    port map (
            in0 => \N__33074\,
            in1 => \N__32881\,
            in2 => \N__28385\,
            in3 => \N__32638\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47955\,
            ce => \N__32550\,
            sr => \N__47311\
        );

    \current_shift_inst.PI_CTRL.prop_term_9_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28265\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47955\,
            ce => \N__32550\,
            sr => \N__47311\
        );

    \current_shift_inst.PI_CTRL.integrator_18_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011111111"
        )
    port map (
            in0 => \N__33036\,
            in1 => \N__32838\,
            in2 => \N__28607\,
            in3 => \N__32656\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47946\,
            ce => \N__32553\,
            sr => \N__47317\
        );

    \current_shift_inst.PI_CTRL.integrator_3_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000111110011"
        )
    port map (
            in0 => \N__30117\,
            in1 => \N__32842\,
            in2 => \N__27773\,
            in3 => \N__30074\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47946\,
            ce => \N__32553\,
            sr => \N__47317\
        );

    \current_shift_inst.PI_CTRL.integrator_13_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011111111"
        )
    port map (
            in0 => \N__33034\,
            in1 => \N__32836\,
            in2 => \N__28997\,
            in3 => \N__32653\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47946\,
            ce => \N__32553\,
            sr => \N__47317\
        );

    \current_shift_inst.PI_CTRL.integrator_15_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110111010101"
        )
    port map (
            in0 => \N__32655\,
            in1 => \N__28850\,
            in2 => \N__33073\,
            in3 => \N__32839\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47946\,
            ce => \N__32553\,
            sr => \N__47317\
        );

    \current_shift_inst.PI_CTRL.integrator_14_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011111111"
        )
    port map (
            in0 => \N__33035\,
            in1 => \N__32837\,
            in2 => \N__28925\,
            in3 => \N__32654\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47946\,
            ce => \N__32553\,
            sr => \N__47317\
        );

    \current_shift_inst.PI_CTRL.integrator_1_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__30116\,
            in1 => \N__32840\,
            in2 => \N__27875\,
            in3 => \N__30073\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47946\,
            ce => \N__32553\,
            sr => \N__47317\
        );

    \current_shift_inst.PI_CTRL.integrator_29_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010111010101"
        )
    port map (
            in0 => \N__32657\,
            in1 => \N__33037\,
            in2 => \N__29594\,
            in3 => \N__32841\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47946\,
            ce => \N__32553\,
            sr => \N__47317\
        );

    \current_shift_inst.PI_CTRL.integrator_6_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100010001010"
        )
    port map (
            in0 => \N__32714\,
            in1 => \N__28457\,
            in2 => \N__32861\,
            in3 => \N__33081\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47937\,
            ce => \N__32552\,
            sr => \N__47323\
        );

    \current_shift_inst.PI_CTRL.integrator_11_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011111111"
        )
    port map (
            in0 => \N__33076\,
            in1 => \N__32811\,
            in2 => \N__28082\,
            in3 => \N__32710\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47937\,
            ce => \N__32552\,
            sr => \N__47323\
        );

    \current_shift_inst.PI_CTRL.integrator_12_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110111010101"
        )
    port map (
            in0 => \N__32711\,
            in1 => \N__28004\,
            in2 => \N__32859\,
            in3 => \N__33079\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47937\,
            ce => \N__32552\,
            sr => \N__47323\
        );

    \current_shift_inst.PI_CTRL.integrator_9_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000100000000"
        )
    port map (
            in0 => \N__33078\,
            in1 => \N__32825\,
            in2 => \N__28232\,
            in3 => \N__32716\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47937\,
            ce => \N__32552\,
            sr => \N__47323\
        );

    \current_shift_inst.PI_CTRL.integrator_26_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110111010101"
        )
    port map (
            in0 => \N__32713\,
            in1 => \N__29072\,
            in2 => \N__32860\,
            in3 => \N__33080\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47937\,
            ce => \N__32552\,
            sr => \N__47323\
        );

    \current_shift_inst.PI_CTRL.integrator_21_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011111111"
        )
    port map (
            in0 => \N__33077\,
            in1 => \N__32815\,
            in2 => \N__29309\,
            in3 => \N__32712\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47937\,
            ce => \N__32552\,
            sr => \N__47323\
        );

    \current_shift_inst.PI_CTRL.integrator_8_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100010001010"
        )
    port map (
            in0 => \N__32715\,
            in1 => \N__28316\,
            in2 => \N__32862\,
            in3 => \N__33082\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47937\,
            ce => \N__32552\,
            sr => \N__47323\
        );

    \current_shift_inst.PI_CTRL.integrator_10_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011111111"
        )
    port map (
            in0 => \N__33075\,
            in1 => \N__32810\,
            in2 => \N__28157\,
            in3 => \N__32709\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47937\,
            ce => \N__32552\,
            sr => \N__47323\
        );

    \current_shift_inst.timer_s1.running_RNIUKI8_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27575\,
            lcout => \current_shift_inst.timer_s1.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_4_c_RNO_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \N__25460\,
            in1 => \_gnd_net_\,
            in2 => \N__25612\,
            in3 => \N__26397\,
            lcout => \current_shift_inst.un38_control_input_0_cry_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_5_c_RNO_0_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__26398\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25605\,
            lcout => \current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_1_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__41279\,
            in1 => \N__35303\,
            in2 => \N__40730\,
            in3 => \N__40831\,
            lcout => measured_delay_hc_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47928\,
            ce => 'H',
            sr => \N__47335\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQKU1_5_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__25643\,
            in1 => \N__25503\,
            in2 => \N__26372\,
            in3 => \N__26337\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIVQKU1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILORI_11_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30890\,
            in2 => \_gnd_net_\,
            in3 => \N__30801\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNILORI_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIN7DV_8_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25742\,
            in2 => \_gnd_net_\,
            in3 => \N__26771\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIN7DV_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOSSI_12_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30764\,
            in2 => \_gnd_net_\,
            in3 => \N__30843\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIOSSI_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1PG21_9_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__25770\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26730\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI1PG21_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIER9V_5_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25642\,
            in2 => \_gnd_net_\,
            in3 => \N__26367\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIER9V_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIP5T51_13_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__26647\,
            in1 => \N__25836\,
            in2 => \N__25688\,
            in3 => \N__26599\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIP5T51_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_5_c_RNO_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__26399\,
            in1 => \N__25641\,
            in2 => \N__25613\,
            in3 => \N__26368\,
            lcout => \current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5M161_15_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__26566\,
            in1 => \N__26194\,
            in2 => \N__26150\,
            in3 => \N__26538\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5M161_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIIKQI_10_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25933\,
            in2 => \_gnd_net_\,
            in3 => \N__26689\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIIKQI_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4D1J_16_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26195\,
            in2 => \_gnd_net_\,
            in3 => \N__26539\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI4D1J_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVDV51_14_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__25841\,
            in1 => \N__26146\,
            in2 => \N__26606\,
            in3 => \N__26565\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIVDV51_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIK3CV_7_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__26304\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25890\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIK3CV_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI53NU1_6_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__25505\,
            in1 => \N__25891\,
            in2 => \N__26342\,
            in3 => \N__26305\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI53NU1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHVAV_6_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25504\,
            in2 => \_gnd_net_\,
            in3 => \N__26338\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIHVAV_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7DM51_10_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__25934\,
            in1 => \N__30805\,
            in2 => \N__26693\,
            in3 => \N__30886\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI7DM51_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4H5J_19_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__26878\,
            in1 => \_gnd_net_\,
            in2 => \N__26239\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI4H5J_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJDBL1_10_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__26734\,
            in1 => \N__25932\,
            in2 => \N__25781\,
            in3 => \N__26688\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJDBL1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBBPU1_7_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__25892\,
            in1 => \N__26769\,
            in2 => \N__26309\,
            in3 => \N__25740\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIBBPU1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU4VI_14_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25837\,
            in2 => \_gnd_net_\,
            in3 => \N__26598\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIU4VI_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIO0U12_8_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110100101"
        )
    port map (
            in0 => \N__25777\,
            in1 => \N__25741\,
            in2 => \N__26735\,
            in3 => \N__26770\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIO0U12_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIE6961_18_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__25989\,
            in1 => \N__26877\,
            in2 => \N__26921\,
            in3 => \N__26232\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIE6961_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJ3381_21_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \N__26813\,
            in1 => \N__26069\,
            in2 => \N__30515\,
            in3 => \N__30465\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJ3381_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOV0K_21_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__26068\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26812\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIOV0K_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAL3J_18_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__26913\,
            in1 => \_gnd_net_\,
            in2 => \N__25994\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIAL3J_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7H2J_17_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26024\,
            in3 => \N__26952\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI7H2J_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILRVJ_20_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26102\,
            in3 => \N__26841\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNILRVJ_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPC571_19_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100110011001"
        )
    port map (
            in0 => \N__26842\,
            in1 => \N__26097\,
            in2 => \N__26885\,
            in3 => \N__26240\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPC571_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBU361_16_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001111000011"
        )
    port map (
            in0 => \N__26540\,
            in1 => \N__26019\,
            in2 => \N__26959\,
            in3 => \N__26188\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIBU361_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI190J_15_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__26140\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26567\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI190J_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDR081_20_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__26101\,
            in1 => \N__26067\,
            in2 => \N__26846\,
            in3 => \N__26806\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIDR081_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIH6661_17_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__26023\,
            in1 => \N__25990\,
            in2 => \N__26960\,
            in3 => \N__26914\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIH6661_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_RNI48NB_31_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29735\,
            in2 => \N__29767\,
            in3 => \N__29763\,
            lcout => \current_shift_inst.un38_control_input_0\,
            ltout => OPEN,
            carryin => \bfn_10_17_0_\,
            carryout => \current_shift_inst.un4_control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_1_c_RNIJF2G_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29723\,
            in2 => \_gnd_net_\,
            in3 => \N__26459\,
            lcout => \current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_1\,
            carryout => \current_shift_inst.un4_control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_2_c_RNILI3G_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29711\,
            in2 => \_gnd_net_\,
            in3 => \N__26423\,
            lcout => \current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_2\,
            carryout => \current_shift_inst.un4_control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_3_c_RNINL4G_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29834\,
            in2 => \_gnd_net_\,
            in3 => \N__26402\,
            lcout => \current_shift_inst.un4_control_input_cry_3_c_RNINL4GZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_3\,
            carryout => \current_shift_inst.un4_control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_4_c_RNIPO5G_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29828\,
            in2 => \_gnd_net_\,
            in3 => \N__26375\,
            lcout => \current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_4\,
            carryout => \current_shift_inst.un4_control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_5_c_RNIRR6G_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29822\,
            in2 => \_gnd_net_\,
            in3 => \N__26345\,
            lcout => \current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_5\,
            carryout => \current_shift_inst.un4_control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_6_c_RNITU7G_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29816\,
            in3 => \N__26312\,
            lcout => \current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_6\,
            carryout => \current_shift_inst.un4_control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_7_c_RNIV19G_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29807\,
            in3 => \N__26279\,
            lcout => \current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_7\,
            carryout => \current_shift_inst.un4_control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_8_c_RNI15AG_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29786\,
            in2 => \_gnd_net_\,
            in3 => \N__26738\,
            lcout => \current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0\,
            ltout => OPEN,
            carryin => \bfn_10_18_0_\,
            carryout => \current_shift_inst.un4_control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_9_c_RNIALDJ_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29780\,
            in2 => \_gnd_net_\,
            in3 => \N__26696\,
            lcout => \current_shift_inst.un4_control_input_cry_9_c_RNIALDJZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_9\,
            carryout => \current_shift_inst.un4_control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_10_c_RNIJLTG_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29774\,
            in2 => \_gnd_net_\,
            in3 => \N__26657\,
            lcout => \current_shift_inst.un4_control_input_cry_10_c_RNIJLTGZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_10\,
            carryout => \current_shift_inst.un4_control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_11_c_RNILOUG_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29888\,
            in2 => \_gnd_net_\,
            in3 => \N__26654\,
            lcout => \current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_11\,
            carryout => \current_shift_inst.un4_control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_12_c_RNINRVG_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29798\,
            in2 => \_gnd_net_\,
            in3 => \N__26651\,
            lcout => \current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_12\,
            carryout => \current_shift_inst.un4_control_input_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_13_c_RNIPU0H_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29717\,
            in2 => \_gnd_net_\,
            in3 => \N__26609\,
            lcout => \current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_13\,
            carryout => \current_shift_inst.un4_control_input_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_14_c_RNIR12H_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29792\,
            in2 => \_gnd_net_\,
            in3 => \N__26570\,
            lcout => \current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_14\,
            carryout => \current_shift_inst.un4_control_input_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_15_c_RNIT43H_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29882\,
            in2 => \_gnd_net_\,
            in3 => \N__26543\,
            lcout => \current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_15\,
            carryout => \current_shift_inst.un4_control_input_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_16_c_RNIV74H_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29993\,
            in2 => \_gnd_net_\,
            in3 => \N__26513\,
            lcout => \current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0\,
            ltout => OPEN,
            carryin => \bfn_10_19_0_\,
            carryout => \current_shift_inst.un4_control_input_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_17_c_RNI1B5H_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29870\,
            in2 => \_gnd_net_\,
            in3 => \N__26924\,
            lcout => \current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_17\,
            carryout => \current_shift_inst.un4_control_input_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_18_c_RNI3E6H_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29858\,
            in2 => \_gnd_net_\,
            in3 => \N__26888\,
            lcout => \current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_18\,
            carryout => \current_shift_inst.un4_control_input_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_19_c_RNIS88H_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29876\,
            in2 => \_gnd_net_\,
            in3 => \N__26849\,
            lcout => \current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_19\,
            carryout => \current_shift_inst.un4_control_input_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_20_c_RNILQ1I_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29987\,
            in2 => \_gnd_net_\,
            in3 => \N__26816\,
            lcout => \current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_20\,
            carryout => \current_shift_inst.un4_control_input_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_21_c_RNINT2I_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29846\,
            in2 => \_gnd_net_\,
            in3 => \N__26786\,
            lcout => \current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_21\,
            carryout => \current_shift_inst.un4_control_input_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_22_c_RNIP04I_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29864\,
            in2 => \_gnd_net_\,
            in3 => \N__26783\,
            lcout => \current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_22\,
            carryout => \current_shift_inst.un4_control_input_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_23_c_RNIR35I_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29840\,
            in2 => \_gnd_net_\,
            in3 => \N__26780\,
            lcout => \current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_23\,
            carryout => \current_shift_inst.un4_control_input_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_24_c_RNIT66I_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29852\,
            in2 => \_gnd_net_\,
            in3 => \N__26777\,
            lcout => \current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0\,
            ltout => OPEN,
            carryin => \bfn_10_20_0_\,
            carryout => \current_shift_inst.un4_control_input_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_25_c_RNIV97I_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29978\,
            in2 => \_gnd_net_\,
            in3 => \N__26774\,
            lcout => \current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_25\,
            carryout => \current_shift_inst.un4_control_input_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_26_c_RNI1D8I_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29915\,
            in2 => \_gnd_net_\,
            in3 => \N__27179\,
            lcout => \current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_26\,
            carryout => \current_shift_inst.un4_control_input_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_27_c_RNI3G9I_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29897\,
            in2 => \_gnd_net_\,
            in3 => \N__27176\,
            lcout => \current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_27\,
            carryout => \current_shift_inst.un4_control_input_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_28_c_RNI5JAI_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29906\,
            in2 => \_gnd_net_\,
            in3 => \N__27173\,
            lcout => \current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_28\,
            carryout => \current_shift_inst.un4_control_input_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_29_c_RNIUDCI_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29924\,
            in2 => \_gnd_net_\,
            in3 => \N__27149\,
            lcout => \current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_29\,
            carryout => \current_shift_inst.un4_control_input_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_30_c_RNINV5J_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27134\,
            in2 => \_gnd_net_\,
            in3 => \N__27068\,
            lcout => \current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNINKG81_27_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__30697\,
            in1 => \N__27044\,
            in2 => \N__30655\,
            in3 => \N__27000\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNINKG81_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.counter_0_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27335\,
            in1 => \N__31086\,
            in2 => \_gnd_net_\,
            in3 => \N__26966\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_10_21_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_0\,
            clk => \N__47877\,
            ce => \N__27517\,
            sr => \N__47399\
        );

    \current_shift_inst.timer_s1.counter_1_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27330\,
            in1 => \N__31047\,
            in2 => \_gnd_net_\,
            in3 => \N__26963\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_0\,
            carryout => \current_shift_inst.timer_s1.counter_cry_1\,
            clk => \N__47877\,
            ce => \N__27517\,
            sr => \N__47399\
        );

    \current_shift_inst.timer_s1.counter_2_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27336\,
            in1 => \N__31017\,
            in2 => \_gnd_net_\,
            in3 => \N__27206\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_1\,
            carryout => \current_shift_inst.timer_s1.counter_cry_2\,
            clk => \N__47877\,
            ce => \N__27517\,
            sr => \N__47399\
        );

    \current_shift_inst.timer_s1.counter_3_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27331\,
            in1 => \N__30987\,
            in2 => \_gnd_net_\,
            in3 => \N__27203\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_2\,
            carryout => \current_shift_inst.timer_s1.counter_cry_3\,
            clk => \N__47877\,
            ce => \N__27517\,
            sr => \N__47399\
        );

    \current_shift_inst.timer_s1.counter_4_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27337\,
            in1 => \N__30946\,
            in2 => \_gnd_net_\,
            in3 => \N__27200\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_3\,
            carryout => \current_shift_inst.timer_s1.counter_cry_4\,
            clk => \N__47877\,
            ce => \N__27517\,
            sr => \N__47399\
        );

    \current_shift_inst.timer_s1.counter_5_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27332\,
            in1 => \N__30910\,
            in2 => \_gnd_net_\,
            in3 => \N__27197\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_4\,
            carryout => \current_shift_inst.timer_s1.counter_cry_5\,
            clk => \N__47877\,
            ce => \N__27517\,
            sr => \N__47399\
        );

    \current_shift_inst.timer_s1.counter_6_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27334\,
            in1 => \N__31615\,
            in2 => \_gnd_net_\,
            in3 => \N__27194\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_5\,
            carryout => \current_shift_inst.timer_s1.counter_cry_6\,
            clk => \N__47877\,
            ce => \N__27517\,
            sr => \N__47399\
        );

    \current_shift_inst.timer_s1.counter_7_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27333\,
            in1 => \N__31585\,
            in2 => \_gnd_net_\,
            in3 => \N__27191\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_6\,
            carryout => \current_shift_inst.timer_s1.counter_cry_7\,
            clk => \N__47877\,
            ce => \N__27517\,
            sr => \N__47399\
        );

    \current_shift_inst.timer_s1.counter_8_LC_10_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27341\,
            in1 => \N__31551\,
            in2 => \_gnd_net_\,
            in3 => \N__27188\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_10_22_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_8\,
            clk => \N__47870\,
            ce => \N__27518\,
            sr => \N__47403\
        );

    \current_shift_inst.timer_s1.counter_9_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27345\,
            in1 => \N__31509\,
            in2 => \_gnd_net_\,
            in3 => \N__27185\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_8\,
            carryout => \current_shift_inst.timer_s1.counter_cry_9\,
            clk => \N__47870\,
            ce => \N__27518\,
            sr => \N__47403\
        );

    \current_shift_inst.timer_s1.counter_10_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27338\,
            in1 => \N__31470\,
            in2 => \_gnd_net_\,
            in3 => \N__27182\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_9\,
            carryout => \current_shift_inst.timer_s1.counter_cry_10\,
            clk => \N__47870\,
            ce => \N__27518\,
            sr => \N__47403\
        );

    \current_shift_inst.timer_s1.counter_11_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27342\,
            in1 => \N__31434\,
            in2 => \_gnd_net_\,
            in3 => \N__27236\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_10\,
            carryout => \current_shift_inst.timer_s1.counter_cry_11\,
            clk => \N__47870\,
            ce => \N__27518\,
            sr => \N__47403\
        );

    \current_shift_inst.timer_s1.counter_12_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27339\,
            in1 => \N__31396\,
            in2 => \_gnd_net_\,
            in3 => \N__27233\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_11\,
            carryout => \current_shift_inst.timer_s1.counter_cry_12\,
            clk => \N__47870\,
            ce => \N__27518\,
            sr => \N__47403\
        );

    \current_shift_inst.timer_s1.counter_13_LC_10_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27343\,
            in1 => \N__31900\,
            in2 => \_gnd_net_\,
            in3 => \N__27230\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_12\,
            carryout => \current_shift_inst.timer_s1.counter_cry_13\,
            clk => \N__47870\,
            ce => \N__27518\,
            sr => \N__47403\
        );

    \current_shift_inst.timer_s1.counter_14_LC_10_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27340\,
            in1 => \N__31864\,
            in2 => \_gnd_net_\,
            in3 => \N__27227\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_13\,
            carryout => \current_shift_inst.timer_s1.counter_cry_14\,
            clk => \N__47870\,
            ce => \N__27518\,
            sr => \N__47403\
        );

    \current_shift_inst.timer_s1.counter_15_LC_10_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27344\,
            in1 => \N__31828\,
            in2 => \_gnd_net_\,
            in3 => \N__27224\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_14\,
            carryout => \current_shift_inst.timer_s1.counter_cry_15\,
            clk => \N__47870\,
            ce => \N__27518\,
            sr => \N__47403\
        );

    \current_shift_inst.timer_s1.counter_16_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27350\,
            in1 => \N__31797\,
            in2 => \_gnd_net_\,
            in3 => \N__27221\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_10_23_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_16\,
            clk => \N__47864\,
            ce => \N__27507\,
            sr => \N__47406\
        );

    \current_shift_inst.timer_s1.counter_17_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27346\,
            in1 => \N__31758\,
            in2 => \_gnd_net_\,
            in3 => \N__27218\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_16\,
            carryout => \current_shift_inst.timer_s1.counter_cry_17\,
            clk => \N__47864\,
            ce => \N__27507\,
            sr => \N__47406\
        );

    \current_shift_inst.timer_s1.counter_18_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27351\,
            in1 => \N__31719\,
            in2 => \_gnd_net_\,
            in3 => \N__27215\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_17\,
            carryout => \current_shift_inst.timer_s1.counter_cry_18\,
            clk => \N__47864\,
            ce => \N__27507\,
            sr => \N__47406\
        );

    \current_shift_inst.timer_s1.counter_19_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27347\,
            in1 => \N__31683\,
            in2 => \_gnd_net_\,
            in3 => \N__27212\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_18\,
            carryout => \current_shift_inst.timer_s1.counter_cry_19\,
            clk => \N__47864\,
            ce => \N__27507\,
            sr => \N__47406\
        );

    \current_shift_inst.timer_s1.counter_20_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27352\,
            in1 => \N__31648\,
            in2 => \_gnd_net_\,
            in3 => \N__27209\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_19\,
            carryout => \current_shift_inst.timer_s1.counter_cry_20\,
            clk => \N__47864\,
            ce => \N__27507\,
            sr => \N__47406\
        );

    \current_shift_inst.timer_s1.counter_21_LC_10_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27348\,
            in1 => \N__32239\,
            in2 => \_gnd_net_\,
            in3 => \N__27383\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_20\,
            carryout => \current_shift_inst.timer_s1.counter_cry_21\,
            clk => \N__47864\,
            ce => \N__27507\,
            sr => \N__47406\
        );

    \current_shift_inst.timer_s1.counter_22_LC_10_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27353\,
            in1 => \N__32203\,
            in2 => \_gnd_net_\,
            in3 => \N__27380\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_21\,
            carryout => \current_shift_inst.timer_s1.counter_cry_22\,
            clk => \N__47864\,
            ce => \N__27507\,
            sr => \N__47406\
        );

    \current_shift_inst.timer_s1.counter_23_LC_10_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27349\,
            in1 => \N__32167\,
            in2 => \_gnd_net_\,
            in3 => \N__27377\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_22\,
            carryout => \current_shift_inst.timer_s1.counter_cry_23\,
            clk => \N__47864\,
            ce => \N__27507\,
            sr => \N__47406\
        );

    \current_shift_inst.timer_s1.counter_24_LC_10_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27354\,
            in1 => \N__32136\,
            in2 => \_gnd_net_\,
            in3 => \N__27374\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_10_24_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_24\,
            clk => \N__47859\,
            ce => \N__27506\,
            sr => \N__47410\
        );

    \current_shift_inst.timer_s1.counter_25_LC_10_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27358\,
            in1 => \N__32097\,
            in2 => \_gnd_net_\,
            in3 => \N__27371\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_24\,
            carryout => \current_shift_inst.timer_s1.counter_cry_25\,
            clk => \N__47859\,
            ce => \N__27506\,
            sr => \N__47410\
        );

    \current_shift_inst.timer_s1.counter_26_LC_10_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27355\,
            in1 => \N__32040\,
            in2 => \_gnd_net_\,
            in3 => \N__27368\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_25\,
            carryout => \current_shift_inst.timer_s1.counter_cry_26\,
            clk => \N__47859\,
            ce => \N__27506\,
            sr => \N__47410\
        );

    \current_shift_inst.timer_s1.counter_27_LC_10_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27359\,
            in1 => \N__31986\,
            in2 => \_gnd_net_\,
            in3 => \N__27365\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_26\,
            carryout => \current_shift_inst.timer_s1.counter_cry_27\,
            clk => \N__47859\,
            ce => \N__27506\,
            sr => \N__47410\
        );

    \current_shift_inst.timer_s1.counter_28_LC_10_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27356\,
            in1 => \N__32062\,
            in2 => \_gnd_net_\,
            in3 => \N__27362\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_27\,
            carryout => \current_shift_inst.timer_s1.counter_cry_28\,
            clk => \N__47859\,
            ce => \N__27506\,
            sr => \N__47410\
        );

    \current_shift_inst.timer_s1.counter_29_LC_10_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__32008\,
            in1 => \N__27357\,
            in2 => \_gnd_net_\,
            in3 => \N__27239\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47859\,
            ce => \N__27506\,
            sr => \N__47410\
        );

    \current_shift_inst.timer_s1.running_RNIEOIK_LC_10_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__27601\,
            in1 => \N__27567\,
            in2 => \_gnd_net_\,
            in3 => \N__27540\,
            lcout => \current_shift_inst.timer_s1.N_192_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.stop_timer_phase_LC_10_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110100000"
        )
    port map (
            in0 => \N__30285\,
            in1 => \N__30233\,
            in2 => \N__32305\,
            in3 => \N__27451\,
            lcout => \current_shift_inst.stop_timer_phaseZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47853\,
            ce => \N__35836\,
            sr => \_gnd_net_\
        );

    \reset_ibuf_gb_io_RNI79U7_LC_10_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__47460\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => red_c_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.running_RNIC90O_LC_10_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27470\,
            in2 => \_gnd_net_\,
            in3 => \N__27446\,
            lcout => \current_shift_inst.timer_phase.N_188_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MAX_D1_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27410\,
            lcout => \il_max_comp2_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47973\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MIN_D1_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__27398\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_min_comp2_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47964\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_16_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011111111"
        )
    port map (
            in0 => \N__32896\,
            in1 => \N__33007\,
            in2 => \N__28766\,
            in3 => \N__32691\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47947\,
            ce => \N__32551\,
            sr => \N__47304\
        );

    \current_shift_inst.PI_CTRL.integrator_5_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000010100010"
        )
    port map (
            in0 => \N__32694\,
            in1 => \N__33010\,
            in2 => \N__27626\,
            in3 => \N__32899\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47947\,
            ce => \N__32551\,
            sr => \N__47304\
        );

    \current_shift_inst.PI_CTRL.integrator_4_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010111010101"
        )
    port map (
            in0 => \N__32693\,
            in1 => \N__33009\,
            in2 => \N__27704\,
            in3 => \N__32898\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47947\,
            ce => \N__32551\,
            sr => \N__47304\
        );

    \current_shift_inst.PI_CTRL.integrator_28_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011111111"
        )
    port map (
            in0 => \N__32897\,
            in1 => \N__33008\,
            in2 => \N__29654\,
            in3 => \N__32692\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47947\,
            ce => \N__32551\,
            sr => \N__47304\
        );

    \current_shift_inst.PI_CTRL.integrator_0_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__30125\,
            in1 => \N__32895\,
            in2 => \N__27938\,
            in3 => \N__30082\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47947\,
            ce => \N__32551\,
            sr => \N__47304\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_0_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27984\,
            in2 => \N__27964\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.un1_integrator_axb_0\,
            ltout => OPEN,
            carryin => \bfn_11_10_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27918\,
            in2 => \N__27899\,
            in3 => \N__27866\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30024\,
            in2 => \N__27863\,
            in3 => \N__27839\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27832\,
            in2 => \N__27803\,
            in3 => \N__27764\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27744\,
            in2 => \N__27728\,
            in3 => \N__27695\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27677\,
            in2 => \N__27655\,
            in3 => \N__27617\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28505\,
            in2 => \N__28484\,
            in3 => \N__28451\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28423\,
            in2 => \N__28411\,
            in3 => \N__28376\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28361\,
            in2 => \N__28340\,
            in3 => \N__28307\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \bfn_11_11_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28286\,
            in2 => \N__28261\,
            in3 => \N__28223\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28195\,
            in2 => \N__28183\,
            in3 => \N__28148\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28134\,
            in2 => \N__28109\,
            in3 => \N__28073\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28050\,
            in2 => \N__28034\,
            in3 => \N__27995\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29045\,
            in2 => \N__29024\,
            in3 => \N__28988\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28980\,
            in2 => \N__28955\,
            in3 => \N__28913\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28902\,
            in2 => \N__28877\,
            in3 => \N__28844\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28826\,
            in2 => \N__28793\,
            in3 => \N__28754\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \bfn_11_12_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28743\,
            in2 => \N__28712\,
            in3 => \N__28673\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28663\,
            in2 => \N__28634\,
            in3 => \N__28595\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28590\,
            in2 => \N__28556\,
            in3 => \N__28520\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29446\,
            in2 => \N__29422\,
            in3 => \N__29369\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29356\,
            in2 => \N__29336\,
            in3 => \N__29300\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29291\,
            in2 => \N__29258\,
            in3 => \N__29225\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29218\,
            in2 => \N__29186\,
            in3 => \N__29150\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30403\,
            in2 => \N__29147\,
            in3 => \N__29120\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \bfn_11_13_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30349\,
            in2 => \N__29506\,
            in3 => \N__29117\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29491\,
            in2 => \N__29107\,
            in3 => \N__29063\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32597\,
            in2 => \N__29507\,
            in3 => \N__29060\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29495\,
            in2 => \N__29704\,
            in3 => \N__29639\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29632\,
            in2 => \N__29508\,
            in3 => \N__29579\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29499\,
            in2 => \N__29575\,
            in3 => \N__29513\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__33041\,
            in1 => \_gnd_net_\,
            in2 => \N__29509\,
            in3 => \N__29453\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_14_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010001010101010"
        )
    port map (
            in0 => \N__34844\,
            in1 => \N__34768\,
            in2 => \N__39728\,
            in3 => \N__34856\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47910\,
            ce => \N__33561\,
            sr => \N__47344\
        );

    \phase_controller_inst1.stoper_hc.target_time_13_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__34963\,
            in1 => \N__40529\,
            in2 => \_gnd_net_\,
            in3 => \N__35143\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47910\,
            ce => \N__33561\,
            sr => \N__47344\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto31_c_0_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40510\,
            in2 => \_gnd_net_\,
            in3 => \N__33142\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto31_cZ0Z_0\,
            ltout => \phase_controller_inst1.stoper_hc.un1_startlto31_cZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_16_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100000001"
        )
    port map (
            in0 => \N__40511\,
            in1 => \N__35604\,
            in2 => \N__29450\,
            in3 => \N__34816\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47904\,
            ce => \N__33565\,
            sr => \N__47354\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31099\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47897\,
            ce => \N__31958\,
            sr => \N__47362\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31060\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47897\,
            ce => \N__31958\,
            sr => \N__47362\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31927\,
            lcout => \current_shift_inst.elapsed_time_ns_1_fast_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47897\,
            ce => \N__31958\,
            sr => \N__47362\
        );

    \phase_controller_inst1.stoper_hc.target_time_5_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__34988\,
            in1 => \_gnd_net_\,
            in2 => \N__40558\,
            in3 => \N__34517\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47891\,
            ce => \N__33556\,
            sr => \N__47372\
        );

    \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000110011"
        )
    port map (
            in0 => \N__35057\,
            in1 => \N__40547\,
            in2 => \_gnd_net_\,
            in3 => \N__34987\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ1Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47891\,
            ce => \N__33556\,
            sr => \N__47372\
        );

    \phase_controller_inst1.stoper_hc.target_time_19_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__40546\,
            in1 => \N__36800\,
            in2 => \_gnd_net_\,
            in3 => \N__35228\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47891\,
            ce => \N__33556\,
            sr => \N__47372\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29741\,
            lcout => \current_shift_inst.un4_control_input_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29729\,
            lcout => \current_shift_inst.un4_control_input_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31415\,
            lcout => \current_shift_inst.un4_control_input_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31067\,
            lcout => \current_shift_inst.un4_control_input_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31028\,
            lcout => \current_shift_inst.un4_control_input_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30998\,
            lcout => \current_shift_inst.un4_control_input_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30968\,
            lcout => \current_shift_inst.un4_control_input_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30932\,
            lcout => \current_shift_inst.un4_control_input_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30896\,
            lcout => \current_shift_inst.un4_control_input_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31451\,
            lcout => \current_shift_inst.un4_control_input_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31382\,
            lcout => \current_shift_inst.un4_control_input_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31601\,
            lcout => \current_shift_inst.un4_control_input_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31571\,
            lcout => \current_shift_inst.un4_control_input_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31529\,
            lcout => \current_shift_inst.un4_control_input_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31487\,
            lcout => \current_shift_inst.un4_control_input_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31886\,
            lcout => \current_shift_inst.un4_control_input_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31736\,
            lcout => \current_shift_inst.un4_control_input_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31814\,
            lcout => \current_shift_inst.un4_control_input_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31634\,
            lcout => \current_shift_inst.un4_control_input_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31775\,
            lcout => \current_shift_inst.un4_control_input_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32189\,
            lcout => \current_shift_inst.un4_control_input_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31664\,
            lcout => \current_shift_inst.un4_control_input_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32225\,
            lcout => \current_shift_inst.un4_control_input_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31850\,
            lcout => \current_shift_inst.un4_control_input_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31700\,
            lcout => \current_shift_inst.un4_control_input_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32153\,
            lcout => \current_shift_inst.un4_control_input_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_i_31_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29968\,
            lcout => \current_shift_inst.z_i_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31967\,
            lcout => \current_shift_inst.un4_control_input_axb_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32114\,
            lcout => \current_shift_inst.un4_control_input_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32021\,
            lcout => \current_shift_inst.un4_control_input_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_11_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32075\,
            lcout => \current_shift_inst.un4_control_input_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.S1_rise_LC_11_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30314\,
            in2 => \_gnd_net_\,
            in3 => \N__30301\,
            lcout => \current_shift_inst.S1_riseZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47854\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.S1_sync0_LC_11_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32317\,
            lcout => \current_shift_inst.S1_syncZ0Z0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47854\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.S1_sync_prev_LC_11_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__30302\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.S1_sync_prevZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47854\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.S1_sync1_LC_11_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30308\,
            lcout => \current_shift_inst.S1_syncZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47854\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.phase_valid_LC_11_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100011101010"
        )
    port map (
            in0 => \N__30184\,
            in1 => \N__30293\,
            in2 => \N__32292\,
            in3 => \N__30232\,
            lcout => \current_shift_inst.phase_validZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47851\,
            ce => 'H',
            sr => \N__47411\
        );

    \SB_DFF_inst_PH1_MIN_D2_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30137\,
            lcout => \il_min_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47962\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MIN_D1_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__30152\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_min_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47962\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MIN_D2_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30131\,
            lcout => \il_min_comp2_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47954\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_2_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__30124\,
            in1 => \N__32909\,
            in2 => \N__30086\,
            in3 => \N__30047\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47936\,
            ce => \N__32554\,
            sr => \N__47297\
        );

    \current_shift_inst.PI_CTRL.integrator_31_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011111111"
        )
    port map (
            in0 => \N__33003\,
            in1 => \N__32900\,
            in2 => \N__30008\,
            in3 => \N__32720\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47927\,
            ce => \N__32555\,
            sr => \N__47305\
        );

    \current_shift_inst.PI_CTRL.integrator_24_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011111111"
        )
    port map (
            in0 => \N__33004\,
            in1 => \N__32891\,
            in2 => \N__30419\,
            in3 => \N__32721\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47921\,
            ce => \N__32530\,
            sr => \N__47312\
        );

    \current_shift_inst.PI_CTRL.integrator_25_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110111010101"
        )
    port map (
            in0 => \N__32722\,
            in1 => \N__30365\,
            in2 => \N__32907\,
            in3 => \N__33005\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47921\,
            ce => \N__32530\,
            sr => \N__47312\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__39958\,
            in1 => \N__40232\,
            in2 => \N__40127\,
            in3 => \N__37220\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47914\,
            ce => 'H',
            sr => \N__47318\
        );

    \phase_controller_inst1.stoper_hc.un1_m5_i_1_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110000"
        )
    port map (
            in0 => \N__35039\,
            in1 => \N__33119\,
            in2 => \N__36419\,
            in3 => \N__33113\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un1_m5_iZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_m5_i_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101110101010"
        )
    port map (
            in0 => \N__35180\,
            in1 => \N__32333\,
            in2 => \N__30320\,
            in3 => \N__39724\,
            lcout => \phase_controller_inst1.stoper_hc.un1_N_4\,
            ltout => \phase_controller_inst1.stoper_hc.un1_N_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto30_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34893\,
            in2 => \N__30317\,
            in3 => \N__33130\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlt31_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_11_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__40519\,
            in1 => \N__34648\,
            in2 => \_gnd_net_\,
            in3 => \N__34948\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47909\,
            ce => \N__33540\,
            sr => \N__47324\
        );

    \phase_controller_inst1.stoper_hc.target_time_2_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__35448\,
            in1 => \N__35542\,
            in2 => \N__34607\,
            in3 => \N__40524\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47909\,
            ce => \N__33540\,
            sr => \N__47324\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__35541\,
            in1 => \N__34561\,
            in2 => \N__40552\,
            in3 => \N__35450\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47909\,
            ce => \N__33540\,
            sr => \N__47324\
        );

    \phase_controller_inst1.stoper_hc.target_time_3_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__35449\,
            in1 => \N__35543\,
            in2 => \N__35278\,
            in3 => \N__40525\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47909\,
            ce => \N__33540\,
            sr => \N__47324\
        );

    \phase_controller_inst1.stoper_hc.target_time_1_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111110"
        )
    port map (
            in0 => \N__35540\,
            in1 => \N__35311\,
            in2 => \N__40551\,
            in3 => \N__35447\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47909\,
            ce => \N__33540\,
            sr => \N__47324\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__34949\,
            in1 => \N__40520\,
            in2 => \_gnd_net_\,
            in3 => \N__39766\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47909\,
            ce => \N__33540\,
            sr => \N__47324\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011010000"
        )
    port map (
            in0 => \N__40062\,
            in1 => \N__40200\,
            in2 => \N__36926\,
            in3 => \N__39936\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47903\,
            ce => 'H',
            sr => \N__47336\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__40199\,
            in1 => \N__40065\,
            in2 => \N__39961\,
            in3 => \N__37166\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47903\,
            ce => 'H',
            sr => \N__47336\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__40061\,
            in1 => \N__39937\,
            in2 => \N__37136\,
            in3 => \N__40201\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47903\,
            ce => 'H',
            sr => \N__47336\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__40197\,
            in1 => \N__40063\,
            in2 => \N__39959\,
            in3 => \N__33440\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47903\,
            ce => 'H',
            sr => \N__47336\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__40198\,
            in1 => \N__40064\,
            in2 => \N__39960\,
            in3 => \N__36890\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47903\,
            ce => 'H',
            sr => \N__47336\
        );

    \phase_controller_inst1.state_3_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110111010"
        )
    port map (
            in0 => \N__33851\,
            in1 => \N__34410\,
            in2 => \N__34450\,
            in3 => \N__33749\,
            lcout => \phase_controller_inst1.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47896\,
            ce => 'H',
            sr => \N__47345\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34321\,
            in2 => \_gnd_net_\,
            in3 => \N__34285\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.stoper_state_RNI38A6_0_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37774\,
            in2 => \_gnd_net_\,
            in3 => \N__38047\,
            lcout => \phase_controller_slave.stoper_tr.time_passed11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__38048\,
            in1 => \N__37973\,
            in2 => \_gnd_net_\,
            in3 => \N__37780\,
            lcout => \phase_controller_slave.stoper_tr.time_passed_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto30_3_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100000011"
        )
    port map (
            in0 => \N__34904\,
            in1 => \N__33146\,
            in2 => \N__40509\,
            in3 => \N__34873\,
            lcout => \phase_controller_inst1.stoper_hc.un1_start\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDLO51_11_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__30885\,
            in1 => \N__30844\,
            in2 => \N__30809\,
            in3 => \N__30763\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIDLO51_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.start_timer_tr_RNO_0_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33950\,
            in2 => \_gnd_net_\,
            in3 => \N__33987\,
            lcout => \phase_controller_slave.start_timer_tr_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1C4K_24_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31283\,
            in2 => \_gnd_net_\,
            in3 => \N__31188\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI1C4K_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHCE81_26_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__31373\,
            in1 => \N__30698\,
            in2 => \N__31337\,
            in3 => \N__30654\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIHCE81_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPB581_22_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__30508\,
            in1 => \N__30602\,
            in2 => \N__30470\,
            in3 => \N__30561\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPB581_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR32K_22_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30507\,
            in2 => \_gnd_net_\,
            in3 => \N__30466\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIR32K_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7K6K_26_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31372\,
            in2 => \_gnd_net_\,
            in3 => \N__31332\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI7K6K_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5S981_24_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__31282\,
            in1 => \N__31230\,
            in2 => \N__31193\,
            in3 => \N__31145\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5S981_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31018\,
            in2 => \N__31100\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_3\,
            ltout => OPEN,
            carryin => \bfn_12_19_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            clk => \N__47876\,
            ce => \N__31957\,
            sr => \N__47377\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30988\,
            in2 => \N__31061\,
            in3 => \N__31022\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            clk => \N__47876\,
            ce => \N__31957\,
            sr => \N__47377\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31019\,
            in2 => \N__30958\,
            in3 => \N__30992\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            clk => \N__47876\,
            ce => \N__31957\,
            sr => \N__47377\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30989\,
            in2 => \N__30922\,
            in3 => \N__30962\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            clk => \N__47876\,
            ce => \N__31957\,
            sr => \N__47377\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31621\,
            in2 => \N__30959\,
            in3 => \N__30926\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            clk => \N__47876\,
            ce => \N__31957\,
            sr => \N__47377\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31591\,
            in2 => \N__30923\,
            in3 => \N__31625\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            clk => \N__47876\,
            ce => \N__31957\,
            sr => \N__47377\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31622\,
            in2 => \N__31562\,
            in3 => \N__31595\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            clk => \N__47876\,
            ce => \N__31957\,
            sr => \N__47377\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31592\,
            in2 => \N__31520\,
            in3 => \N__31565\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            clk => \N__47876\,
            ce => \N__31957\,
            sr => \N__47377\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31561\,
            in2 => \N__31477\,
            in3 => \N__31523\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_11\,
            ltout => OPEN,
            carryin => \bfn_12_20_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            clk => \N__47869\,
            ce => \N__31956\,
            sr => \N__47383\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31519\,
            in2 => \N__31441\,
            in3 => \N__31481\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            clk => \N__47869\,
            ce => \N__31956\,
            sr => \N__47383\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31402\,
            in2 => \N__31478\,
            in3 => \N__31445\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            clk => \N__47869\,
            ce => \N__31956\,
            sr => \N__47383\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31906\,
            in2 => \N__31442\,
            in3 => \N__31406\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            clk => \N__47869\,
            ce => \N__31956\,
            sr => \N__47383\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31403\,
            in2 => \N__31876\,
            in3 => \N__31376\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            clk => \N__47869\,
            ce => \N__31956\,
            sr => \N__47383\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31907\,
            in2 => \N__31840\,
            in3 => \N__31880\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            clk => \N__47869\,
            ce => \N__31956\,
            sr => \N__47383\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31804\,
            in2 => \N__31877\,
            in3 => \N__31844\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            clk => \N__47869\,
            ce => \N__31956\,
            sr => \N__47383\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31765\,
            in2 => \N__31841\,
            in3 => \N__31808\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            clk => \N__47869\,
            ce => \N__31956\,
            sr => \N__47383\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_12_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31805\,
            in2 => \N__31726\,
            in3 => \N__31769\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_19\,
            ltout => OPEN,
            carryin => \bfn_12_21_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            clk => \N__47863\,
            ce => \N__31955\,
            sr => \N__47391\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31766\,
            in2 => \N__31690\,
            in3 => \N__31730\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            clk => \N__47863\,
            ce => \N__31955\,
            sr => \N__47391\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31654\,
            in2 => \N__31727\,
            in3 => \N__31694\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            clk => \N__47863\,
            ce => \N__31955\,
            sr => \N__47391\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32245\,
            in2 => \N__31691\,
            in3 => \N__31658\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            clk => \N__47863\,
            ce => \N__31955\,
            sr => \N__47391\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31655\,
            in2 => \N__32215\,
            in3 => \N__31628\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            clk => \N__47863\,
            ce => \N__31955\,
            sr => \N__47391\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32246\,
            in2 => \N__32179\,
            in3 => \N__32219\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            clk => \N__47863\,
            ce => \N__31955\,
            sr => \N__47391\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_12_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32143\,
            in2 => \N__32216\,
            in3 => \N__32183\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            clk => \N__47863\,
            ce => \N__31955\,
            sr => \N__47391\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32104\,
            in2 => \N__32180\,
            in3 => \N__32147\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            clk => \N__47863\,
            ce => \N__31955\,
            sr => \N__47391\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32144\,
            in2 => \N__32047\,
            in3 => \N__32108\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_27\,
            ltout => OPEN,
            carryin => \bfn_12_22_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            clk => \N__47858\,
            ce => \N__31954\,
            sr => \N__47395\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_12_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32105\,
            in2 => \N__31993\,
            in3 => \N__32069\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            clk => \N__47858\,
            ce => \N__31954\,
            sr => \N__47395\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_12_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32066\,
            in2 => \N__32048\,
            in3 => \N__32015\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            clk => \N__47858\,
            ce => \N__31954\,
            sr => \N__47395\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_12_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32012\,
            in2 => \N__31994\,
            in3 => \N__31961\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\,
            clk => \N__47858\,
            ce => \N__31954\,
            sr => \N__47395\
        );

    \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_12_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31934\,
            lcout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_12_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__36102\,
            in1 => \N__36054\,
            in2 => \_gnd_net_\,
            in3 => \N__36279\,
            lcout => \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.S1_LC_12_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34457\,
            lcout => s1_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47850\,
            ce => 'H',
            sr => \N__47404\
        );

    \phase_controller_inst1.stoper_tr.target_time_16_LC_12_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__48338\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47849\,
            ce => \N__43111\,
            sr => \N__47407\
        );

    \current_shift_inst.S3_rise_LC_12_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32267\,
            in2 => \_gnd_net_\,
            in3 => \N__32254\,
            lcout => \current_shift_inst.S3_riseZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47848\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.S3_sync0_LC_12_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33895\,
            lcout => \current_shift_inst.S3_syncZ0Z0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47848\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.S3_sync_prev_LC_12_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32255\,
            lcout => \current_shift_inst.S3_sync_prevZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47848\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_12_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36017\,
            in2 => \_gnd_net_\,
            in3 => \N__36278\,
            lcout => \phase_controller_inst1.stoper_tr.time_passed11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.S3_sync1_LC_12_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32261\,
            lcout => \current_shift_inst.S3_syncZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47848\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.hc_state_0_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__36574\,
            in1 => \N__36552\,
            in2 => \_gnd_net_\,
            in3 => \N__36452\,
            lcout => \delay_measurement_inst.hc_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47965\,
            ce => \N__35897\,
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MAX_D2_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33095\,
            lcout => \il_max_comp2_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47957\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_9_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__34641\,
            in1 => \N__36403\,
            in2 => \N__35350\,
            in3 => \N__35046\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_16_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101110011"
        )
    port map (
            in0 => \N__40718\,
            in1 => \N__36698\,
            in2 => \N__34807\,
            in3 => \N__44228\,
            lcout => measured_delay_hc_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47948\,
            ce => 'H',
            sr => \N__47292\
        );

    \delay_measurement_inst.delay_hc_reg_17_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101110011"
        )
    port map (
            in0 => \N__40719\,
            in1 => \N__36699\,
            in2 => \N__34732\,
            in3 => \N__44285\,
            lcout => measured_delay_hc_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47948\,
            ce => 'H',
            sr => \N__47292\
        );

    \delay_measurement_inst.delay_hc_reg_13_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__35131\,
            in1 => \N__40720\,
            in2 => \N__41396\,
            in3 => \N__40853\,
            lcout => measured_delay_hc_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47948\,
            ce => 'H',
            sr => \N__47292\
        );

    \delay_measurement_inst.delay_hc_reg_15_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__40717\,
            in1 => \N__35176\,
            in2 => \N__42016\,
            in3 => \N__36700\,
            lcout => measured_delay_hc_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47948\,
            ce => 'H',
            sr => \N__47292\
        );

    \current_shift_inst.PI_CTRL.integrator_27_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011111111"
        )
    port map (
            in0 => \N__33006\,
            in1 => \N__32908\,
            in2 => \N__32738\,
            in3 => \N__32723\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47938\,
            ce => \N__32561\,
            sr => \N__47298\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto13_3_1_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__34673\,
            in1 => \N__34636\,
            in2 => \N__35368\,
            in3 => \N__35136\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto13_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_11_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__34640\,
            in1 => \N__40722\,
            in2 => \N__41495\,
            in3 => \N__40844\,
            lcout => measured_delay_hc_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47929\,
            ce => 'H',
            sr => \N__47306\
        );

    \delay_measurement_inst.delay_hc_reg_6_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111100010"
        )
    port map (
            in0 => \N__35045\,
            in1 => \N__40723\,
            in2 => \N__44021\,
            in3 => \N__40845\,
            lcout => measured_delay_hc_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47929\,
            ce => 'H',
            sr => \N__47306\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_12_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__33155\,
            in1 => \N__34208\,
            in2 => \N__39723\,
            in3 => \N__34220\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto30_2_0_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__36823\,
            in1 => \N__36724\,
            in2 => \N__36767\,
            in3 => \N__35213\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto30_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto8_0_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__35489\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34556\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto8Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_m2_e_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__39591\,
            in1 => \N__34201\,
            in2 => \N__35274\,
            in3 => \N__34219\,
            lcout => \phase_controller_inst1.stoper_hc.un1_m2_eZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_11_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__34202\,
            in1 => \N__34193\,
            in2 => \_gnd_net_\,
            in3 => \N__35267\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__36792\,
            in1 => \N__33107\,
            in2 => \N__33101\,
            in3 => \N__35214\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlt31\,
            ltout => \phase_controller_inst1.stoper_hc.un2_startlt31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto31_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33098\,
            in3 => \N__40461\,
            lcout => \phase_controller_inst1.stoper_hc.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__39938\,
            in1 => \N__40006\,
            in2 => \_gnd_net_\,
            in3 => \N__40202\,
            lcout => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.start_timer_hc_RNO_0_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42785\,
            in2 => \_gnd_net_\,
            in3 => \N__42989\,
            lcout => \phase_controller_slave.start_timer_hc_RNO_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33293\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_13_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33266\,
            in2 => \N__33275\,
            in3 => \N__37026\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33251\,
            in2 => \N__33260\,
            in3 => \N__37009\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33236\,
            in2 => \N__33245\,
            in3 => \N__36964\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33230\,
            in2 => \N__33224\,
            in3 => \N__36937\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33200\,
            in2 => \N__33215\,
            in3 => \N__36901\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33179\,
            in2 => \N__33194\,
            in3 => \N__36874\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33161\,
            in2 => \N__33173\,
            in3 => \N__37231\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33422\,
            in2 => \N__33434\,
            in3 => \N__37204\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \bfn_13_14_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33392\,
            in2 => \N__33416\,
            in3 => \N__37177\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33368\,
            in2 => \N__33386\,
            in3 => \N__40301\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33350\,
            in2 => \N__33362\,
            in3 => \N__37147\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33344\,
            in2 => \N__33599\,
            in3 => \N__37120\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__40280\,
            in1 => \N__33323\,
            in2 => \N__33338\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33305\,
            in2 => \N__33317\,
            in3 => \N__37096\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33299\,
            in2 => \N__33614\,
            in3 => \N__40259\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33482\,
            in2 => \N__33494\,
            in3 => \N__37373\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \bfn_13_15_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33476\,
            in2 => \N__33587\,
            in3 => \N__37346\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37321\,
            in1 => \N__33470\,
            in2 => \N__33578\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33449\,
            in2 => \N__33464\,
            in3 => \N__39836\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33443\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__40060\,
            in1 => \N__39923\,
            in2 => \_gnd_net_\,
            in3 => \N__40193\,
            lcout => \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34322\,
            in1 => \N__37030\,
            in2 => \_gnd_net_\,
            in3 => \N__34286\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_8_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__35414\,
            in1 => \N__35597\,
            in2 => \N__40536\,
            in3 => \N__35499\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47898\,
            ce => \N__33557\,
            sr => \N__47346\
        );

    \phase_controller_inst1.stoper_hc.target_time_15_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__35594\,
            in1 => \N__40488\,
            in2 => \N__35194\,
            in3 => \N__35412\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47898\,
            ce => \N__33557\,
            sr => \N__47346\
        );

    \phase_controller_inst1.stoper_hc.target_time_12_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__35369\,
            in1 => \N__40487\,
            in2 => \_gnd_net_\,
            in3 => \N__34992\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47898\,
            ce => \N__33557\,
            sr => \N__47346\
        );

    \phase_controller_inst1.stoper_hc.target_time_17_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000000010001"
        )
    port map (
            in0 => \N__40489\,
            in1 => \N__35595\,
            in2 => \N__34742\,
            in3 => \N__34775\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47898\,
            ce => \N__33557\,
            sr => \N__47346\
        );

    \phase_controller_inst1.stoper_hc.target_time_18_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001100000010"
        )
    port map (
            in0 => \N__35413\,
            in1 => \N__35596\,
            in2 => \N__40535\,
            in3 => \N__35096\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47898\,
            ce => \N__33557\,
            sr => \N__47346\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_0_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__39915\,
            in1 => \N__40184\,
            in2 => \N__40100\,
            in3 => \N__34294\,
            lcout => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47892\,
            ce => \N__35887\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_1_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001010000"
        )
    port map (
            in0 => \N__34295\,
            in1 => \N__40066\,
            in2 => \N__40229\,
            in3 => \N__39916\,
            lcout => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47892\,
            ce => \N__35887\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_0_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__36065\,
            in1 => \N__36245\,
            in2 => \N__36204\,
            in3 => \N__39219\,
            lcout => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47892\,
            ce => \N__35887\,
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.stoper_state_0_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__43519\,
            in1 => \N__43032\,
            in2 => \N__43733\,
            in3 => \N__43790\,
            lcout => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47892\,
            ce => \N__35887\,
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.stoper_state_1_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001010000"
        )
    port map (
            in0 => \N__43033\,
            in1 => \N__43728\,
            in2 => \N__43833\,
            in3 => \N__43520\,
            lcout => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47892\,
            ce => \N__35887\,
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.stoper_state_0_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__37792\,
            in1 => \N__37974\,
            in2 => \N__38104\,
            in3 => \N__38698\,
            lcout => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47892\,
            ce => \N__35887\,
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.stoper_state_1_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000001000100"
        )
    port map (
            in0 => \N__38699\,
            in1 => \N__38062\,
            in2 => \N__38008\,
            in3 => \N__37793\,
            lcout => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47892\,
            ce => \N__35887\,
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_16_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__37791\,
            in1 => \N__38058\,
            in2 => \N__37972\,
            in3 => \N__35630\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47885\,
            ce => 'H',
            sr => \N__47363\
        );

    \phase_controller_slave.stoper_tr.time_passed_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__33778\,
            in1 => \N__38189\,
            in2 => \N__33794\,
            in3 => \N__38697\,
            lcout => \phase_controller_slave.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47885\,
            ce => 'H',
            sr => \N__47363\
        );

    \phase_controller_slave.state_0_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111000001010"
        )
    port map (
            in0 => \N__33761\,
            in1 => \N__33994\,
            in2 => \N__33779\,
            in3 => \N__33945\,
            lcout => \phase_controller_slave.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47885\,
            ce => 'H',
            sr => \N__47363\
        );

    \phase_controller_slave.state_RNIVDE2_0_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33774\,
            in2 => \_gnd_net_\,
            in3 => \N__33760\,
            lcout => \phase_controller_slave.state_RNIVDE2Z0Z_0\,
            ltout => \phase_controller_slave.state_RNIVDE2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.state_3_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__42813\,
            in1 => \N__42861\,
            in2 => \N__33752\,
            in3 => \N__33742\,
            lcout => \phase_controller_slave.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47885\,
            ce => 'H',
            sr => \N__47363\
        );

    \phase_controller_slave.state_ns_i_a2_1_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33718\,
            in2 => \_gnd_net_\,
            in3 => \N__42891\,
            lcout => state_ns_i_a2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_4_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__33729\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42892\,
            lcout => phase_controller_inst1_state_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47882\,
            ce => 'H',
            sr => \N__47373\
        );

    \phase_controller_slave.S2_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101100001000"
        )
    port map (
            in0 => \N__33625\,
            in1 => \N__42812\,
            in2 => \N__33872\,
            in3 => \N__33941\,
            lcout => s4_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47882\,
            ce => 'H',
            sr => \N__47373\
        );

    \phase_controller_slave.state_1_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__33995\,
            in1 => \N__42781\,
            in2 => \N__33949\,
            in3 => \N__42988\,
            lcout => \phase_controller_slave.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47882\,
            ce => 'H',
            sr => \N__47373\
        );

    \phase_controller_slave.start_timer_tr_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__42893\,
            in1 => \N__37921\,
            in2 => \N__33920\,
            in3 => \N__33908\,
            lcout => \phase_controller_slave.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47882\,
            ce => 'H',
            sr => \N__47373\
        );

    \phase_controller_slave.S1_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010100000"
        )
    port map (
            in0 => \N__42817\,
            in1 => \_gnd_net_\,
            in2 => \N__33871\,
            in3 => \N__33883\,
            lcout => s3_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47878\,
            ce => 'H',
            sr => \N__47378\
        );

    \phase_controller_inst1.T23_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__34142\,
            in1 => \N__33864\,
            in2 => \_gnd_net_\,
            in3 => \N__34453\,
            lcout => shift_flag_start,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47878\,
            ce => 'H',
            sr => \N__47378\
        );

    \phase_controller_inst1.start_timer_tr_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__33844\,
            in1 => \N__33824\,
            in2 => \N__36176\,
            in3 => \N__42904\,
            lcout => \phase_controller_inst1.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47865\,
            ce => 'H',
            sr => \N__47392\
        );

    \phase_controller_inst1.state_RNI7NN7_0_LC_13_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33813\,
            in2 => \_gnd_net_\,
            in3 => \N__33802\,
            lcout => \phase_controller_inst1.state_RNI7NN7Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.time_passed_LC_13_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__33817\,
            in1 => \N__34252\,
            in2 => \N__33833\,
            in3 => \N__39220\,
            lcout => \phase_controller_inst1.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47860\,
            ce => 'H',
            sr => \N__47396\
        );

    \phase_controller_inst1.start_timer_tr_RNO_0_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34136\,
            in2 => \_gnd_net_\,
            in3 => \N__34177\,
            lcout => \phase_controller_inst1.start_timer_tr_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_0_LC_13_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111000001010"
        )
    port map (
            in0 => \N__33803\,
            in1 => \N__34178\,
            in2 => \N__33818\,
            in3 => \N__34140\,
            lcout => \phase_controller_inst1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47860\,
            ce => 'H',
            sr => \N__47396\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_13_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__36060\,
            in1 => \N__36255\,
            in2 => \N__36180\,
            in3 => \N__34037\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47860\,
            ce => 'H',
            sr => \N__47396\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34091\,
            in2 => \N__38620\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_24_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38591\,
            in2 => \_gnd_net_\,
            in3 => \N__34019\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_13_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34082\,
            in2 => \N__38570\,
            in3 => \N__34016\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_13_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38909\,
            in2 => \_gnd_net_\,
            in3 => \N__34013\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_13_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38891\,
            in2 => \_gnd_net_\,
            in3 => \N__34010\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_13_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38873\,
            in2 => \_gnd_net_\,
            in3 => \N__34007\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_13_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38852\,
            in2 => \_gnd_net_\,
            in3 => \N__34004\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_13_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38834\,
            in2 => \_gnd_net_\,
            in3 => \N__34001\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_13_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38816\,
            in3 => \N__33998\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9\,
            ltout => OPEN,
            carryin => \bfn_13_25_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_13_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38789\,
            in2 => \_gnd_net_\,
            in3 => \N__34055\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_13_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39074\,
            in2 => \_gnd_net_\,
            in3 => \N__34052\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_13_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39056\,
            in2 => \_gnd_net_\,
            in3 => \N__34049\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_13_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39038\,
            in2 => \_gnd_net_\,
            in3 => \N__34046\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_13_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39020\,
            in2 => \_gnd_net_\,
            in3 => \N__34043\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_13_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39002\,
            in2 => \_gnd_net_\,
            in3 => \N__34040\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_13_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38968\,
            in2 => \_gnd_net_\,
            in3 => \N__34028\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_13_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38945\,
            in2 => \_gnd_net_\,
            in3 => \N__34025\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17\,
            ltout => OPEN,
            carryin => \bfn_13_26_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_13_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38927\,
            in2 => \_gnd_net_\,
            in3 => \N__34022\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_13_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39242\,
            in2 => \_gnd_net_\,
            in3 => \N__34094\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_13_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34238\,
            in2 => \_gnd_net_\,
            in3 => \N__39205\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_13_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__39206\,
            in1 => \_gnd_net_\,
            in2 => \N__34248\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.S2_LC_13_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34141\,
            lcout => s2_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47847\,
            ce => 'H',
            sr => \N__47421\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_14_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__39104\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39127\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_335_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.prev_hc_sig_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__36451\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.prev_hc_sigZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47982\,
            ce => 'H',
            sr => \N__47273\
        );

    \delay_measurement_inst.stop_timer_hc_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__36573\,
            in1 => \N__36553\,
            in2 => \N__47464\,
            in3 => \N__36441\,
            lcout => \delay_measurement_inst.stop_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47974\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_5_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__41205\,
            in1 => \N__34511\,
            in2 => \N__40729\,
            in3 => \N__40852\,
            lcout => measured_delay_hc_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47958\,
            ce => 'H',
            sr => \N__47289\
        );

    \delay_measurement_inst.delay_hc_reg_12_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__40709\,
            in1 => \N__41447\,
            in2 => \N__35360\,
            in3 => \N__40850\,
            lcout => measured_delay_hc_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47958\,
            ce => 'H',
            sr => \N__47289\
        );

    \delay_measurement_inst.delay_hc_reg_3_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000011001010"
        )
    port map (
            in0 => \N__35252\,
            in1 => \N__42436\,
            in2 => \N__40728\,
            in3 => \N__40851\,
            lcout => measured_delay_hc_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47958\,
            ce => 'H',
            sr => \N__47289\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41550\,
            in1 => \N__41442\,
            in2 => \N__41395\,
            in3 => \N__41488\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_11_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41487\,
            in1 => \N__44284\,
            in2 => \N__41446\,
            in3 => \N__44305\,
            lcout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITRKR_5_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41207\,
            in2 => \_gnd_net_\,
            in3 => \N__42475\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQI9C2_13_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__41391\,
            in1 => \N__34187\,
            in2 => \N__34181\,
            in3 => \N__44227\,
            lcout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_18_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111011000"
        )
    port map (
            in0 => \N__40666\,
            in1 => \N__44309\,
            in2 => \N__35095\,
            in3 => \N__40846\,
            lcout => measured_delay_hc_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47949\,
            ce => 'H',
            sr => \N__47293\
        );

    \delay_measurement_inst.delay_hc_reg_2_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__40847\,
            in1 => \N__44357\,
            in2 => \N__34606\,
            in3 => \N__40670\,
            lcout => measured_delay_hc_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47949\,
            ce => 'H',
            sr => \N__47293\
        );

    \delay_measurement_inst.delay_hc_reg_7_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__40848\,
            in1 => \N__34543\,
            in2 => \N__41711\,
            in3 => \N__40671\,
            lcout => measured_delay_hc_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47949\,
            ce => 'H',
            sr => \N__47293\
        );

    \delay_measurement_inst.delay_hc_reg_8_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001010"
        )
    port map (
            in0 => \N__35488\,
            in1 => \N__41644\,
            in2 => \N__40716\,
            in3 => \N__40849\,
            lcout => measured_delay_hc_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47949\,
            ce => 'H',
            sr => \N__47293\
        );

    \phase_controller_inst1.state_1_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__34176\,
            in1 => \N__34379\,
            in2 => \N__34123\,
            in3 => \N__34346\,
            lcout => \phase_controller_inst1.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47939\,
            ce => 'H',
            sr => \N__47299\
        );

    \delay_measurement_inst.delay_hc_reg_10_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__40653\,
            in1 => \N__34680\,
            in2 => \N__41555\,
            in3 => \N__40842\,
            lcout => measured_delay_hc_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47939\,
            ce => 'H',
            sr => \N__47299\
        );

    \delay_measurement_inst.delay_hc_reg_23_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__40652\,
            in1 => \N__34486\,
            in2 => \_gnd_net_\,
            in3 => \N__40843\,
            lcout => measured_delay_hc_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47939\,
            ce => 'H',
            sr => \N__47299\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__37064\,
            in1 => \N__39659\,
            in2 => \N__39641\,
            in3 => \N__34472\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34259\,
            in1 => \N__38624\,
            in2 => \_gnd_net_\,
            in3 => \N__39221\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_m2_e_1_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34512\,
            in2 => \_gnd_net_\,
            in3 => \N__39759\,
            lcout => \phase_controller_inst1.stoper_hc.un1_m2_eZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35090\,
            in1 => \N__34736\,
            in2 => \N__36746\,
            in3 => \N__34809\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__34557\,
            in1 => \N__34672\,
            in2 => \N__35500\,
            in3 => \N__35089\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_m2_e_2_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34595\,
            in2 => \_gnd_net_\,
            in3 => \N__35304\,
            lcout => \phase_controller_inst1.stoper_hc.un1_m2_eZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_8_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__34808\,
            in1 => \N__35187\,
            in2 => \N__34741\,
            in3 => \N__35132\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_3_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39677\,
            in2 => \_gnd_net_\,
            in3 => \N__34487\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_RNO_1_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34451\,
            in2 => \_gnd_net_\,
            in3 => \N__34411\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.start_timer_hc_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011110010"
        )
    port map (
            in0 => \N__40024\,
            in1 => \N__34463\,
            in2 => \N__34466\,
            in3 => \N__42908\,
            lcout => \phase_controller_inst1.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47922\,
            ce => 'H',
            sr => \N__47313\
        );

    \phase_controller_inst1.start_timer_hc_RNO_0_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34371\,
            in2 => \_gnd_net_\,
            in3 => \N__34340\,
            lcout => \phase_controller_inst1.start_timer_hc_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_2_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101000110000"
        )
    port map (
            in0 => \N__34452\,
            in1 => \N__34345\,
            in2 => \N__34378\,
            in3 => \N__34412\,
            lcout => \phase_controller_inst1.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47922\,
            ce => 'H',
            sr => \N__47313\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__39957\,
            in1 => \N__40025\,
            in2 => \N__37358\,
            in3 => \N__40231\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47922\,
            ce => 'H',
            sr => \N__47313\
        );

    \phase_controller_inst1.stoper_hc.time_passed_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__34341\,
            in1 => \N__34314\,
            in2 => \N__34358\,
            in3 => \N__34293\,
            lcout => \phase_controller_inst1.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47922\,
            ce => 'H',
            sr => \N__47313\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39956\,
            in2 => \_gnd_net_\,
            in3 => \N__40230\,
            lcout => \phase_controller_inst1.stoper_hc.time_passed11\,
            ltout => \phase_controller_inst1.stoper_hc.time_passed11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34298\,
            in3 => \N__34292\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__39950\,
            in1 => \N__40239\,
            in2 => \N__40125\,
            in3 => \N__37331\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47915\,
            ce => 'H',
            sr => \N__47319\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__40233\,
            in1 => \N__40113\,
            in2 => \N__37310\,
            in3 => \N__39952\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47915\,
            ce => 'H',
            sr => \N__47319\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__39949\,
            in1 => \N__40238\,
            in2 => \N__40124\,
            in3 => \N__37085\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47915\,
            ce => 'H',
            sr => \N__47319\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__40234\,
            in1 => \N__40114\,
            in2 => \N__36998\,
            in3 => \N__39953\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47915\,
            ce => 'H',
            sr => \N__47319\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__39951\,
            in1 => \N__40240\,
            in2 => \N__40126\,
            in3 => \N__36953\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47915\,
            ce => 'H',
            sr => \N__47319\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__40236\,
            in1 => \N__40116\,
            in2 => \N__37193\,
            in3 => \N__39955\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47915\,
            ce => 'H',
            sr => \N__47319\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__39948\,
            in1 => \N__40237\,
            in2 => \N__40123\,
            in3 => \N__37109\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47915\,
            ce => 'H',
            sr => \N__47319\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__40235\,
            in1 => \N__40115\,
            in2 => \N__36863\,
            in3 => \N__39954\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47915\,
            ce => 'H',
            sr => \N__47319\
        );

    \phase_controller_slave.stoper_hc.target_time_0_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__34986\,
            in1 => \N__40463\,
            in2 => \N__35615\,
            in3 => \N__39592\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47911\,
            ce => \N__39801\,
            sr => \N__47325\
        );

    \phase_controller_slave.stoper_hc.target_time_9_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001000000011"
        )
    port map (
            in0 => \N__36417\,
            in1 => \N__35600\,
            in2 => \N__40531\,
            in3 => \N__34985\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47911\,
            ce => \N__39801\,
            sr => \N__47325\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto31_d_0_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__40462\,
            in1 => \N__34903\,
            in2 => \_gnd_net_\,
            in3 => \N__34877\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto31_dZ0Z_0\,
            ltout => \phase_controller_inst1.stoper_hc.un1_startlto31_dZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.target_time_14_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000110011001100"
        )
    port map (
            in0 => \N__39722\,
            in1 => \N__34843\,
            in2 => \N__34823\,
            in3 => \N__34771\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47911\,
            ce => \N__39801\,
            sr => \N__47325\
        );

    \phase_controller_slave.stoper_hc.target_time_16_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000000010001"
        )
    port map (
            in0 => \N__35598\,
            in1 => \N__40464\,
            in2 => \N__34820\,
            in3 => \N__34769\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47911\,
            ce => \N__39801\,
            sr => \N__47325\
        );

    \phase_controller_slave.stoper_hc.target_time_17_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001100000001"
        )
    port map (
            in0 => \N__34770\,
            in1 => \N__35599\,
            in2 => \N__40530\,
            in3 => \N__34737\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47911\,
            ce => \N__39801\,
            sr => \N__47325\
        );

    \phase_controller_slave.stoper_hc.target_time_10_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__40475\,
            in1 => \N__34681\,
            in2 => \_gnd_net_\,
            in3 => \N__35009\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47905\,
            ce => \N__39817\,
            sr => \N__47337\
        );

    \phase_controller_slave.stoper_hc.target_time_11_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__35010\,
            in1 => \N__40476\,
            in2 => \_gnd_net_\,
            in3 => \N__34649\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47905\,
            ce => \N__39817\,
            sr => \N__47337\
        );

    \phase_controller_slave.stoper_hc.target_time_2_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__35584\,
            in1 => \N__34596\,
            in2 => \N__40534\,
            in3 => \N__35437\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47905\,
            ce => \N__39817\,
            sr => \N__47337\
        );

    \phase_controller_slave.stoper_hc.target_time_7_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__35439\,
            in1 => \N__35586\,
            in2 => \N__34565\,
            in3 => \N__40486\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47905\,
            ce => \N__39817\,
            sr => \N__47337\
        );

    \phase_controller_slave.stoper_hc.target_time_5_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__40478\,
            in1 => \N__35012\,
            in2 => \_gnd_net_\,
            in3 => \N__34513\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47905\,
            ce => \N__39817\,
            sr => \N__47337\
        );

    \phase_controller_slave.stoper_hc.target_time_12_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__35011\,
            in1 => \N__40477\,
            in2 => \_gnd_net_\,
            in3 => \N__35364\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47905\,
            ce => \N__39817\,
            sr => \N__47337\
        );

    \phase_controller_slave.stoper_hc.target_time_1_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111110"
        )
    port map (
            in0 => \N__35583\,
            in1 => \N__35315\,
            in2 => \N__40533\,
            in3 => \N__35436\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47905\,
            ce => \N__39817\,
            sr => \N__47337\
        );

    \phase_controller_slave.stoper_hc.target_time_3_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__35438\,
            in1 => \N__35585\,
            in2 => \N__35279\,
            in3 => \N__40485\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47905\,
            ce => \N__39817\,
            sr => \N__47337\
        );

    \phase_controller_slave.stoper_hc.target_time_19_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100110011"
        )
    port map (
            in0 => \N__35221\,
            in1 => \N__40471\,
            in2 => \_gnd_net_\,
            in3 => \N__36799\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47899\,
            ce => \N__39818\,
            sr => \N__47347\
        );

    \phase_controller_slave.stoper_hc.target_time_15_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__35451\,
            in1 => \N__35611\,
            in2 => \N__40537\,
            in3 => \N__35195\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47899\,
            ce => \N__39818\,
            sr => \N__47347\
        );

    \phase_controller_slave.stoper_hc.target_time_13_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__35014\,
            in1 => \N__40497\,
            in2 => \_gnd_net_\,
            in3 => \N__35144\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47899\,
            ce => \N__39818\,
            sr => \N__47347\
        );

    \phase_controller_slave.stoper_hc.target_time_4_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__40498\,
            in1 => \N__35015\,
            in2 => \_gnd_net_\,
            in3 => \N__39767\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47899\,
            ce => \N__39818\,
            sr => \N__47347\
        );

    \phase_controller_slave.stoper_hc.target_time_18_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001100000010"
        )
    port map (
            in0 => \N__35091\,
            in1 => \N__40502\,
            in2 => \N__35618\,
            in3 => \N__35452\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47899\,
            ce => \N__39818\,
            sr => \N__47347\
        );

    \phase_controller_slave.stoper_hc.target_timeZ0Z_6_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__40496\,
            in1 => \N__35056\,
            in2 => \_gnd_net_\,
            in3 => \N__35013\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ1Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47899\,
            ce => \N__39818\,
            sr => \N__47347\
        );

    \phase_controller_slave.stoper_hc.target_time_8_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__35610\,
            in1 => \N__35501\,
            in2 => \N__40532\,
            in3 => \N__35453\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47899\,
            ce => \N__39818\,
            sr => \N__47347\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37649\,
            in2 => \N__37733\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_18_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38381\,
            in2 => \_gnd_net_\,
            in3 => \N__35390\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37685\,
            in2 => \N__38360\,
            in3 => \N__35387\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38336\,
            in2 => \_gnd_net_\,
            in3 => \N__35384\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38315\,
            in2 => \_gnd_net_\,
            in3 => \N__35381\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38294\,
            in3 => \N__35378\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38269\,
            in2 => \_gnd_net_\,
            in3 => \N__35375\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38239\,
            in2 => \_gnd_net_\,
            in3 => \N__35372\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38218\,
            in2 => \_gnd_net_\,
            in3 => \N__35651\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9\,
            ltout => OPEN,
            carryin => \bfn_14_19_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38548\,
            in2 => \_gnd_net_\,
            in3 => \N__35648\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38527\,
            in2 => \_gnd_net_\,
            in3 => \N__35645\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38506\,
            in2 => \_gnd_net_\,
            in3 => \N__35642\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38485\,
            in2 => \_gnd_net_\,
            in3 => \N__35639\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38464\,
            in2 => \_gnd_net_\,
            in3 => \N__35636\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38443\,
            in2 => \_gnd_net_\,
            in3 => \N__35633\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38407\,
            in3 => \N__35624\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38767\,
            in2 => \_gnd_net_\,
            in3 => \N__35621\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17\,
            ltout => OPEN,
            carryin => \bfn_14_20_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38743\,
            in2 => \_gnd_net_\,
            in3 => \N__35711\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38722\,
            in2 => \_gnd_net_\,
            in3 => \N__35708\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_17_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__37842\,
            in1 => \N__38117\,
            in2 => \N__38012\,
            in3 => \N__35705\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47879\,
            ce => 'H',
            sr => \N__47379\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_18_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__38113\,
            in1 => \N__37991\,
            in2 => \N__37869\,
            in3 => \N__35699\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47879\,
            ce => 'H',
            sr => \N__47379\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_19_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__37843\,
            in1 => \N__38118\,
            in2 => \N__38013\,
            in3 => \N__35693\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47879\,
            ce => 'H',
            sr => \N__47379\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_2_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__38114\,
            in1 => \N__37992\,
            in2 => \N__37870\,
            in3 => \N__35687\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47879\,
            ce => 'H',
            sr => \N__47379\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_3_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010000100"
        )
    port map (
            in0 => \N__37844\,
            in1 => \N__35678\,
            in2 => \N__38014\,
            in3 => \N__38120\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47879\,
            ce => 'H',
            sr => \N__47379\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_4_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__38115\,
            in1 => \N__37993\,
            in2 => \N__37871\,
            in3 => \N__35669\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47879\,
            ce => 'H',
            sr => \N__47379\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_5_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__37845\,
            in1 => \N__38119\,
            in2 => \N__38015\,
            in3 => \N__35660\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47879\,
            ce => 'H',
            sr => \N__47379\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_6_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__38116\,
            in1 => \N__37994\,
            in2 => \N__37872\,
            in3 => \N__35759\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47879\,
            ce => 'H',
            sr => \N__47379\
        );

    \phase_controller_slave.stoper_tr.target_time_16_LC_14_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48334\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47871\,
            ce => \N__43354\,
            sr => \N__47384\
        );

    \phase_controller_slave.stoper_tr.target_time_8_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43445\,
            in2 => \_gnd_net_\,
            in3 => \N__46823\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47871\,
            ce => \N__43354\,
            sr => \N__47384\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__36316\,
            in1 => \N__36104\,
            in2 => \N__36055\,
            in3 => \N__35750\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47866\,
            ce => 'H',
            sr => \N__47393\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_14_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__36317\,
            in1 => \N__36105\,
            in2 => \N__36056\,
            in3 => \N__35744\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47866\,
            ce => 'H',
            sr => \N__47393\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_14_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__36103\,
            in1 => \N__36021\,
            in2 => \_gnd_net_\,
            in3 => \N__36315\,
            lcout => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_1_LC_14_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__43585\,
            in1 => \N__43853\,
            in2 => \N__43732\,
            in3 => \N__37679\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47866\,
            ce => 'H',
            sr => \N__47393\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_14_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__36294\,
            in1 => \N__36155\,
            in2 => \N__36064\,
            in3 => \N__35735\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47861\,
            ce => 'H',
            sr => \N__47397\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_14_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__36034\,
            in1 => \N__36287\,
            in2 => \N__36181\,
            in3 => \N__35729\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47861\,
            ce => 'H',
            sr => \N__47397\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_14_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__36289\,
            in1 => \N__36144\,
            in2 => \N__36062\,
            in3 => \N__35723\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47861\,
            ce => 'H',
            sr => \N__47397\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_14_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__36035\,
            in1 => \N__36290\,
            in2 => \N__36182\,
            in3 => \N__35813\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47861\,
            ce => 'H',
            sr => \N__47397\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_14_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__36291\,
            in1 => \N__36148\,
            in2 => \N__36063\,
            in3 => \N__35807\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47861\,
            ce => 'H',
            sr => \N__47397\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_14_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__36036\,
            in1 => \N__36292\,
            in2 => \N__36183\,
            in3 => \N__35801\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47861\,
            ce => 'H',
            sr => \N__47397\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_14_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__36288\,
            in1 => \N__36143\,
            in2 => \N__36061\,
            in3 => \N__35795\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47861\,
            ce => 'H',
            sr => \N__47397\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_14_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__36037\,
            in1 => \N__36293\,
            in2 => \N__36184\,
            in3 => \N__35789\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47861\,
            ce => 'H',
            sr => \N__47397\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_14_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010000100"
        )
    port map (
            in0 => \N__36000\,
            in1 => \N__35783\,
            in2 => \N__36205\,
            in3 => \N__36318\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47855\,
            ce => 'H',
            sr => \N__47400\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_14_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__36322\,
            in1 => \N__36193\,
            in2 => \N__36052\,
            in3 => \N__35777\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47855\,
            ce => 'H',
            sr => \N__47400\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_14_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__36003\,
            in1 => \N__36325\,
            in2 => \N__36208\,
            in3 => \N__35771\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47855\,
            ce => 'H',
            sr => \N__47400\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_14_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__36324\,
            in1 => \N__36197\,
            in2 => \N__36053\,
            in3 => \N__35765\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47855\,
            ce => 'H',
            sr => \N__47400\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_14_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__36002\,
            in1 => \N__36323\,
            in2 => \N__36207\,
            in3 => \N__36350\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47855\,
            ce => 'H',
            sr => \N__47400\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_14_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__36321\,
            in1 => \N__36192\,
            in2 => \N__36051\,
            in3 => \N__36344\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47855\,
            ce => 'H',
            sr => \N__47400\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_14_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__36001\,
            in1 => \N__36319\,
            in2 => \N__36206\,
            in3 => \N__36338\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47855\,
            ce => 'H',
            sr => \N__47400\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_14_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__36320\,
            in1 => \N__36191\,
            in2 => \N__36050\,
            in3 => \N__36332\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47855\,
            ce => 'H',
            sr => \N__47400\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_1_LC_14_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000001100010"
        )
    port map (
            in0 => \N__36326\,
            in1 => \N__36016\,
            in2 => \N__36209\,
            in3 => \N__39201\,
            lcout => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47852\,
            ce => \N__35861\,
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_DELAY_TR1_LC_15_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35912\,
            lcout => delay_tr_d1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47993\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_DELAY_TR2_LC_15_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35903\,
            lcout => delay_tr_d2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47993\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.tr_state_0_LC_15_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001100110"
        )
    port map (
            in0 => \N__36525\,
            in1 => \N__36507\,
            in2 => \_gnd_net_\,
            in3 => \N__36491\,
            lcout => \delay_measurement_inst.tr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47990\,
            ce => \N__35879\,
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.prev_tr_sig_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36535\,
            lcout => \delay_measurement_inst.prev_tr_sigZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47983\,
            ce => 'H',
            sr => \N__47274\
        );

    \delay_measurement_inst.start_timer_hc_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__36575\,
            in1 => \N__36557\,
            in2 => \_gnd_net_\,
            in3 => \N__36440\,
            lcout => \delay_measurement_inst.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47983\,
            ce => 'H',
            sr => \N__47274\
        );

    \delay_measurement_inst.delay_hc_timer.running_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__39140\,
            in1 => \N__39126\,
            in2 => \_gnd_net_\,
            in3 => \N__39103\,
            lcout => \delay_measurement_inst.delay_hc_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47983\,
            ce => 'H',
            sr => \N__47274\
        );

    \delay_measurement_inst.start_timer_tr_LC_15_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001100110"
        )
    port map (
            in0 => \N__36534\,
            in1 => \N__36508\,
            in2 => \_gnd_net_\,
            in3 => \N__36489\,
            lcout => \delay_measurement_inst.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47983\,
            ce => 'H',
            sr => \N__47274\
        );

    \delay_measurement_inst.stop_timer_tr_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__36536\,
            in1 => \N__36512\,
            in2 => \N__47465\,
            in3 => \N__36490\,
            lcout => \delay_measurement_inst.stop_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47975\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_DELAY_HC1_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36473\,
            lcout => delay_hc_d1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47975\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_DELAY_HC2_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36458\,
            lcout => delay_hc_d2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47975\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_9_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011111111"
        )
    port map (
            in0 => \N__40693\,
            in1 => \N__44078\,
            in2 => \N__36413\,
            in3 => \N__36704\,
            lcout => measured_delay_hc_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47966\,
            ce => 'H',
            sr => \N__47286\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__36645\,
            in1 => \N__36364\,
            in2 => \_gnd_net_\,
            in3 => \N__36596\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_338_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__36597\,
            in1 => \N__36365\,
            in2 => \_gnd_net_\,
            in3 => \N__36646\,
            lcout => \delay_measurement_inst.delay_tr_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47966\,
            ce => 'H',
            sr => \N__47286\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOKRB1_10_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__44355\,
            in1 => \N__44257\,
            in2 => \N__41554\,
            in3 => \N__42432\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITLCJ3_7_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__36629\,
            in1 => \N__41643\,
            in2 => \N__36650\,
            in3 => \N__41707\,
            lcout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36647\,
            in2 => \_gnd_net_\,
            in3 => \N__36598\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_337_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_15_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__44080\,
            in1 => \N__44138\,
            in2 => \N__42010\,
            in3 => \N__44020\,
            lcout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINVQV2_14_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100000000"
        )
    port map (
            in0 => \N__42369\,
            in1 => \N__44081\,
            in2 => \N__36833\,
            in3 => \N__44149\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt15_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINAE19_13_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000000000000"
        )
    port map (
            in0 => \N__36620\,
            in1 => \N__36614\,
            in2 => \N__39380\,
            in3 => \N__39365\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOVQ9D_15_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000011110000"
        )
    port map (
            in0 => \N__36608\,
            in1 => \N__42011\,
            in2 => \N__36602\,
            in3 => \N__43956\,
            lcout => \delay_measurement_inst.un1_elapsed_time_hc\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36599\,
            lcout => \delay_measurement_inst.delay_tr_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIB9F91_3_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111111111"
        )
    port map (
            in0 => \N__42470\,
            in1 => \N__42431\,
            in2 => \_gnd_net_\,
            in3 => \N__44014\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto6_c_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIEB452_7_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41638\,
            in2 => \N__36851\,
            in3 => \N__41705\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto6_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINH8A4_6_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101000001010"
        )
    port map (
            in0 => \N__44079\,
            in1 => \N__42391\,
            in2 => \N__36848\,
            in3 => \N__44015\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJHF91_7_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__41706\,
            in1 => \_gnd_net_\,
            in2 => \N__41645\,
            in3 => \N__44016\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI64F91_1_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__41206\,
            in1 => \N__44356\,
            in2 => \_gnd_net_\,
            in3 => \N__41272\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_26_1_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__36824\,
            in1 => \N__36762\,
            in2 => \N__36728\,
            in3 => \N__36741\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_20_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__36763\,
            in1 => \N__40681\,
            in2 => \_gnd_net_\,
            in3 => \N__36696\,
            lcout => measured_delay_hc_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47940\,
            ce => 'H',
            sr => \N__47300\
        );

    \delay_measurement_inst.delay_hc_reg_19_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111100010"
        )
    port map (
            in0 => \N__36742\,
            in1 => \N__40684\,
            in2 => \N__44261\,
            in3 => \N__40792\,
            lcout => measured_delay_hc_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47940\,
            ce => 'H',
            sr => \N__47300\
        );

    \delay_measurement_inst.delay_hc_reg_22_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__40793\,
            in1 => \_gnd_net_\,
            in2 => \N__40721\,
            in3 => \N__36723\,
            lcout => measured_delay_hc_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47940\,
            ce => 'H',
            sr => \N__47300\
        );

    \delay_measurement_inst.delay_hc_reg_29_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__37076\,
            in1 => \N__40683\,
            in2 => \_gnd_net_\,
            in3 => \N__36697\,
            lcout => measured_delay_hc_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47940\,
            ce => 'H',
            sr => \N__47300\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_4_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__37075\,
            in1 => \N__39619\,
            in2 => \N__37058\,
            in3 => \N__39607\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_27_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__37057\,
            in1 => \N__40682\,
            in2 => \_gnd_net_\,
            in3 => \N__40794\,
            lcout => measured_delay_hc_27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47940\,
            ce => 'H',
            sr => \N__47300\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37043\,
            in2 => \N__37037\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_13_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37010\,
            in2 => \_gnd_net_\,
            in3 => \N__36983\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36980\,
            in2 => \N__36968\,
            in3 => \N__36947\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36944\,
            in2 => \_gnd_net_\,
            in3 => \N__36911\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36908\,
            in2 => \_gnd_net_\,
            in3 => \N__36878\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36875\,
            in2 => \_gnd_net_\,
            in3 => \N__36854\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37238\,
            in2 => \_gnd_net_\,
            in3 => \N__37208\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37205\,
            in2 => \_gnd_net_\,
            in3 => \N__37184\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37181\,
            in2 => \_gnd_net_\,
            in3 => \N__37157\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_15_14_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40300\,
            in2 => \_gnd_net_\,
            in3 => \N__37154\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37151\,
            in2 => \_gnd_net_\,
            in3 => \N__37124\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37121\,
            in2 => \_gnd_net_\,
            in3 => \N__37103\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40279\,
            in2 => \_gnd_net_\,
            in3 => \N__37100\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37097\,
            in2 => \_gnd_net_\,
            in3 => \N__37079\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40258\,
            in2 => \_gnd_net_\,
            in3 => \N__37376\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37372\,
            in2 => \_gnd_net_\,
            in3 => \N__37349\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37345\,
            in2 => \_gnd_net_\,
            in3 => \N__37325\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \bfn_15_15_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37322\,
            in2 => \_gnd_net_\,
            in3 => \N__37301\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39832\,
            in2 => \_gnd_net_\,
            in3 => \N__37298\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0_c_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__37295\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_16_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37274\,
            in2 => \N__37286\,
            in3 => \N__45327\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37259\,
            in2 => \N__37268\,
            in3 => \N__45295\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37244\,
            in2 => \N__37253\,
            in3 => \N__45253\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37481\,
            in2 => \N__37490\,
            in3 => \N__45220\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37466\,
            in2 => \N__37475\,
            in3 => \N__45187\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37451\,
            in2 => \N__37460\,
            in3 => \N__45151\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__45643\,
            in1 => \N__37436\,
            in2 => \N__37445\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37418\,
            in2 => \N__37430\,
            in3 => \N__45610\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \bfn_15_17_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37400\,
            in2 => \N__37412\,
            in3 => \N__45581\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37382\,
            in2 => \N__37394\,
            in3 => \N__45547\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37628\,
            in2 => \N__37643\,
            in3 => \N__45518\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37610\,
            in2 => \N__37622\,
            in3 => \N__45491\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37592\,
            in2 => \N__37604\,
            in3 => \N__45464\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__45889\,
            in1 => \N__37571\,
            in2 => \N__37586\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37553\,
            in2 => \N__37565\,
            in3 => \N__45863\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37532\,
            in2 => \N__37547\,
            in3 => \N__45836\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \bfn_15_18_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37511\,
            in2 => \N__37526\,
            in3 => \N__45809\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37496\,
            in2 => \N__37505\,
            in3 => \N__45782\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37703\,
            in2 => \N__37697\,
            in3 => \N__45755\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37688\,
            lcout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1B6_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38191\,
            in2 => \_gnd_net_\,
            in3 => \N__38681\,
            lcout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__43063\,
            in1 => \N__45328\,
            in2 => \_gnd_net_\,
            in3 => \N__43015\,
            lcout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_7_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010100010"
        )
    port map (
            in0 => \N__37667\,
            in1 => \N__37841\,
            in2 => \N__38131\,
            in3 => \N__37938\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47893\,
            ce => 'H',
            sr => \N__47355\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_8_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__37840\,
            in1 => \N__38106\,
            in2 => \N__37978\,
            in3 => \N__37661\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47893\,
            ce => 'H',
            sr => \N__47355\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_9_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__37839\,
            in1 => \N__37934\,
            in2 => \N__38130\,
            in3 => \N__37655\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47893\,
            ce => 'H',
            sr => \N__47355\
        );

    \phase_controller_slave.stoper_tr.stoper_state_RNII60D_0_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__37933\,
            in1 => \N__37838\,
            in2 => \_gnd_net_\,
            in3 => \N__38105\,
            lcout => \phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38190\,
            in2 => \_gnd_net_\,
            in3 => \N__38680\,
            lcout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_10_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__37858\,
            in1 => \N__38123\,
            in2 => \N__38009\,
            in3 => \N__38198\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47886\,
            ce => 'H',
            sr => \N__47364\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__38192\,
            in1 => \N__37729\,
            in2 => \_gnd_net_\,
            in3 => \N__38682\,
            lcout => OPEN,
            ltout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_1_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__37861\,
            in1 => \N__38007\,
            in2 => \N__38159\,
            in3 => \N__38129\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47886\,
            ce => 'H',
            sr => \N__47364\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_11_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010100010"
        )
    port map (
            in0 => \N__38156\,
            in1 => \N__37979\,
            in2 => \N__38132\,
            in3 => \N__37862\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47886\,
            ce => 'H',
            sr => \N__47364\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_12_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__37859\,
            in1 => \N__38124\,
            in2 => \N__38010\,
            in3 => \N__38150\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47886\,
            ce => 'H',
            sr => \N__47364\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_13_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__38121\,
            in1 => \N__37980\,
            in2 => \N__37873\,
            in3 => \N__38144\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47886\,
            ce => 'H',
            sr => \N__47364\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_14_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__37860\,
            in1 => \N__38125\,
            in2 => \N__38011\,
            in3 => \N__38138\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47886\,
            ce => 'H',
            sr => \N__47364\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_15_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__38122\,
            in1 => \N__37981\,
            in2 => \N__37874\,
            in3 => \N__37739\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47886\,
            ce => 'H',
            sr => \N__47364\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37709\,
            in2 => \N__40892\,
            in3 => \N__37725\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_15_21_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38366\,
            in2 => \N__40910\,
            in3 => \N__38377\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38342\,
            in2 => \N__41006\,
            in3 => \N__38353\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38321\,
            in2 => \N__40862\,
            in3 => \N__38332\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38300\,
            in2 => \N__40997\,
            in3 => \N__38311\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38276\,
            in2 => \N__40883\,
            in3 => \N__38287\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38255\,
            in2 => \N__40871\,
            in3 => \N__38270\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38225\,
            in2 => \N__38249\,
            in3 => \N__38240\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38204\,
            in2 => \N__40937\,
            in3 => \N__38219\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_15_22_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38549\,
            in1 => \N__38534\,
            in2 => \N__40985\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38513\,
            in2 => \N__40973\,
            in3 => \N__38528\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38492\,
            in2 => \N__40949\,
            in3 => \N__38507\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38486\,
            in1 => \N__38471\,
            in2 => \N__40958\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38450\,
            in2 => \N__43373\,
            in3 => \N__38465\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_15_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38444\,
            in1 => \N__40898\,
            in2 => \N__38429\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38387\,
            in2 => \N__38420\,
            in3 => \N__38408\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38753\,
            in2 => \N__38642\,
            in3 => \N__38771\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_15_23_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38729\,
            in2 => \N__38633\,
            in3 => \N__38747\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_15_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38723\,
            in1 => \N__38708\,
            in2 => \N__40928\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38702\,
            lcout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.target_time_17_LC_15_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48373\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47872\,
            ce => \N__43353\,
            sr => \N__47385\
        );

    \phase_controller_slave.stoper_tr.target_time_18_LC_15_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48409\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47872\,
            ce => \N__43353\,
            sr => \N__47385\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_15_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38597\,
            in2 => \N__41114\,
            in3 => \N__38613\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_15_24_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_15_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40919\,
            in2 => \N__38579\,
            in3 => \N__38590\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_15_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38555\,
            in2 => \N__41129\,
            in3 => \N__38566\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_15_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38897\,
            in2 => \N__41141\,
            in3 => \N__38908\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_15_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38890\,
            in1 => \N__38879\,
            in2 => \N__41036\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_15_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41147\,
            in2 => \N__38861\,
            in3 => \N__38872\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_15_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38851\,
            in1 => \N__38840\,
            in2 => \N__41105\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_15_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38833\,
            in1 => \N__38822\,
            in2 => \N__41045\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_15_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38795\,
            in2 => \N__41339\,
            in3 => \N__38812\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_15_25_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_15_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38788\,
            in1 => \N__38777\,
            in2 => \N__41057\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_15_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39062\,
            in2 => \N__41090\,
            in3 => \N__39073\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_15_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__39055\,
            in1 => \N__39044\,
            in2 => \N__41288\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_15_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39026\,
            in2 => \N__41330\,
            in3 => \N__39037\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_15_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39008\,
            in2 => \N__41321\,
            in3 => \N__39019\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_15_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43136\,
            in2 => \N__38990\,
            in3 => \N__39001\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_15_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38951\,
            in2 => \N__38981\,
            in3 => \N__38969\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_15_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38933\,
            in2 => \N__39167\,
            in3 => \N__38944\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_15_26_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_15_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38915\,
            in2 => \N__39158\,
            in3 => \N__38926\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_15_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39230\,
            in2 => \N__39149\,
            in3 => \N__39241\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_15_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39224\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_17_LC_15_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48377\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47856\,
            ce => \N__43103\,
            sr => \N__47401\
        );

    \phase_controller_inst1.stoper_tr.target_time_18_LC_15_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__48410\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47856\,
            ce => \N__43103\,
            sr => \N__47401\
        );

    \phase_controller_inst1.stoper_tr.target_time_19_LC_15_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48059\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47856\,
            ce => \N__43103\,
            sr => \N__47401\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_16_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__39102\,
            in1 => \N__39139\,
            in2 => \_gnd_net_\,
            in3 => \N__39128\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_336_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_16_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39101\,
            lcout => \delay_measurement_inst.delay_hc_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.counter_0_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39548\,
            in1 => \N__41247\,
            in2 => \_gnd_net_\,
            in3 => \N__39080\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_16_7_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            clk => \N__47984\,
            ce => \N__39405\,
            sr => \N__47275\
        );

    \delay_measurement_inst.delay_hc_timer.counter_1_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39504\,
            in1 => \N__44373\,
            in2 => \_gnd_net_\,
            in3 => \N__39077\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            clk => \N__47984\,
            ce => \N__39405\,
            sr => \N__47275\
        );

    \delay_measurement_inst.delay_hc_timer.counter_2_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39549\,
            in1 => \N__41226\,
            in2 => \_gnd_net_\,
            in3 => \N__39269\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            clk => \N__47984\,
            ce => \N__39405\,
            sr => \N__47275\
        );

    \delay_measurement_inst.delay_hc_timer.counter_3_LC_16_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39505\,
            in1 => \N__41169\,
            in2 => \_gnd_net_\,
            in3 => \N__39266\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            clk => \N__47984\,
            ce => \N__39405\,
            sr => \N__47275\
        );

    \delay_measurement_inst.delay_hc_timer.counter_4_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39550\,
            in1 => \N__41730\,
            in2 => \_gnd_net_\,
            in3 => \N__39263\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            clk => \N__47984\,
            ce => \N__39405\,
            sr => \N__47275\
        );

    \delay_measurement_inst.delay_hc_timer.counter_5_LC_16_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39506\,
            in1 => \N__41664\,
            in2 => \_gnd_net_\,
            in3 => \N__39260\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            clk => \N__47984\,
            ce => \N__39405\,
            sr => \N__47275\
        );

    \delay_measurement_inst.delay_hc_timer.counter_6_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39551\,
            in1 => \N__41598\,
            in2 => \_gnd_net_\,
            in3 => \N__39257\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            clk => \N__47984\,
            ce => \N__39405\,
            sr => \N__47275\
        );

    \delay_measurement_inst.delay_hc_timer.counter_7_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39507\,
            in1 => \N__41574\,
            in2 => \_gnd_net_\,
            in3 => \N__39254\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            clk => \N__47984\,
            ce => \N__39405\,
            sr => \N__47275\
        );

    \delay_measurement_inst.delay_hc_timer.counter_8_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39539\,
            in1 => \N__41514\,
            in2 => \_gnd_net_\,
            in3 => \N__39251\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_16_8_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            clk => \N__47976\,
            ce => \N__39423\,
            sr => \N__47278\
        );

    \delay_measurement_inst.delay_hc_timer.counter_9_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39517\,
            in1 => \N__41466\,
            in2 => \_gnd_net_\,
            in3 => \N__39248\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            clk => \N__47976\,
            ce => \N__39423\,
            sr => \N__47278\
        );

    \delay_measurement_inst.delay_hc_timer.counter_10_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39536\,
            in1 => \N__41415\,
            in2 => \_gnd_net_\,
            in3 => \N__39245\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            clk => \N__47976\,
            ce => \N__39423\,
            sr => \N__47278\
        );

    \delay_measurement_inst.delay_hc_timer.counter_11_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39514\,
            in1 => \N__41361\,
            in2 => \_gnd_net_\,
            in3 => \N__39296\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            clk => \N__47976\,
            ce => \N__39423\,
            sr => \N__47278\
        );

    \delay_measurement_inst.delay_hc_timer.counter_12_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39537\,
            in1 => \N__42045\,
            in2 => \_gnd_net_\,
            in3 => \N__39293\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            clk => \N__47976\,
            ce => \N__39423\,
            sr => \N__47278\
        );

    \delay_measurement_inst.delay_hc_timer.counter_13_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39515\,
            in1 => \N__41958\,
            in2 => \_gnd_net_\,
            in3 => \N__39290\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            clk => \N__47976\,
            ce => \N__39423\,
            sr => \N__47278\
        );

    \delay_measurement_inst.delay_hc_timer.counter_14_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39538\,
            in1 => \N__41934\,
            in2 => \_gnd_net_\,
            in3 => \N__39287\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            clk => \N__47976\,
            ce => \N__39423\,
            sr => \N__47278\
        );

    \delay_measurement_inst.delay_hc_timer.counter_15_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39516\,
            in1 => \N__41910\,
            in2 => \_gnd_net_\,
            in3 => \N__39284\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            clk => \N__47976\,
            ce => \N__39423\,
            sr => \N__47278\
        );

    \delay_measurement_inst.delay_hc_timer.counter_16_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39544\,
            in1 => \N__41886\,
            in2 => \_gnd_net_\,
            in3 => \N__39281\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_16_9_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            clk => \N__47967\,
            ce => \N__39425\,
            sr => \N__47287\
        );

    \delay_measurement_inst.delay_hc_timer.counter_17_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39540\,
            in1 => \N__41862\,
            in2 => \_gnd_net_\,
            in3 => \N__39278\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            clk => \N__47967\,
            ce => \N__39425\,
            sr => \N__47287\
        );

    \delay_measurement_inst.delay_hc_timer.counter_18_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39545\,
            in1 => \N__41820\,
            in2 => \_gnd_net_\,
            in3 => \N__39275\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            clk => \N__47967\,
            ce => \N__39425\,
            sr => \N__47287\
        );

    \delay_measurement_inst.delay_hc_timer.counter_19_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39541\,
            in1 => \N__41775\,
            in2 => \_gnd_net_\,
            in3 => \N__39272\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            clk => \N__47967\,
            ce => \N__39425\,
            sr => \N__47287\
        );

    \delay_measurement_inst.delay_hc_timer.counter_20_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39546\,
            in1 => \N__42318\,
            in2 => \_gnd_net_\,
            in3 => \N__39323\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            clk => \N__47967\,
            ce => \N__39425\,
            sr => \N__47287\
        );

    \delay_measurement_inst.delay_hc_timer.counter_21_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39542\,
            in1 => \N__42288\,
            in2 => \_gnd_net_\,
            in3 => \N__39320\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            clk => \N__47967\,
            ce => \N__39425\,
            sr => \N__47287\
        );

    \delay_measurement_inst.delay_hc_timer.counter_22_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39547\,
            in1 => \N__42258\,
            in2 => \_gnd_net_\,
            in3 => \N__39317\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            clk => \N__47967\,
            ce => \N__39425\,
            sr => \N__47287\
        );

    \delay_measurement_inst.delay_hc_timer.counter_23_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39543\,
            in1 => \N__42228\,
            in2 => \_gnd_net_\,
            in3 => \N__39314\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            clk => \N__47967\,
            ce => \N__39425\,
            sr => \N__47287\
        );

    \delay_measurement_inst.delay_hc_timer.counter_24_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39508\,
            in1 => \N__42198\,
            in2 => \_gnd_net_\,
            in3 => \N__39311\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_16_10_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            clk => \N__47959\,
            ce => \N__39424\,
            sr => \N__47290\
        );

    \delay_measurement_inst.delay_hc_timer.counter_25_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39512\,
            in1 => \N__42168\,
            in2 => \_gnd_net_\,
            in3 => \N__39308\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            clk => \N__47959\,
            ce => \N__39424\,
            sr => \N__47290\
        );

    \delay_measurement_inst.delay_hc_timer.counter_26_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39509\,
            in1 => \N__42138\,
            in2 => \_gnd_net_\,
            in3 => \N__39305\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            clk => \N__47959\,
            ce => \N__39424\,
            sr => \N__47290\
        );

    \delay_measurement_inst.delay_hc_timer.counter_27_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39513\,
            in1 => \N__42093\,
            in2 => \_gnd_net_\,
            in3 => \N__39302\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            clk => \N__47959\,
            ce => \N__39424\,
            sr => \N__47290\
        );

    \delay_measurement_inst.delay_hc_timer.counter_28_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39510\,
            in1 => \N__42118\,
            in2 => \_gnd_net_\,
            in3 => \N__39299\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_28\,
            clk => \N__47959\,
            ce => \N__39424\,
            sr => \N__47290\
        );

    \delay_measurement_inst.delay_hc_timer.counter_29_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__42073\,
            in1 => \N__39511\,
            in2 => \_gnd_net_\,
            in3 => \N__39428\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47959\,
            ce => \N__39424\,
            sr => \N__47290\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVU8G_23_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42269\,
            in2 => \_gnd_net_\,
            in3 => \N__42299\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBC512_25_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__42209\,
            in1 => \N__42239\,
            in2 => \N__39389\,
            in3 => \N__39371\,
            lcout => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII0UL_14_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__44071\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44134\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_a1_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJHOP1_7_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100000"
        )
    port map (
            in0 => \N__41698\,
            in1 => \N__41642\,
            in2 => \N__39386\,
            in3 => \N__44182\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_a1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRLFA3_15_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010000000000"
        )
    port map (
            in0 => \N__44184\,
            in1 => \N__42012\,
            in2 => \N__39383\,
            in3 => \N__43950\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILLI01_20_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41797\,
            in1 => \N__41836\,
            in2 => \N__41752\,
            in3 => \N__44183\,
            lcout => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__42104\,
            in1 => \N__42149\,
            in2 => \N__42059\,
            in3 => \N__42179\,
            lcout => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JIP2_20_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__39364\,
            in1 => \N__41756\,
            in2 => \N__41843\,
            in3 => \N__41801\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto30_2\,
            ltout => \delay_measurement_inst.delay_hc_reg3lto30_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVBSED_31_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101011"
        )
    port map (
            in0 => \N__39779\,
            in1 => \N__44185\,
            in2 => \N__39773\,
            in3 => \N__42344\,
            lcout => \delay_measurement_inst.delay_hc_reg3\,
            ltout => \delay_measurement_inst.delay_hc_reg3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_4_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__40702\,
            in1 => \N__42474\,
            in2 => \N__39770\,
            in3 => \N__39758\,
            lcout => measured_delay_hc_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47950\,
            ce => 'H',
            sr => \N__47294\
        );

    \delay_measurement_inst.delay_hc_reg_14_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111011000"
        )
    port map (
            in0 => \N__40697\,
            in1 => \N__44145\,
            in2 => \N__39712\,
            in3 => \N__40785\,
            lcout => measured_delay_hc_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47941\,
            ce => 'H',
            sr => \N__47301\
        );

    \delay_measurement_inst.delay_hc_reg_24_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__40786\,
            in1 => \N__40698\,
            in2 => \_gnd_net_\,
            in3 => \N__39673\,
            lcout => measured_delay_hc_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47941\,
            ce => 'H',
            sr => \N__47301\
        );

    \delay_measurement_inst.delay_hc_reg_25_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__40695\,
            in1 => \N__39655\,
            in2 => \_gnd_net_\,
            in3 => \N__40787\,
            lcout => measured_delay_hc_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47941\,
            ce => 'H',
            sr => \N__47301\
        );

    \delay_measurement_inst.delay_hc_reg_26_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__40788\,
            in1 => \N__40699\,
            in2 => \_gnd_net_\,
            in3 => \N__39634\,
            lcout => measured_delay_hc_26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47941\,
            ce => 'H',
            sr => \N__47301\
        );

    \delay_measurement_inst.delay_hc_reg_28_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__40696\,
            in1 => \N__39620\,
            in2 => \_gnd_net_\,
            in3 => \N__40789\,
            lcout => measured_delay_hc_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47941\,
            ce => 'H',
            sr => \N__47301\
        );

    \delay_measurement_inst.delay_hc_reg_30_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__40790\,
            in1 => \N__40700\,
            in2 => \_gnd_net_\,
            in3 => \N__39608\,
            lcout => measured_delay_hc_30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47941\,
            ce => 'H',
            sr => \N__47301\
        );

    \delay_measurement_inst.delay_hc_reg_0_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__40694\,
            in1 => \N__39581\,
            in2 => \_gnd_net_\,
            in3 => \N__40784\,
            lcout => measured_delay_hc_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47941\,
            ce => 'H',
            sr => \N__47301\
        );

    \delay_measurement_inst.delay_hc_reg_31_LC_16_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__40791\,
            in1 => \N__40701\,
            in2 => \_gnd_net_\,
            in3 => \N__40358\,
            lcout => measured_delay_hc_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47941\,
            ce => 'H',
            sr => \N__47301\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010000100"
        )
    port map (
            in0 => \N__39962\,
            in1 => \N__40307\,
            in2 => \N__40120\,
            in3 => \N__40244\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47930\,
            ce => 'H',
            sr => \N__47307\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__39963\,
            in1 => \N__40242\,
            in2 => \N__40121\,
            in3 => \N__40286\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47930\,
            ce => 'H',
            sr => \N__47307\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__39964\,
            in1 => \N__40243\,
            in2 => \N__40122\,
            in3 => \N__40265\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47930\,
            ce => 'H',
            sr => \N__47307\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__40241\,
            in1 => \N__40090\,
            in2 => \N__39974\,
            in3 => \N__39965\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47930\,
            ce => 'H',
            sr => \N__47307\
        );

    \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_0_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__43714\,
            in1 => \N__43583\,
            in2 => \_gnd_net_\,
            in3 => \N__43852\,
            lcout => \phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_7_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__43854\,
            in1 => \N__43584\,
            in2 => \N__43724\,
            in3 => \N__45632\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47916\,
            ce => 'H',
            sr => \N__47320\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_2_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__43823\,
            in1 => \N__43558\,
            in2 => \N__43721\,
            in3 => \N__45284\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47912\,
            ce => 'H',
            sr => \N__47326\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_8_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__43556\,
            in1 => \N__43703\,
            in2 => \N__45599\,
            in3 => \N__43829\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47912\,
            ce => 'H',
            sr => \N__47326\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_3_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__43824\,
            in1 => \N__43559\,
            in2 => \N__43722\,
            in3 => \N__45242\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47912\,
            ce => 'H',
            sr => \N__47326\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_5_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__43554\,
            in1 => \N__43701\,
            in2 => \N__45176\,
            in3 => \N__43827\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47912\,
            ce => 'H',
            sr => \N__47326\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_14_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__43822\,
            in1 => \N__43557\,
            in2 => \N__43720\,
            in3 => \N__45878\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47912\,
            ce => 'H',
            sr => \N__47326\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_6_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__43555\,
            in1 => \N__43702\,
            in2 => \N__45668\,
            in3 => \N__43828\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47912\,
            ce => 'H',
            sr => \N__47326\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_4_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__43825\,
            in1 => \N__43560\,
            in2 => \N__43723\,
            in3 => \N__45209\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47912\,
            ce => 'H',
            sr => \N__47326\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_10_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__43553\,
            in1 => \N__43700\,
            in2 => \N__45536\,
            in3 => \N__43826\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47912\,
            ce => 'H',
            sr => \N__47326\
        );

    \phase_controller_slave.stoper_hc.stoper_state_RNIDEUE_0_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43564\,
            in2 => \_gnd_net_\,
            in3 => \N__43834\,
            lcout => \phase_controller_slave.stoper_hc.time_passed11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__43835\,
            in1 => \_gnd_net_\,
            in2 => \N__43586\,
            in3 => \N__43660\,
            lcout => \phase_controller_slave.stoper_hc.time_passed_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_esr_10_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__48260\,
            in1 => \N__48505\,
            in2 => \_gnd_net_\,
            in3 => \N__45950\,
            lcout => measured_delay_tr_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47900\,
            ce => \N__47518\,
            sr => \N__47348\
        );

    \delay_measurement_inst.delay_tr_reg_esr_12_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__48506\,
            in1 => \N__48261\,
            in2 => \_gnd_net_\,
            in3 => \N__45968\,
            lcout => measured_delay_tr_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47900\,
            ce => \N__47518\,
            sr => \N__47348\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_6_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41304\,
            in1 => \N__48459\,
            in2 => \N__46678\,
            in3 => \N__41073\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_9_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40913\,
            in3 => \N__41019\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_esr_9_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000100"
        )
    port map (
            in0 => \N__42932\,
            in1 => \N__48504\,
            in2 => \N__48281\,
            in3 => \N__46034\,
            lcout => measured_delay_tr_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47894\,
            ce => \N__47519\,
            sr => \N__47356\
        );

    \phase_controller_slave.stoper_tr.target_time_2_LC_16_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__43244\,
            in1 => \N__43186\,
            in2 => \N__46432\,
            in3 => \N__43407\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47887\,
            ce => \N__43352\,
            sr => \N__47365\
        );

    \phase_controller_slave.stoper_tr.target_time_15_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45712\,
            in2 => \_gnd_net_\,
            in3 => \N__46182\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47887\,
            ce => \N__43352\,
            sr => \N__47365\
        );

    \phase_controller_slave.stoper_tr.target_time_1_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101011101010"
        )
    port map (
            in0 => \N__43243\,
            in1 => \N__43185\,
            in2 => \N__46060\,
            in3 => \N__43406\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47887\,
            ce => \N__43352\,
            sr => \N__47365\
        );

    \phase_controller_slave.stoper_tr.target_time_6_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__43411\,
            in1 => \N__46615\,
            in2 => \_gnd_net_\,
            in3 => \N__43190\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47887\,
            ce => \N__43352\,
            sr => \N__47365\
        );

    \phase_controller_slave.stoper_tr.target_time_7_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46759\,
            in2 => \_gnd_net_\,
            in3 => \N__43412\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47887\,
            ce => \N__43352\,
            sr => \N__47365\
        );

    \phase_controller_slave.stoper_tr.target_time_4_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__43409\,
            in1 => \N__43188\,
            in2 => \_gnd_net_\,
            in3 => \N__46564\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47887\,
            ce => \N__43352\,
            sr => \N__47365\
        );

    \phase_controller_slave.stoper_tr.target_time_3_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__43187\,
            in1 => \N__43408\,
            in2 => \N__46888\,
            in3 => \N__43263\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47887\,
            ce => \N__43352\,
            sr => \N__47365\
        );

    \phase_controller_slave.stoper_tr.target_time_5_LC_16_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__43410\,
            in1 => \N__43189\,
            in2 => \_gnd_net_\,
            in3 => \N__46945\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47887\,
            ce => \N__43352\,
            sr => \N__47365\
        );

    \phase_controller_slave.stoper_tr.target_time_10_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43299\,
            in2 => \_gnd_net_\,
            in3 => \N__41080\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47883\,
            ce => \N__43348\,
            sr => \N__47374\
        );

    \phase_controller_slave.stoper_tr.target_time_11_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__43300\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48466\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47883\,
            ce => \N__43348\,
            sr => \N__47374\
        );

    \phase_controller_slave.stoper_tr.target_time_13_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__43302\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46674\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47883\,
            ce => \N__43348\,
            sr => \N__47374\
        );

    \phase_controller_slave.stoper_tr.target_time_12_LC_16_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__41311\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43301\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47883\,
            ce => \N__43348\,
            sr => \N__47374\
        );

    \phase_controller_slave.stoper_tr.target_time_9_LC_16_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110011011101"
        )
    port map (
            in0 => \N__43303\,
            in1 => \N__41027\,
            in2 => \N__46184\,
            in3 => \N__43218\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47883\,
            ce => \N__43348\,
            sr => \N__47374\
        );

    \phase_controller_slave.stoper_tr.target_time_19_LC_16_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48054\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47883\,
            ce => \N__43348\,
            sr => \N__47374\
        );

    \phase_controller_inst1.stoper_tr.target_time_2_LC_16_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011100000"
        )
    port map (
            in0 => \N__43161\,
            in1 => \N__43435\,
            in2 => \N__46433\,
            in3 => \N__43237\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47880\,
            ce => \N__43094\,
            sr => \N__47380\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__43438\,
            in1 => \N__43164\,
            in2 => \_gnd_net_\,
            in3 => \N__46619\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47880\,
            ce => \N__43094\,
            sr => \N__47380\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_LC_16_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__43163\,
            in1 => \N__46568\,
            in2 => \_gnd_net_\,
            in3 => \N__43437\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47880\,
            ce => \N__43094\,
            sr => \N__47380\
        );

    \phase_controller_inst1.stoper_tr.target_time_3_LC_16_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__43436\,
            in1 => \N__43162\,
            in2 => \N__46889\,
            in3 => \N__43265\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47880\,
            ce => \N__43094\,
            sr => \N__47380\
        );

    \phase_controller_inst1.stoper_tr.target_time_1_LC_16_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__43160\,
            in1 => \N__43434\,
            in2 => \N__46067\,
            in3 => \N__43236\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47880\,
            ce => \N__43094\,
            sr => \N__47380\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_LC_16_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43440\,
            in2 => \_gnd_net_\,
            in3 => \N__46763\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47873\,
            ce => \N__43110\,
            sr => \N__47386\
        );

    \phase_controller_inst1.stoper_tr.target_time_11_LC_16_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__43297\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48467\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47873\,
            ce => \N__43110\,
            sr => \N__47386\
        );

    \phase_controller_inst1.stoper_tr.target_time_10_LC_16_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43296\,
            in2 => \_gnd_net_\,
            in3 => \N__41081\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47873\,
            ce => \N__43110\,
            sr => \N__47386\
        );

    \phase_controller_inst1.stoper_tr.target_time_8_LC_16_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__43441\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46822\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47873\,
            ce => \N__43110\,
            sr => \N__47386\
        );

    \phase_controller_inst1.stoper_tr.target_time_5_LC_16_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__43165\,
            in1 => \N__46946\,
            in2 => \_gnd_net_\,
            in3 => \N__43439\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47873\,
            ce => \N__43110\,
            sr => \N__47386\
        );

    \phase_controller_inst1.stoper_tr.target_time_9_LC_16_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111101000101"
        )
    port map (
            in0 => \N__43298\,
            in1 => \N__46183\,
            in2 => \N__43223\,
            in3 => \N__41026\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47873\,
            ce => \N__43110\,
            sr => \N__47386\
        );

    \phase_controller_inst1.stoper_tr.target_time_13_LC_16_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__43310\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46679\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47867\,
            ce => \N__43123\,
            sr => \N__47394\
        );

    \phase_controller_inst1.stoper_tr.target_time_14_LC_16_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__45713\,
            in1 => \N__46181\,
            in2 => \_gnd_net_\,
            in3 => \N__46318\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47867\,
            ce => \N__43123\,
            sr => \N__47394\
        );

    \phase_controller_inst1.stoper_tr.target_time_12_LC_16_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43309\,
            in2 => \_gnd_net_\,
            in3 => \N__41312\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47867\,
            ce => \N__43123\,
            sr => \N__47394\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41249\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.elapsed_time_hc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47991\,
            ce => \N__44328\,
            sr => \N__47272\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41248\,
            in2 => \N__41228\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.elapsed_time_hc_3\,
            ltout => OPEN,
            carryin => \bfn_17_8_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__47985\,
            ce => \N__44329\,
            sr => \N__47276\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44374\,
            in2 => \N__41171\,
            in3 => \N__41231\,
            lcout => \delay_measurement_inst.elapsed_time_hc_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__47985\,
            ce => \N__44329\,
            sr => \N__47276\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41227\,
            in2 => \N__41732\,
            in3 => \N__41174\,
            lcout => \delay_measurement_inst.elapsed_time_hc_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__47985\,
            ce => \N__44329\,
            sr => \N__47276\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41170\,
            in2 => \N__41666\,
            in3 => \N__41150\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__47985\,
            ce => \N__44329\,
            sr => \N__47276\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41731\,
            in2 => \N__41600\,
            in3 => \N__41669\,
            lcout => \delay_measurement_inst.elapsed_time_hc_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__47985\,
            ce => \N__44329\,
            sr => \N__47276\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41665\,
            in2 => \N__41576\,
            in3 => \N__41603\,
            lcout => \delay_measurement_inst.elapsed_time_hc_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__47985\,
            ce => \N__44329\,
            sr => \N__47276\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41599\,
            in2 => \N__41516\,
            in3 => \N__41579\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__47985\,
            ce => \N__44329\,
            sr => \N__47276\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41575\,
            in2 => \N__41468\,
            in3 => \N__41519\,
            lcout => \delay_measurement_inst.elapsed_time_hc_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__47985\,
            ce => \N__44329\,
            sr => \N__47276\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41515\,
            in2 => \N__41417\,
            in3 => \N__41471\,
            lcout => \delay_measurement_inst.elapsed_time_hc_11\,
            ltout => OPEN,
            carryin => \bfn_17_9_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__47977\,
            ce => \N__44330\,
            sr => \N__47279\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41467\,
            in2 => \N__41363\,
            in3 => \N__41420\,
            lcout => \delay_measurement_inst.elapsed_time_hc_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__47977\,
            ce => \N__44330\,
            sr => \N__47279\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41416\,
            in2 => \N__42047\,
            in3 => \N__41366\,
            lcout => \delay_measurement_inst.elapsed_time_hc_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__47977\,
            ce => \N__44330\,
            sr => \N__47279\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41362\,
            in2 => \N__41960\,
            in3 => \N__41342\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__47977\,
            ce => \N__44330\,
            sr => \N__47279\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42046\,
            in2 => \N__41936\,
            in3 => \N__41963\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__47977\,
            ce => \N__44330\,
            sr => \N__47279\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41959\,
            in2 => \N__41912\,
            in3 => \N__41939\,
            lcout => \delay_measurement_inst.elapsed_time_hc_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__47977\,
            ce => \N__44330\,
            sr => \N__47279\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41935\,
            in2 => \N__41888\,
            in3 => \N__41915\,
            lcout => \delay_measurement_inst.elapsed_time_hc_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__47977\,
            ce => \N__44330\,
            sr => \N__47279\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41911\,
            in2 => \N__41864\,
            in3 => \N__41891\,
            lcout => \delay_measurement_inst.elapsed_time_hc_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__47977\,
            ce => \N__44330\,
            sr => \N__47279\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41887\,
            in2 => \N__41822\,
            in3 => \N__41867\,
            lcout => \delay_measurement_inst.elapsed_time_hc_19\,
            ltout => OPEN,
            carryin => \bfn_17_10_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__47968\,
            ce => \N__44331\,
            sr => \N__47288\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41863\,
            in2 => \N__41777\,
            in3 => \N__41825\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__47968\,
            ce => \N__44331\,
            sr => \N__47288\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41821\,
            in2 => \N__42320\,
            in3 => \N__41780\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__47968\,
            ce => \N__44331\,
            sr => \N__47288\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41776\,
            in2 => \N__42290\,
            in3 => \N__41735\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__47968\,
            ce => \N__44331\,
            sr => \N__47288\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42319\,
            in2 => \N__42260\,
            in3 => \N__42293\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__47968\,
            ce => \N__44331\,
            sr => \N__47288\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42289\,
            in2 => \N__42230\,
            in3 => \N__42263\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__47968\,
            ce => \N__44331\,
            sr => \N__47288\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42259\,
            in2 => \N__42200\,
            in3 => \N__42233\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__47968\,
            ce => \N__44331\,
            sr => \N__47288\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42229\,
            in2 => \N__42170\,
            in3 => \N__42203\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__47968\,
            ce => \N__44331\,
            sr => \N__47288\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42199\,
            in2 => \N__42140\,
            in3 => \N__42173\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\,
            ltout => OPEN,
            carryin => \bfn_17_11_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__47960\,
            ce => \N__44333\,
            sr => \N__47291\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42169\,
            in2 => \N__42095\,
            in3 => \N__42143\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__47960\,
            ce => \N__44333\,
            sr => \N__47291\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42139\,
            in2 => \N__42119\,
            in3 => \N__42098\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__47960\,
            ce => \N__44333\,
            sr => \N__47291\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42094\,
            in2 => \N__42074\,
            in3 => \N__42050\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hcZ0Z_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__47960\,
            ce => \N__44333\,
            sr => \N__47291\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42479\,
            lcout => \delay_measurement_inst.elapsed_time_hc_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47960\,
            ce => \N__44333\,
            sr => \N__47291\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIB3GH4_3_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__42476\,
            in1 => \N__42437\,
            in2 => \N__42401\,
            in3 => \N__43907\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIB3GH4Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4KK27_3_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__44090\,
            in1 => \N__42379\,
            in2 => \N__42347\,
            in3 => \N__43943\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42717\,
            in1 => \N__43896\,
            in2 => \_gnd_net_\,
            in3 => \N__42338\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_17_13_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            clk => \N__47951\,
            ce => \N__42590\,
            sr => \N__47295\
        );

    \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42733\,
            in1 => \N__43875\,
            in2 => \_gnd_net_\,
            in3 => \N__42335\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            clk => \N__47951\,
            ce => \N__42590\,
            sr => \N__47295\
        );

    \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42718\,
            in1 => \N__44619\,
            in2 => \_gnd_net_\,
            in3 => \N__42332\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            clk => \N__47951\,
            ce => \N__42590\,
            sr => \N__47295\
        );

    \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42734\,
            in1 => \N__44592\,
            in2 => \_gnd_net_\,
            in3 => \N__42329\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            clk => \N__47951\,
            ce => \N__42590\,
            sr => \N__47295\
        );

    \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42719\,
            in1 => \N__44566\,
            in2 => \_gnd_net_\,
            in3 => \N__42326\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            clk => \N__47951\,
            ce => \N__42590\,
            sr => \N__47295\
        );

    \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42735\,
            in1 => \N__44542\,
            in2 => \_gnd_net_\,
            in3 => \N__42323\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            clk => \N__47951\,
            ce => \N__42590\,
            sr => \N__47295\
        );

    \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42716\,
            in1 => \N__44514\,
            in2 => \_gnd_net_\,
            in3 => \N__42506\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            clk => \N__47951\,
            ce => \N__42590\,
            sr => \N__47295\
        );

    \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42736\,
            in1 => \N__44482\,
            in2 => \_gnd_net_\,
            in3 => \N__42503\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            clk => \N__47951\,
            ce => \N__42590\,
            sr => \N__47295\
        );

    \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42711\,
            in1 => \N__44457\,
            in2 => \_gnd_net_\,
            in3 => \N__42500\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_17_14_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            clk => \N__47942\,
            ce => \N__42591\,
            sr => \N__47302\
        );

    \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42723\,
            in1 => \N__44431\,
            in2 => \_gnd_net_\,
            in3 => \N__42497\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            clk => \N__47942\,
            ce => \N__42591\,
            sr => \N__47302\
        );

    \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42708\,
            in1 => \N__44400\,
            in2 => \_gnd_net_\,
            in3 => \N__42494\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            clk => \N__47942\,
            ce => \N__42591\,
            sr => \N__47302\
        );

    \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42720\,
            in1 => \N__44835\,
            in2 => \_gnd_net_\,
            in3 => \N__42491\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            clk => \N__47942\,
            ce => \N__42591\,
            sr => \N__47302\
        );

    \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42709\,
            in1 => \N__44808\,
            in2 => \_gnd_net_\,
            in3 => \N__42488\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            clk => \N__47942\,
            ce => \N__42591\,
            sr => \N__47302\
        );

    \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42721\,
            in1 => \N__44781\,
            in2 => \_gnd_net_\,
            in3 => \N__42485\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            clk => \N__47942\,
            ce => \N__42591\,
            sr => \N__47302\
        );

    \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42710\,
            in1 => \N__44760\,
            in2 => \_gnd_net_\,
            in3 => \N__42482\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            clk => \N__47942\,
            ce => \N__42591\,
            sr => \N__47302\
        );

    \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42722\,
            in1 => \N__44739\,
            in2 => \_gnd_net_\,
            in3 => \N__42533\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            clk => \N__47942\,
            ce => \N__42591\,
            sr => \N__47302\
        );

    \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42712\,
            in1 => \N__44715\,
            in2 => \_gnd_net_\,
            in3 => \N__42530\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_17_15_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            clk => \N__47931\,
            ce => \N__42599\,
            sr => \N__47308\
        );

    \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42737\,
            in1 => \N__44688\,
            in2 => \_gnd_net_\,
            in3 => \N__42527\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            clk => \N__47931\,
            ce => \N__42599\,
            sr => \N__47308\
        );

    \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42713\,
            in1 => \N__44652\,
            in2 => \_gnd_net_\,
            in3 => \N__42524\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            clk => \N__47931\,
            ce => \N__42599\,
            sr => \N__47308\
        );

    \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42738\,
            in1 => \N__45132\,
            in2 => \_gnd_net_\,
            in3 => \N__42521\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            clk => \N__47931\,
            ce => \N__42599\,
            sr => \N__47308\
        );

    \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42714\,
            in1 => \N__45100\,
            in2 => \_gnd_net_\,
            in3 => \N__42518\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            clk => \N__47931\,
            ce => \N__42599\,
            sr => \N__47308\
        );

    \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42739\,
            in1 => \N__45066\,
            in2 => \_gnd_net_\,
            in3 => \N__42515\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            clk => \N__47931\,
            ce => \N__42599\,
            sr => \N__47308\
        );

    \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42715\,
            in1 => \N__45027\,
            in2 => \_gnd_net_\,
            in3 => \N__42512\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            clk => \N__47931\,
            ce => \N__42599\,
            sr => \N__47308\
        );

    \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42740\,
            in1 => \N__45000\,
            in2 => \_gnd_net_\,
            in3 => \N__42509\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            clk => \N__47931\,
            ce => \N__42599\,
            sr => \N__47308\
        );

    \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42702\,
            in1 => \N__44967\,
            in2 => \_gnd_net_\,
            in3 => \N__42755\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_17_16_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            clk => \N__47923\,
            ce => \N__42595\,
            sr => \N__47314\
        );

    \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42706\,
            in1 => \N__44931\,
            in2 => \_gnd_net_\,
            in3 => \N__42752\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            clk => \N__47923\,
            ce => \N__42595\,
            sr => \N__47314\
        );

    \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42703\,
            in1 => \N__44871\,
            in2 => \_gnd_net_\,
            in3 => \N__42749\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            clk => \N__47923\,
            ce => \N__42595\,
            sr => \N__47314\
        );

    \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42707\,
            in1 => \N__45435\,
            in2 => \_gnd_net_\,
            in3 => \N__42746\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            clk => \N__47923\,
            ce => \N__42595\,
            sr => \N__47314\
        );

    \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42704\,
            in1 => \N__44893\,
            in2 => \_gnd_net_\,
            in3 => \N__42743\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_28\,
            clk => \N__47923\,
            ce => \N__42595\,
            sr => \N__47314\
        );

    \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__45415\,
            in1 => \N__42705\,
            in2 => \_gnd_net_\,
            in3 => \N__42602\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47923\,
            ce => \N__42595\,
            sr => \N__47314\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6O9B2_14_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101010101"
        )
    port map (
            in0 => \N__46348\,
            in1 => \N__46028\,
            in2 => \_gnd_net_\,
            in3 => \N__45925\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_293\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__44948\,
            in1 => \N__44984\,
            in2 => \N__44909\,
            in3 => \N__45011\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__45086\,
            in1 => \N__45116\,
            in2 => \N__45050\,
            in3 => \N__44636\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__44669\,
            in1 => \N__42956\,
            in2 => \N__42950\,
            in3 => \N__42938\,
            lcout => \delay_measurement_inst.N_358\,
            ltout => \delay_measurement_inst.N_358_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2EEG9_15_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000100"
        )
    port map (
            in0 => \N__46277\,
            in1 => \N__42947\,
            in2 => \N__42941\,
            in3 => \N__46213\,
            lcout => \delay_measurement_inst.N_324\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO4MS_29_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45401\,
            in2 => \_gnd_net_\,
            in3 => \N__44855\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__43061\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43022\,
            lcout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSR_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__43062\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43023\,
            lcout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_esr_RNO_0_9_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__46029\,
            in1 => \N__45926\,
            in2 => \N__46276\,
            in3 => \N__48080\,
            lcout => \delay_measurement_inst.N_307\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.start_timer_hc_RNO_1_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42823\,
            in2 => \_gnd_net_\,
            in3 => \N__42862\,
            lcout => OPEN,
            ltout => \phase_controller_slave.start_timer_hc_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.start_timer_hc_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011110010"
        )
    port map (
            in0 => \N__43664\,
            in1 => \N__42923\,
            in2 => \N__42911\,
            in3 => \N__42903\,
            lcout => \phase_controller_slave.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47906\,
            ce => 'H',
            sr => \N__47338\
        );

    \phase_controller_slave.state_2_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__42863\,
            in1 => \N__42774\,
            in2 => \N__42827\,
            in3 => \N__42980\,
            lcout => \phase_controller_slave.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47906\,
            ce => 'H',
            sr => \N__47338\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_11_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__43568\,
            in1 => \N__43665\,
            in2 => \N__43856\,
            in3 => \N__45500\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47906\,
            ce => 'H',
            sr => \N__47338\
        );

    \phase_controller_slave.stoper_hc.time_passed_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__42981\,
            in1 => \N__43064\,
            in2 => \N__43043\,
            in3 => \N__43034\,
            lcout => \phase_controller_slave.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47906\,
            ce => 'H',
            sr => \N__47338\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_12_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__43569\,
            in1 => \N__43842\,
            in2 => \N__43710\,
            in3 => \N__45473\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47901\,
            ce => 'H',
            sr => \N__47349\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_9_LC_17_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010100010"
        )
    port map (
            in0 => \N__45563\,
            in1 => \N__43573\,
            in2 => \N__43855\,
            in3 => \N__43681\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47901\,
            ce => 'H',
            sr => \N__47349\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_15_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__43571\,
            in1 => \N__43844\,
            in2 => \N__43712\,
            in3 => \N__45845\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47901\,
            ce => 'H',
            sr => \N__47349\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_16_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__43839\,
            in1 => \N__43666\,
            in2 => \N__43587\,
            in3 => \N__45818\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47901\,
            ce => 'H',
            sr => \N__47349\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_13_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__43570\,
            in1 => \N__43843\,
            in2 => \N__43711\,
            in3 => \N__45446\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47901\,
            ce => 'H',
            sr => \N__47349\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_17_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__43840\,
            in1 => \N__43667\,
            in2 => \N__43588\,
            in3 => \N__45791\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47901\,
            ce => 'H',
            sr => \N__47349\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_18_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__43572\,
            in1 => \N__43845\,
            in2 => \N__43713\,
            in3 => \N__45764\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47901\,
            ce => 'H',
            sr => \N__47349\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_19_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__43841\,
            in1 => \N__43668\,
            in2 => \N__43589\,
            in3 => \N__45734\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47901\,
            ce => 'H',
            sr => \N__47349\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4_3_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__46312\,
            in1 => \N__46941\,
            in2 => \N__46177\,
            in3 => \N__46563\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__48299\,
            in1 => \N__45724\,
            in2 => \N__43463\,
            in3 => \N__43456\,
            lcout => \phase_controller_inst1.stoper_tr.N_279\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_6_LC_17_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010111011"
        )
    port map (
            in0 => \N__45693\,
            in1 => \N__46155\,
            in2 => \N__43460\,
            in3 => \N__46313\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.target_time_14_LC_17_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__45695\,
            in1 => \N__46173\,
            in2 => \_gnd_net_\,
            in3 => \N__46317\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47888\,
            ce => \N__43358\,
            sr => \N__47366\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_9_LC_17_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__45694\,
            in1 => \N__46179\,
            in2 => \_gnd_net_\,
            in3 => \N__46319\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a3_1_LC_17_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__46884\,
            in1 => \N__46422\,
            in2 => \_gnd_net_\,
            in3 => \N__43264\,
            lcout => \phase_controller_inst1.stoper_tr.N_262\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0_6_LC_17_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__45728\,
            in1 => \N__43222\,
            in2 => \_gnd_net_\,
            in3 => \N__46178\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_15_LC_17_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45708\,
            in2 => \_gnd_net_\,
            in3 => \N__46180\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47874\,
            ce => \N__43124\,
            sr => \N__47387\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44381\,
            lcout => \delay_measurement_inst.elapsed_time_hc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47986\,
            ce => \N__44332\,
            sr => \N__47277\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__44298\,
            in1 => \N__44277\,
            in2 => \N__44250\,
            in3 => \N__44220\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITS8G_14_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44181\,
            in2 => \_gnd_net_\,
            in3 => \N__44133\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_a0_1\,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_a0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA5CC2_6_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__44067\,
            in1 => \N__44013\,
            in2 => \N__43970\,
            in3 => \N__43928\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto31_a0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43900\,
            lcout => \delay_measurement_inst.elapsed_time_tr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47952\,
            ce => \N__45373\,
            sr => \N__47296\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_18_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43879\,
            lcout => \delay_measurement_inst.elapsed_time_tr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47952\,
            ce => \N__45373\,
            sr => \N__47296\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43901\,
            in2 => \N__44626\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.elapsed_time_tr_3\,
            ltout => OPEN,
            carryin => \bfn_18_15_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__47943\,
            ce => \N__45389\,
            sr => \N__47303\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43880\,
            in2 => \N__44599\,
            in3 => \N__43859\,
            lcout => \delay_measurement_inst.elapsed_time_tr_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__47943\,
            ce => \N__45389\,
            sr => \N__47303\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44572\,
            in2 => \N__44627\,
            in3 => \N__44603\,
            lcout => \delay_measurement_inst.elapsed_time_tr_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__47943\,
            ce => \N__45389\,
            sr => \N__47303\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44548\,
            in2 => \N__44600\,
            in3 => \N__44576\,
            lcout => \delay_measurement_inst.delay_tr_reg3lto6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__47943\,
            ce => \N__45389\,
            sr => \N__47303\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44573\,
            in2 => \N__44525\,
            in3 => \N__44552\,
            lcout => \delay_measurement_inst.elapsed_time_tr_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__47943\,
            ce => \N__45389\,
            sr => \N__47303\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44549\,
            in2 => \N__44494\,
            in3 => \N__44528\,
            lcout => \delay_measurement_inst.elapsed_time_tr_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__47943\,
            ce => \N__45389\,
            sr => \N__47303\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44524\,
            in2 => \N__44461\,
            in3 => \N__44498\,
            lcout => \delay_measurement_inst.delay_tr_reg3lto9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__47943\,
            ce => \N__45389\,
            sr => \N__47303\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_18_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44430\,
            in2 => \N__44495\,
            in3 => \N__44468\,
            lcout => \delay_measurement_inst.elapsed_time_tr_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__47943\,
            ce => \N__45389\,
            sr => \N__47303\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44465\,
            in2 => \N__44411\,
            in3 => \N__44438\,
            lcout => \delay_measurement_inst.elapsed_time_tr_11\,
            ltout => OPEN,
            carryin => \bfn_18_16_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__47932\,
            ce => \N__45377\,
            sr => \N__47309\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44435\,
            in2 => \N__44846\,
            in3 => \N__44414\,
            lcout => \delay_measurement_inst.elapsed_time_tr_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__47932\,
            ce => \N__45377\,
            sr => \N__47309\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44410\,
            in2 => \N__44815\,
            in3 => \N__44384\,
            lcout => \delay_measurement_inst.elapsed_time_tr_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__47932\,
            ce => \N__45377\,
            sr => \N__47309\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44845\,
            in2 => \N__44788\,
            in3 => \N__44819\,
            lcout => \delay_measurement_inst.delay_tr_reg3lto14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__47932\,
            ce => \N__45377\,
            sr => \N__47309\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44761\,
            in2 => \N__44816\,
            in3 => \N__44792\,
            lcout => \delay_measurement_inst.delay_tr_reg3lto15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__47932\,
            ce => \N__45377\,
            sr => \N__47309\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44740\,
            in2 => \N__44789\,
            in3 => \N__44765\,
            lcout => \delay_measurement_inst.elapsed_time_tr_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__47932\,
            ce => \N__45377\,
            sr => \N__47309\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44762\,
            in2 => \N__44720\,
            in3 => \N__44744\,
            lcout => \delay_measurement_inst.elapsed_time_tr_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__47932\,
            ce => \N__45377\,
            sr => \N__47309\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_18_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44741\,
            in2 => \N__44692\,
            in3 => \N__44723\,
            lcout => \delay_measurement_inst.elapsed_time_tr_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__47932\,
            ce => \N__45377\,
            sr => \N__47309\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44719\,
            in2 => \N__44659\,
            in3 => \N__44696\,
            lcout => \delay_measurement_inst.elapsed_time_tr_19\,
            ltout => OPEN,
            carryin => \bfn_18_17_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__47924\,
            ce => \N__45387\,
            sr => \N__47315\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44693\,
            in2 => \N__45139\,
            in3 => \N__44663\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__47924\,
            ce => \N__45387\,
            sr => \N__47315\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45106\,
            in2 => \N__44660\,
            in3 => \N__44630\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__47924\,
            ce => \N__45387\,
            sr => \N__47315\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45073\,
            in2 => \N__45140\,
            in3 => \N__45110\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__47924\,
            ce => \N__45387\,
            sr => \N__47315\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45107\,
            in2 => \N__45038\,
            in3 => \N__45080\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__47924\,
            ce => \N__45387\,
            sr => \N__47315\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45001\,
            in2 => \N__45077\,
            in3 => \N__45041\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__47924\,
            ce => \N__45387\,
            sr => \N__47315\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45037\,
            in2 => \N__44971\,
            in3 => \N__45005\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__47924\,
            ce => \N__45387\,
            sr => \N__47315\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_18_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45002\,
            in2 => \N__44932\,
            in3 => \N__44978\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__47924\,
            ce => \N__45387\,
            sr => \N__47315\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_18_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44975\,
            in2 => \N__44878\,
            in3 => \N__44942\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\,
            ltout => OPEN,
            carryin => \bfn_18_18_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__47917\,
            ce => \N__45388\,
            sr => \N__47321\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45436\,
            in2 => \N__44939\,
            in3 => \N__44897\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__47917\,
            ce => \N__45388\,
            sr => \N__47321\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44894\,
            in2 => \N__44879\,
            in3 => \N__44849\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__47917\,
            ce => \N__45388\,
            sr => \N__47321\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_18_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45437\,
            in2 => \N__45419\,
            in3 => \N__45395\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__47917\,
            ce => \N__45388\,
            sr => \N__47321\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45392\,
            lcout => \delay_measurement_inst.elapsed_time_tr_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47917\,
            ce => \N__45388\,
            sr => \N__47321\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_18_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45338\,
            in2 => \N__45332\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_19_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45302\,
            in2 => \_gnd_net_\,
            in3 => \N__45272\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_18_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45269\,
            in2 => \N__45263\,
            in3 => \N__45230\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45227\,
            in2 => \_gnd_net_\,
            in3 => \N__45197\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_18_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45194\,
            in2 => \_gnd_net_\,
            in3 => \N__45161\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_18_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45158\,
            in2 => \_gnd_net_\,
            in3 => \N__45653\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45650\,
            in2 => \_gnd_net_\,
            in3 => \N__45620\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_18_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45617\,
            in2 => \_gnd_net_\,
            in3 => \N__45584\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45577\,
            in2 => \_gnd_net_\,
            in3 => \N__45557\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9\,
            ltout => OPEN,
            carryin => \bfn_18_20_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45554\,
            in2 => \_gnd_net_\,
            in3 => \N__45521\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45514\,
            in2 => \_gnd_net_\,
            in3 => \N__45494\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_18_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45487\,
            in2 => \_gnd_net_\,
            in3 => \N__45467\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_18_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45460\,
            in2 => \_gnd_net_\,
            in3 => \N__45440\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_18_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45896\,
            in2 => \_gnd_net_\,
            in3 => \N__45866\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_18_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45859\,
            in2 => \_gnd_net_\,
            in3 => \N__45839\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_18_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45832\,
            in2 => \_gnd_net_\,
            in3 => \N__45812\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_18_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45805\,
            in2 => \_gnd_net_\,
            in3 => \N__45785\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17\,
            ltout => OPEN,
            carryin => \bfn_18_21_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_18_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45778\,
            in2 => \_gnd_net_\,
            in3 => \N__45758\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_18_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45751\,
            in2 => \_gnd_net_\,
            in3 => \N__45737\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1_6_LC_18_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__46815\,
            in1 => \N__46758\,
            in2 => \_gnd_net_\,
            in3 => \N__46614\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_i_o2_15_LC_18_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__48402\,
            in1 => \N__48366\,
            in2 => \N__48055\,
            in3 => \N__48327\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6FAF_1_LC_20_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__46090\,
            in1 => \N__46021\,
            in2 => \N__46468\,
            in3 => \N__46637\,
            lcout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI86841_2_LC_20_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000101"
        )
    port map (
            in0 => \N__48543\,
            in1 => \N__46914\,
            in2 => \N__46734\,
            in3 => \N__46467\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIOKG82_18_LC_20_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__48154\,
            in1 => \N__48438\,
            in2 => \N__46037\,
            in3 => \N__45983\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI61PC3_6_LC_20_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__46030\,
            in1 => \N__46375\,
            in2 => \N__45986\,
            in3 => \N__46647\,
            lcout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_20_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46969\,
            in2 => \_gnd_net_\,
            in3 => \N__46591\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_320_4\,
            ltout => \delay_measurement_inst.delay_tr_timer.N_320_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRN391_3_LC_20_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__46341\,
            in1 => \N__46915\,
            in2 => \N__45977\,
            in3 => \N__45974\,
            lcout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILUIS_14_LC_20_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__46340\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46254\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILUISZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_20_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__45964\,
            in1 => \N__48520\,
            in2 => \N__46699\,
            in3 => \N__45949\,
            lcout => \delay_measurement_inst.N_328\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_20_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__48442\,
            in1 => \N__46735\,
            in2 => \N__48147\,
            in3 => \N__48550\,
            lcout => \delay_measurement_inst.elapsed_time_ns_1_RNIM96P1_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6_7_LC_20_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__46786\,
            in1 => \N__45912\,
            in2 => \N__46850\,
            in3 => \N__48090\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_331\,
            ltout => \delay_measurement_inst.delay_tr_timer.N_331_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC3FA_15_LC_20_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__46272\,
            in1 => \N__46204\,
            in2 => \N__46394\,
            in3 => \N__46391\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.N_321_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_20_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000101"
        )
    port map (
            in0 => \N__48252\,
            in1 => \N__46385\,
            in2 => \N__46379\,
            in3 => \N__46363\,
            lcout => \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_esr_RNO_0_14_LC_20_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__46273\,
            in1 => \N__48253\,
            in2 => \_gnd_net_\,
            in3 => \N__46206\,
            lcout => \delay_measurement_inst.delay_tr_reg_esr_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_20_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__48091\,
            in1 => \N__46376\,
            in2 => \_gnd_net_\,
            in3 => \N__46205\,
            lcout => \delay_measurement_inst.N_301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI80KG7_6_LC_20_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__46274\,
            in1 => \N__46648\,
            in2 => \_gnd_net_\,
            in3 => \N__46364\,
            lcout => \delay_measurement_inst.elapsed_time_ns_1_RNI80KG7_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_esr_14_LC_20_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__48121\,
            in1 => \N__46355\,
            in2 => \N__48257\,
            in3 => \N__46349\,
            lcout => measured_delay_tr_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47933\,
            ce => \N__47490\,
            sr => \N__47322\
        );

    \delay_measurement_inst.delay_tr_reg_esr_15_LC_20_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010101000"
        )
    port map (
            in0 => \N__46275\,
            in1 => \N__48215\,
            in2 => \N__46217\,
            in3 => \N__48122\,
            lcout => measured_delay_tr_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47933\,
            ce => \N__47490\,
            sr => \N__47322\
        );

    \delay_measurement_inst.delay_tr_reg_ess_1_LC_20_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__46488\,
            in1 => \N__46536\,
            in2 => \N__48258\,
            in3 => \N__46091\,
            lcout => measured_delay_tr_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47933\,
            ce => \N__47490\,
            sr => \N__47322\
        );

    \delay_measurement_inst.delay_tr_reg_esr_5_LC_20_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__46534\,
            in1 => \N__46487\,
            in2 => \N__46973\,
            in3 => \N__48216\,
            lcout => measured_delay_tr_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47933\,
            ce => \N__47490\,
            sr => \N__47322\
        );

    \delay_measurement_inst.delay_tr_reg_ess_3_LC_20_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__46489\,
            in1 => \N__46537\,
            in2 => \N__48259\,
            in3 => \N__46916\,
            lcout => measured_delay_tr_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47933\,
            ce => \N__47490\,
            sr => \N__47322\
        );

    \delay_measurement_inst.delay_tr_reg_esr_8_LC_20_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__46535\,
            in1 => \N__48211\,
            in2 => \_gnd_net_\,
            in3 => \N__46849\,
            lcout => measured_delay_tr_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47933\,
            ce => \N__47490\,
            sr => \N__47322\
        );

    \delay_measurement_inst.delay_tr_reg_esr_7_LC_20_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__46541\,
            in1 => \N__48274\,
            in2 => \_gnd_net_\,
            in3 => \N__46787\,
            lcout => measured_delay_tr_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47925\,
            ce => \N__47492\,
            sr => \N__47327\
        );

    \delay_measurement_inst.delay_tr_reg_esr_17_LC_20_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__48273\,
            in1 => \N__46736\,
            in2 => \_gnd_net_\,
            in3 => \N__48107\,
            lcout => measured_delay_tr_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47925\,
            ce => \N__47492\,
            sr => \N__47327\
        );

    \delay_measurement_inst.delay_tr_reg_esr_13_LC_20_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__46700\,
            in1 => \N__48265\,
            in2 => \_gnd_net_\,
            in3 => \N__48494\,
            lcout => measured_delay_tr_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47925\,
            ce => \N__47492\,
            sr => \N__47327\
        );

    \delay_measurement_inst.delay_tr_reg_esr_6_LC_20_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000001"
        )
    port map (
            in0 => \N__46540\,
            in1 => \N__46499\,
            in2 => \N__48283\,
            in3 => \N__46649\,
            lcout => measured_delay_tr_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47925\,
            ce => \N__47492\,
            sr => \N__47327\
        );

    \delay_measurement_inst.delay_tr_reg_esr_4_LC_20_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__46498\,
            in1 => \N__46539\,
            in2 => \N__48284\,
            in3 => \N__46592\,
            lcout => measured_delay_tr_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47925\,
            ce => \N__47492\,
            sr => \N__47327\
        );

    \delay_measurement_inst.delay_tr_reg_esr_2_LC_20_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__46538\,
            in1 => \N__46497\,
            in2 => \N__48282\,
            in3 => \N__46472\,
            lcout => measured_delay_tr_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47925\,
            ce => \N__47492\,
            sr => \N__47327\
        );

    \delay_measurement_inst.delay_tr_reg_esr_16_LC_20_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__48551\,
            in1 => \N__48266\,
            in2 => \_gnd_net_\,
            in3 => \N__48106\,
            lcout => measured_delay_tr_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47925\,
            ce => \N__47492\,
            sr => \N__47327\
        );

    \delay_measurement_inst.delay_tr_reg_esr_11_LC_20_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000100010"
        )
    port map (
            in0 => \N__48524\,
            in1 => \N__48495\,
            in2 => \_gnd_net_\,
            in3 => \N__48278\,
            lcout => measured_delay_tr_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47918\,
            ce => \N__47511\,
            sr => \N__47339\
        );

    \delay_measurement_inst.delay_tr_reg_esr_18_LC_20_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__48279\,
            in1 => \N__48443\,
            in2 => \_gnd_net_\,
            in3 => \N__48119\,
            lcout => measured_delay_tr_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47918\,
            ce => \N__47511\,
            sr => \N__47339\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_3_LC_20_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__48388\,
            in1 => \N__48357\,
            in2 => \N__48044\,
            in3 => \N__48318\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_31_LC_21_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47459\,
            in2 => \_gnd_net_\,
            in3 => \N__48290\,
            lcout => \delay_measurement_inst.un3_elapsed_time_tr_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_esr_19_LC_21_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__48280\,
            in1 => \N__48155\,
            in2 => \_gnd_net_\,
            in3 => \N__48120\,
            lcout => measured_delay_tr_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47934\,
            ce => \N__47491\,
            sr => \N__47340\
        );
end \INTERFACE\;
