// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Oct 8 2025 23:18:14

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "MAIN" view "INTERFACE"

module MAIN (
    s3_phy,
    il_min_comp2,
    il_max_comp1,
    s1_phy,
    reset,
    il_min_comp1,
    delay_tr_input,
    s4_phy,
    rgb_g,
    start_stop,
    s2_phy,
    rgb_r,
    rgb_b,
    pwm_output,
    il_max_comp2,
    delay_hc_input);

    output s3_phy;
    input il_min_comp2;
    input il_max_comp1;
    output s1_phy;
    input reset;
    input il_min_comp1;
    input delay_tr_input;
    output s4_phy;
    output rgb_g;
    input start_stop;
    output s2_phy;
    output rgb_r;
    output rgb_b;
    output pwm_output;
    input il_max_comp2;
    input delay_hc_input;

    wire N__48353;
    wire N__48352;
    wire N__48351;
    wire N__48342;
    wire N__48341;
    wire N__48340;
    wire N__48333;
    wire N__48332;
    wire N__48331;
    wire N__48324;
    wire N__48323;
    wire N__48322;
    wire N__48315;
    wire N__48314;
    wire N__48313;
    wire N__48306;
    wire N__48305;
    wire N__48304;
    wire N__48297;
    wire N__48296;
    wire N__48295;
    wire N__48288;
    wire N__48287;
    wire N__48286;
    wire N__48279;
    wire N__48278;
    wire N__48277;
    wire N__48270;
    wire N__48269;
    wire N__48268;
    wire N__48261;
    wire N__48260;
    wire N__48259;
    wire N__48252;
    wire N__48251;
    wire N__48250;
    wire N__48243;
    wire N__48242;
    wire N__48241;
    wire N__48224;
    wire N__48221;
    wire N__48218;
    wire N__48215;
    wire N__48214;
    wire N__48211;
    wire N__48208;
    wire N__48205;
    wire N__48202;
    wire N__48197;
    wire N__48196;
    wire N__48195;
    wire N__48192;
    wire N__48189;
    wire N__48186;
    wire N__48185;
    wire N__48184;
    wire N__48183;
    wire N__48182;
    wire N__48181;
    wire N__48180;
    wire N__48179;
    wire N__48178;
    wire N__48177;
    wire N__48176;
    wire N__48175;
    wire N__48174;
    wire N__48173;
    wire N__48164;
    wire N__48159;
    wire N__48158;
    wire N__48157;
    wire N__48156;
    wire N__48155;
    wire N__48154;
    wire N__48153;
    wire N__48150;
    wire N__48149;
    wire N__48146;
    wire N__48145;
    wire N__48142;
    wire N__48139;
    wire N__48126;
    wire N__48121;
    wire N__48118;
    wire N__48115;
    wire N__48110;
    wire N__48093;
    wire N__48088;
    wire N__48085;
    wire N__48074;
    wire N__48073;
    wire N__48072;
    wire N__48071;
    wire N__48068;
    wire N__48067;
    wire N__48066;
    wire N__48065;
    wire N__48064;
    wire N__48063;
    wire N__48062;
    wire N__48061;
    wire N__48060;
    wire N__48059;
    wire N__48056;
    wire N__48053;
    wire N__48050;
    wire N__48049;
    wire N__48048;
    wire N__48047;
    wire N__48042;
    wire N__48039;
    wire N__48036;
    wire N__48033;
    wire N__48030;
    wire N__48029;
    wire N__48028;
    wire N__48027;
    wire N__48026;
    wire N__48025;
    wire N__48024;
    wire N__48015;
    wire N__48002;
    wire N__47999;
    wire N__47998;
    wire N__47997;
    wire N__47988;
    wire N__47983;
    wire N__47974;
    wire N__47969;
    wire N__47966;
    wire N__47961;
    wire N__47948;
    wire N__47947;
    wire N__47946;
    wire N__47943;
    wire N__47942;
    wire N__47941;
    wire N__47940;
    wire N__47937;
    wire N__47934;
    wire N__47933;
    wire N__47930;
    wire N__47923;
    wire N__47916;
    wire N__47915;
    wire N__47914;
    wire N__47913;
    wire N__47912;
    wire N__47911;
    wire N__47910;
    wire N__47903;
    wire N__47898;
    wire N__47895;
    wire N__47894;
    wire N__47893;
    wire N__47892;
    wire N__47891;
    wire N__47890;
    wire N__47889;
    wire N__47888;
    wire N__47887;
    wire N__47886;
    wire N__47879;
    wire N__47874;
    wire N__47873;
    wire N__47872;
    wire N__47867;
    wire N__47850;
    wire N__47845;
    wire N__47840;
    wire N__47831;
    wire N__47828;
    wire N__47825;
    wire N__47824;
    wire N__47821;
    wire N__47818;
    wire N__47813;
    wire N__47810;
    wire N__47807;
    wire N__47806;
    wire N__47803;
    wire N__47800;
    wire N__47797;
    wire N__47794;
    wire N__47791;
    wire N__47788;
    wire N__47783;
    wire N__47782;
    wire N__47781;
    wire N__47780;
    wire N__47779;
    wire N__47776;
    wire N__47773;
    wire N__47770;
    wire N__47767;
    wire N__47764;
    wire N__47761;
    wire N__47756;
    wire N__47753;
    wire N__47750;
    wire N__47745;
    wire N__47742;
    wire N__47735;
    wire N__47732;
    wire N__47729;
    wire N__47726;
    wire N__47725;
    wire N__47724;
    wire N__47723;
    wire N__47720;
    wire N__47713;
    wire N__47708;
    wire N__47707;
    wire N__47706;
    wire N__47701;
    wire N__47698;
    wire N__47695;
    wire N__47694;
    wire N__47691;
    wire N__47688;
    wire N__47685;
    wire N__47684;
    wire N__47681;
    wire N__47678;
    wire N__47673;
    wire N__47666;
    wire N__47665;
    wire N__47664;
    wire N__47663;
    wire N__47660;
    wire N__47657;
    wire N__47652;
    wire N__47649;
    wire N__47642;
    wire N__47641;
    wire N__47638;
    wire N__47637;
    wire N__47634;
    wire N__47631;
    wire N__47628;
    wire N__47625;
    wire N__47622;
    wire N__47615;
    wire N__47612;
    wire N__47609;
    wire N__47606;
    wire N__47605;
    wire N__47604;
    wire N__47599;
    wire N__47598;
    wire N__47597;
    wire N__47596;
    wire N__47595;
    wire N__47594;
    wire N__47593;
    wire N__47590;
    wire N__47587;
    wire N__47578;
    wire N__47573;
    wire N__47570;
    wire N__47567;
    wire N__47564;
    wire N__47561;
    wire N__47558;
    wire N__47555;
    wire N__47552;
    wire N__47547;
    wire N__47540;
    wire N__47539;
    wire N__47538;
    wire N__47537;
    wire N__47536;
    wire N__47535;
    wire N__47534;
    wire N__47531;
    wire N__47530;
    wire N__47527;
    wire N__47524;
    wire N__47521;
    wire N__47520;
    wire N__47513;
    wire N__47510;
    wire N__47507;
    wire N__47502;
    wire N__47499;
    wire N__47496;
    wire N__47493;
    wire N__47488;
    wire N__47487;
    wire N__47484;
    wire N__47481;
    wire N__47478;
    wire N__47475;
    wire N__47472;
    wire N__47469;
    wire N__47466;
    wire N__47463;
    wire N__47456;
    wire N__47447;
    wire N__47444;
    wire N__47443;
    wire N__47442;
    wire N__47439;
    wire N__47436;
    wire N__47435;
    wire N__47432;
    wire N__47429;
    wire N__47426;
    wire N__47421;
    wire N__47418;
    wire N__47413;
    wire N__47410;
    wire N__47407;
    wire N__47402;
    wire N__47401;
    wire N__47400;
    wire N__47397;
    wire N__47392;
    wire N__47391;
    wire N__47390;
    wire N__47387;
    wire N__47384;
    wire N__47379;
    wire N__47376;
    wire N__47371;
    wire N__47366;
    wire N__47363;
    wire N__47360;
    wire N__47357;
    wire N__47354;
    wire N__47351;
    wire N__47350;
    wire N__47349;
    wire N__47348;
    wire N__47347;
    wire N__47346;
    wire N__47345;
    wire N__47344;
    wire N__47343;
    wire N__47342;
    wire N__47341;
    wire N__47340;
    wire N__47339;
    wire N__47338;
    wire N__47337;
    wire N__47336;
    wire N__47335;
    wire N__47334;
    wire N__47333;
    wire N__47332;
    wire N__47331;
    wire N__47330;
    wire N__47329;
    wire N__47328;
    wire N__47327;
    wire N__47326;
    wire N__47325;
    wire N__47324;
    wire N__47323;
    wire N__47322;
    wire N__47321;
    wire N__47320;
    wire N__47319;
    wire N__47318;
    wire N__47317;
    wire N__47316;
    wire N__47315;
    wire N__47314;
    wire N__47313;
    wire N__47312;
    wire N__47311;
    wire N__47310;
    wire N__47309;
    wire N__47308;
    wire N__47307;
    wire N__47306;
    wire N__47305;
    wire N__47304;
    wire N__47303;
    wire N__47302;
    wire N__47301;
    wire N__47300;
    wire N__47299;
    wire N__47298;
    wire N__47297;
    wire N__47296;
    wire N__47295;
    wire N__47294;
    wire N__47293;
    wire N__47292;
    wire N__47291;
    wire N__47290;
    wire N__47289;
    wire N__47288;
    wire N__47287;
    wire N__47286;
    wire N__47285;
    wire N__47284;
    wire N__47283;
    wire N__47282;
    wire N__47281;
    wire N__47280;
    wire N__47279;
    wire N__47278;
    wire N__47277;
    wire N__47276;
    wire N__47275;
    wire N__47274;
    wire N__47273;
    wire N__47272;
    wire N__47271;
    wire N__47270;
    wire N__47269;
    wire N__47268;
    wire N__47267;
    wire N__47266;
    wire N__47265;
    wire N__47264;
    wire N__47263;
    wire N__47262;
    wire N__47261;
    wire N__47260;
    wire N__47259;
    wire N__47258;
    wire N__47257;
    wire N__47256;
    wire N__47255;
    wire N__47254;
    wire N__47253;
    wire N__47252;
    wire N__47251;
    wire N__47250;
    wire N__47249;
    wire N__47248;
    wire N__47247;
    wire N__47246;
    wire N__47245;
    wire N__47244;
    wire N__47243;
    wire N__47242;
    wire N__47241;
    wire N__47240;
    wire N__47239;
    wire N__47238;
    wire N__47237;
    wire N__47236;
    wire N__47235;
    wire N__47234;
    wire N__47233;
    wire N__47232;
    wire N__47231;
    wire N__47230;
    wire N__47229;
    wire N__47228;
    wire N__47227;
    wire N__47226;
    wire N__47225;
    wire N__47224;
    wire N__47223;
    wire N__47222;
    wire N__47221;
    wire N__47220;
    wire N__47219;
    wire N__47218;
    wire N__47217;
    wire N__47216;
    wire N__47215;
    wire N__47214;
    wire N__47213;
    wire N__47212;
    wire N__47211;
    wire N__47210;
    wire N__47209;
    wire N__47208;
    wire N__47207;
    wire N__47206;
    wire N__47205;
    wire N__47204;
    wire N__47203;
    wire N__47202;
    wire N__47201;
    wire N__47200;
    wire N__47199;
    wire N__47198;
    wire N__47197;
    wire N__47196;
    wire N__47195;
    wire N__47194;
    wire N__47193;
    wire N__47192;
    wire N__47191;
    wire N__47190;
    wire N__47189;
    wire N__46862;
    wire N__46859;
    wire N__46858;
    wire N__46857;
    wire N__46856;
    wire N__46853;
    wire N__46852;
    wire N__46849;
    wire N__46846;
    wire N__46843;
    wire N__46840;
    wire N__46837;
    wire N__46834;
    wire N__46831;
    wire N__46828;
    wire N__46827;
    wire N__46826;
    wire N__46823;
    wire N__46820;
    wire N__46817;
    wire N__46812;
    wire N__46809;
    wire N__46806;
    wire N__46801;
    wire N__46796;
    wire N__46793;
    wire N__46790;
    wire N__46781;
    wire N__46780;
    wire N__46779;
    wire N__46778;
    wire N__46777;
    wire N__46774;
    wire N__46773;
    wire N__46770;
    wire N__46767;
    wire N__46764;
    wire N__46761;
    wire N__46758;
    wire N__46755;
    wire N__46752;
    wire N__46749;
    wire N__46746;
    wire N__46745;
    wire N__46744;
    wire N__46743;
    wire N__46742;
    wire N__46741;
    wire N__46740;
    wire N__46739;
    wire N__46738;
    wire N__46737;
    wire N__46736;
    wire N__46735;
    wire N__46734;
    wire N__46733;
    wire N__46732;
    wire N__46731;
    wire N__46730;
    wire N__46729;
    wire N__46728;
    wire N__46727;
    wire N__46726;
    wire N__46725;
    wire N__46724;
    wire N__46723;
    wire N__46722;
    wire N__46721;
    wire N__46720;
    wire N__46719;
    wire N__46718;
    wire N__46717;
    wire N__46716;
    wire N__46715;
    wire N__46714;
    wire N__46713;
    wire N__46712;
    wire N__46711;
    wire N__46710;
    wire N__46709;
    wire N__46708;
    wire N__46707;
    wire N__46706;
    wire N__46705;
    wire N__46704;
    wire N__46703;
    wire N__46702;
    wire N__46701;
    wire N__46698;
    wire N__46697;
    wire N__46696;
    wire N__46695;
    wire N__46694;
    wire N__46693;
    wire N__46692;
    wire N__46691;
    wire N__46690;
    wire N__46689;
    wire N__46688;
    wire N__46687;
    wire N__46686;
    wire N__46685;
    wire N__46684;
    wire N__46683;
    wire N__46682;
    wire N__46681;
    wire N__46680;
    wire N__46679;
    wire N__46678;
    wire N__46677;
    wire N__46676;
    wire N__46675;
    wire N__46674;
    wire N__46673;
    wire N__46672;
    wire N__46671;
    wire N__46670;
    wire N__46669;
    wire N__46668;
    wire N__46667;
    wire N__46666;
    wire N__46665;
    wire N__46664;
    wire N__46663;
    wire N__46662;
    wire N__46661;
    wire N__46660;
    wire N__46659;
    wire N__46658;
    wire N__46657;
    wire N__46656;
    wire N__46655;
    wire N__46654;
    wire N__46653;
    wire N__46652;
    wire N__46651;
    wire N__46650;
    wire N__46649;
    wire N__46648;
    wire N__46647;
    wire N__46646;
    wire N__46645;
    wire N__46644;
    wire N__46643;
    wire N__46642;
    wire N__46641;
    wire N__46640;
    wire N__46639;
    wire N__46638;
    wire N__46637;
    wire N__46636;
    wire N__46635;
    wire N__46634;
    wire N__46633;
    wire N__46632;
    wire N__46631;
    wire N__46630;
    wire N__46629;
    wire N__46628;
    wire N__46627;
    wire N__46624;
    wire N__46621;
    wire N__46620;
    wire N__46619;
    wire N__46618;
    wire N__46617;
    wire N__46616;
    wire N__46615;
    wire N__46614;
    wire N__46613;
    wire N__46612;
    wire N__46611;
    wire N__46610;
    wire N__46609;
    wire N__46608;
    wire N__46607;
    wire N__46606;
    wire N__46605;
    wire N__46604;
    wire N__46603;
    wire N__46602;
    wire N__46601;
    wire N__46600;
    wire N__46599;
    wire N__46598;
    wire N__46597;
    wire N__46596;
    wire N__46595;
    wire N__46298;
    wire N__46295;
    wire N__46292;
    wire N__46291;
    wire N__46288;
    wire N__46285;
    wire N__46280;
    wire N__46277;
    wire N__46274;
    wire N__46271;
    wire N__46270;
    wire N__46267;
    wire N__46264;
    wire N__46259;
    wire N__46256;
    wire N__46253;
    wire N__46250;
    wire N__46249;
    wire N__46246;
    wire N__46243;
    wire N__46238;
    wire N__46235;
    wire N__46232;
    wire N__46229;
    wire N__46226;
    wire N__46225;
    wire N__46222;
    wire N__46219;
    wire N__46214;
    wire N__46211;
    wire N__46208;
    wire N__46205;
    wire N__46202;
    wire N__46201;
    wire N__46198;
    wire N__46195;
    wire N__46192;
    wire N__46187;
    wire N__46184;
    wire N__46181;
    wire N__46178;
    wire N__46177;
    wire N__46174;
    wire N__46171;
    wire N__46166;
    wire N__46163;
    wire N__46160;
    wire N__46157;
    wire N__46156;
    wire N__46153;
    wire N__46150;
    wire N__46145;
    wire N__46142;
    wire N__46139;
    wire N__46136;
    wire N__46135;
    wire N__46132;
    wire N__46129;
    wire N__46124;
    wire N__46121;
    wire N__46118;
    wire N__46115;
    wire N__46112;
    wire N__46111;
    wire N__46108;
    wire N__46105;
    wire N__46100;
    wire N__46097;
    wire N__46094;
    wire N__46091;
    wire N__46090;
    wire N__46087;
    wire N__46084;
    wire N__46079;
    wire N__46076;
    wire N__46073;
    wire N__46070;
    wire N__46069;
    wire N__46066;
    wire N__46063;
    wire N__46058;
    wire N__46055;
    wire N__46052;
    wire N__46049;
    wire N__46048;
    wire N__46045;
    wire N__46042;
    wire N__46037;
    wire N__46034;
    wire N__46031;
    wire N__46028;
    wire N__46027;
    wire N__46024;
    wire N__46021;
    wire N__46016;
    wire N__46013;
    wire N__46010;
    wire N__46007;
    wire N__46004;
    wire N__46003;
    wire N__46000;
    wire N__45997;
    wire N__45992;
    wire N__45989;
    wire N__45986;
    wire N__45983;
    wire N__45982;
    wire N__45979;
    wire N__45976;
    wire N__45971;
    wire N__45968;
    wire N__45965;
    wire N__45962;
    wire N__45959;
    wire N__45958;
    wire N__45955;
    wire N__45954;
    wire N__45951;
    wire N__45948;
    wire N__45945;
    wire N__45942;
    wire N__45935;
    wire N__45932;
    wire N__45929;
    wire N__45926;
    wire N__45923;
    wire N__45920;
    wire N__45917;
    wire N__45914;
    wire N__45913;
    wire N__45910;
    wire N__45907;
    wire N__45904;
    wire N__45899;
    wire N__45898;
    wire N__45895;
    wire N__45892;
    wire N__45891;
    wire N__45886;
    wire N__45883;
    wire N__45880;
    wire N__45875;
    wire N__45872;
    wire N__45869;
    wire N__45866;
    wire N__45863;
    wire N__45860;
    wire N__45859;
    wire N__45856;
    wire N__45853;
    wire N__45850;
    wire N__45845;
    wire N__45844;
    wire N__45841;
    wire N__45838;
    wire N__45837;
    wire N__45832;
    wire N__45829;
    wire N__45826;
    wire N__45821;
    wire N__45818;
    wire N__45815;
    wire N__45812;
    wire N__45809;
    wire N__45806;
    wire N__45803;
    wire N__45802;
    wire N__45801;
    wire N__45798;
    wire N__45797;
    wire N__45796;
    wire N__45795;
    wire N__45794;
    wire N__45791;
    wire N__45790;
    wire N__45787;
    wire N__45786;
    wire N__45785;
    wire N__45782;
    wire N__45773;
    wire N__45770;
    wire N__45765;
    wire N__45762;
    wire N__45761;
    wire N__45760;
    wire N__45757;
    wire N__45748;
    wire N__45741;
    wire N__45736;
    wire N__45731;
    wire N__45728;
    wire N__45727;
    wire N__45726;
    wire N__45725;
    wire N__45722;
    wire N__45719;
    wire N__45718;
    wire N__45715;
    wire N__45712;
    wire N__45707;
    wire N__45704;
    wire N__45703;
    wire N__45698;
    wire N__45693;
    wire N__45690;
    wire N__45687;
    wire N__45684;
    wire N__45681;
    wire N__45674;
    wire N__45671;
    wire N__45668;
    wire N__45665;
    wire N__45664;
    wire N__45661;
    wire N__45660;
    wire N__45657;
    wire N__45654;
    wire N__45651;
    wire N__45644;
    wire N__45643;
    wire N__45640;
    wire N__45637;
    wire N__45632;
    wire N__45629;
    wire N__45626;
    wire N__45623;
    wire N__45620;
    wire N__45617;
    wire N__45614;
    wire N__45611;
    wire N__45610;
    wire N__45607;
    wire N__45604;
    wire N__45599;
    wire N__45596;
    wire N__45593;
    wire N__45590;
    wire N__45587;
    wire N__45584;
    wire N__45583;
    wire N__45580;
    wire N__45579;
    wire N__45576;
    wire N__45573;
    wire N__45570;
    wire N__45563;
    wire N__45560;
    wire N__45557;
    wire N__45554;
    wire N__45551;
    wire N__45548;
    wire N__45547;
    wire N__45544;
    wire N__45541;
    wire N__45538;
    wire N__45537;
    wire N__45534;
    wire N__45531;
    wire N__45528;
    wire N__45525;
    wire N__45522;
    wire N__45515;
    wire N__45512;
    wire N__45509;
    wire N__45506;
    wire N__45505;
    wire N__45504;
    wire N__45499;
    wire N__45496;
    wire N__45493;
    wire N__45488;
    wire N__45485;
    wire N__45482;
    wire N__45479;
    wire N__45478;
    wire N__45475;
    wire N__45472;
    wire N__45471;
    wire N__45466;
    wire N__45463;
    wire N__45460;
    wire N__45455;
    wire N__45452;
    wire N__45449;
    wire N__45446;
    wire N__45445;
    wire N__45442;
    wire N__45439;
    wire N__45438;
    wire N__45433;
    wire N__45430;
    wire N__45427;
    wire N__45422;
    wire N__45419;
    wire N__45416;
    wire N__45413;
    wire N__45410;
    wire N__45409;
    wire N__45408;
    wire N__45403;
    wire N__45400;
    wire N__45397;
    wire N__45392;
    wire N__45389;
    wire N__45386;
    wire N__45383;
    wire N__45380;
    wire N__45377;
    wire N__45376;
    wire N__45371;
    wire N__45370;
    wire N__45367;
    wire N__45364;
    wire N__45361;
    wire N__45356;
    wire N__45353;
    wire N__45350;
    wire N__45347;
    wire N__45344;
    wire N__45341;
    wire N__45340;
    wire N__45337;
    wire N__45336;
    wire N__45333;
    wire N__45330;
    wire N__45327;
    wire N__45324;
    wire N__45317;
    wire N__45314;
    wire N__45311;
    wire N__45308;
    wire N__45305;
    wire N__45302;
    wire N__45299;
    wire N__45298;
    wire N__45297;
    wire N__45294;
    wire N__45291;
    wire N__45288;
    wire N__45281;
    wire N__45278;
    wire N__45277;
    wire N__45274;
    wire N__45271;
    wire N__45266;
    wire N__45263;
    wire N__45260;
    wire N__45259;
    wire N__45256;
    wire N__45253;
    wire N__45252;
    wire N__45247;
    wire N__45244;
    wire N__45241;
    wire N__45236;
    wire N__45235;
    wire N__45232;
    wire N__45229;
    wire N__45226;
    wire N__45223;
    wire N__45220;
    wire N__45217;
    wire N__45212;
    wire N__45209;
    wire N__45208;
    wire N__45205;
    wire N__45202;
    wire N__45201;
    wire N__45196;
    wire N__45193;
    wire N__45190;
    wire N__45185;
    wire N__45182;
    wire N__45181;
    wire N__45176;
    wire N__45175;
    wire N__45172;
    wire N__45169;
    wire N__45166;
    wire N__45161;
    wire N__45160;
    wire N__45159;
    wire N__45156;
    wire N__45155;
    wire N__45154;
    wire N__45153;
    wire N__45150;
    wire N__45147;
    wire N__45144;
    wire N__45139;
    wire N__45134;
    wire N__45131;
    wire N__45128;
    wire N__45125;
    wire N__45122;
    wire N__45117;
    wire N__45114;
    wire N__45111;
    wire N__45104;
    wire N__45101;
    wire N__45100;
    wire N__45095;
    wire N__45094;
    wire N__45091;
    wire N__45088;
    wire N__45085;
    wire N__45080;
    wire N__45077;
    wire N__45076;
    wire N__45075;
    wire N__45072;
    wire N__45067;
    wire N__45062;
    wire N__45059;
    wire N__45056;
    wire N__45055;
    wire N__45052;
    wire N__45051;
    wire N__45048;
    wire N__45045;
    wire N__45042;
    wire N__45039;
    wire N__45036;
    wire N__45029;
    wire N__45026;
    wire N__45025;
    wire N__45024;
    wire N__45021;
    wire N__45018;
    wire N__45015;
    wire N__45008;
    wire N__45005;
    wire N__45004;
    wire N__45001;
    wire N__44998;
    wire N__44993;
    wire N__44992;
    wire N__44989;
    wire N__44986;
    wire N__44983;
    wire N__44978;
    wire N__44975;
    wire N__44974;
    wire N__44973;
    wire N__44970;
    wire N__44965;
    wire N__44960;
    wire N__44957;
    wire N__44954;
    wire N__44953;
    wire N__44950;
    wire N__44949;
    wire N__44946;
    wire N__44943;
    wire N__44940;
    wire N__44937;
    wire N__44930;
    wire N__44927;
    wire N__44926;
    wire N__44925;
    wire N__44922;
    wire N__44919;
    wire N__44916;
    wire N__44913;
    wire N__44910;
    wire N__44907;
    wire N__44900;
    wire N__44897;
    wire N__44894;
    wire N__44893;
    wire N__44890;
    wire N__44889;
    wire N__44886;
    wire N__44883;
    wire N__44880;
    wire N__44877;
    wire N__44870;
    wire N__44867;
    wire N__44866;
    wire N__44865;
    wire N__44862;
    wire N__44859;
    wire N__44856;
    wire N__44851;
    wire N__44846;
    wire N__44843;
    wire N__44842;
    wire N__44839;
    wire N__44836;
    wire N__44835;
    wire N__44830;
    wire N__44827;
    wire N__44824;
    wire N__44819;
    wire N__44816;
    wire N__44813;
    wire N__44812;
    wire N__44811;
    wire N__44808;
    wire N__44803;
    wire N__44800;
    wire N__44797;
    wire N__44792;
    wire N__44789;
    wire N__44788;
    wire N__44785;
    wire N__44782;
    wire N__44781;
    wire N__44776;
    wire N__44773;
    wire N__44770;
    wire N__44765;
    wire N__44762;
    wire N__44761;
    wire N__44760;
    wire N__44757;
    wire N__44752;
    wire N__44749;
    wire N__44746;
    wire N__44741;
    wire N__44738;
    wire N__44737;
    wire N__44732;
    wire N__44731;
    wire N__44728;
    wire N__44725;
    wire N__44722;
    wire N__44717;
    wire N__44716;
    wire N__44715;
    wire N__44712;
    wire N__44709;
    wire N__44706;
    wire N__44701;
    wire N__44698;
    wire N__44695;
    wire N__44692;
    wire N__44687;
    wire N__44684;
    wire N__44683;
    wire N__44678;
    wire N__44677;
    wire N__44674;
    wire N__44671;
    wire N__44668;
    wire N__44663;
    wire N__44662;
    wire N__44659;
    wire N__44656;
    wire N__44655;
    wire N__44652;
    wire N__44649;
    wire N__44646;
    wire N__44639;
    wire N__44636;
    wire N__44633;
    wire N__44630;
    wire N__44629;
    wire N__44626;
    wire N__44625;
    wire N__44622;
    wire N__44619;
    wire N__44616;
    wire N__44613;
    wire N__44610;
    wire N__44603;
    wire N__44602;
    wire N__44601;
    wire N__44598;
    wire N__44595;
    wire N__44594;
    wire N__44591;
    wire N__44586;
    wire N__44581;
    wire N__44576;
    wire N__44573;
    wire N__44570;
    wire N__44569;
    wire N__44566;
    wire N__44563;
    wire N__44558;
    wire N__44557;
    wire N__44554;
    wire N__44551;
    wire N__44548;
    wire N__44543;
    wire N__44542;
    wire N__44539;
    wire N__44536;
    wire N__44533;
    wire N__44530;
    wire N__44527;
    wire N__44524;
    wire N__44519;
    wire N__44516;
    wire N__44515;
    wire N__44512;
    wire N__44511;
    wire N__44508;
    wire N__44505;
    wire N__44502;
    wire N__44499;
    wire N__44492;
    wire N__44489;
    wire N__44488;
    wire N__44485;
    wire N__44482;
    wire N__44477;
    wire N__44474;
    wire N__44471;
    wire N__44468;
    wire N__44465;
    wire N__44462;
    wire N__44459;
    wire N__44456;
    wire N__44453;
    wire N__44450;
    wire N__44449;
    wire N__44446;
    wire N__44445;
    wire N__44444;
    wire N__44441;
    wire N__44438;
    wire N__44435;
    wire N__44432;
    wire N__44429;
    wire N__44424;
    wire N__44421;
    wire N__44418;
    wire N__44417;
    wire N__44414;
    wire N__44411;
    wire N__44408;
    wire N__44405;
    wire N__44402;
    wire N__44399;
    wire N__44394;
    wire N__44387;
    wire N__44386;
    wire N__44385;
    wire N__44384;
    wire N__44379;
    wire N__44376;
    wire N__44373;
    wire N__44370;
    wire N__44365;
    wire N__44362;
    wire N__44357;
    wire N__44354;
    wire N__44351;
    wire N__44348;
    wire N__44345;
    wire N__44342;
    wire N__44341;
    wire N__44338;
    wire N__44335;
    wire N__44330;
    wire N__44329;
    wire N__44326;
    wire N__44323;
    wire N__44318;
    wire N__44317;
    wire N__44314;
    wire N__44311;
    wire N__44308;
    wire N__44303;
    wire N__44302;
    wire N__44299;
    wire N__44296;
    wire N__44291;
    wire N__44288;
    wire N__44285;
    wire N__44282;
    wire N__44281;
    wire N__44278;
    wire N__44275;
    wire N__44274;
    wire N__44273;
    wire N__44270;
    wire N__44267;
    wire N__44264;
    wire N__44261;
    wire N__44260;
    wire N__44257;
    wire N__44254;
    wire N__44251;
    wire N__44248;
    wire N__44245;
    wire N__44236;
    wire N__44233;
    wire N__44230;
    wire N__44225;
    wire N__44222;
    wire N__44219;
    wire N__44216;
    wire N__44213;
    wire N__44210;
    wire N__44207;
    wire N__44206;
    wire N__44205;
    wire N__44204;
    wire N__44201;
    wire N__44200;
    wire N__44199;
    wire N__44198;
    wire N__44189;
    wire N__44188;
    wire N__44187;
    wire N__44186;
    wire N__44185;
    wire N__44184;
    wire N__44183;
    wire N__44182;
    wire N__44181;
    wire N__44180;
    wire N__44179;
    wire N__44178;
    wire N__44177;
    wire N__44174;
    wire N__44173;
    wire N__44170;
    wire N__44169;
    wire N__44168;
    wire N__44167;
    wire N__44166;
    wire N__44165;
    wire N__44164;
    wire N__44161;
    wire N__44158;
    wire N__44157;
    wire N__44156;
    wire N__44155;
    wire N__44154;
    wire N__44151;
    wire N__44148;
    wire N__44145;
    wire N__44144;
    wire N__44141;
    wire N__44140;
    wire N__44139;
    wire N__44126;
    wire N__44109;
    wire N__44100;
    wire N__44097;
    wire N__44094;
    wire N__44091;
    wire N__44088;
    wire N__44087;
    wire N__44086;
    wire N__44085;
    wire N__44084;
    wire N__44081;
    wire N__44066;
    wire N__44063;
    wire N__44062;
    wire N__44061;
    wire N__44060;
    wire N__44055;
    wire N__44052;
    wire N__44049;
    wire N__44046;
    wire N__44039;
    wire N__44034;
    wire N__44031;
    wire N__44028;
    wire N__44025;
    wire N__44018;
    wire N__44017;
    wire N__44014;
    wire N__44009;
    wire N__44006;
    wire N__44001;
    wire N__43998;
    wire N__43995;
    wire N__43990;
    wire N__43987;
    wire N__43984;
    wire N__43979;
    wire N__43976;
    wire N__43969;
    wire N__43958;
    wire N__43957;
    wire N__43956;
    wire N__43955;
    wire N__43954;
    wire N__43951;
    wire N__43948;
    wire N__43945;
    wire N__43942;
    wire N__43939;
    wire N__43936;
    wire N__43933;
    wire N__43930;
    wire N__43927;
    wire N__43924;
    wire N__43913;
    wire N__43912;
    wire N__43911;
    wire N__43910;
    wire N__43901;
    wire N__43900;
    wire N__43899;
    wire N__43898;
    wire N__43897;
    wire N__43896;
    wire N__43895;
    wire N__43894;
    wire N__43893;
    wire N__43892;
    wire N__43889;
    wire N__43888;
    wire N__43887;
    wire N__43880;
    wire N__43879;
    wire N__43878;
    wire N__43875;
    wire N__43864;
    wire N__43863;
    wire N__43862;
    wire N__43861;
    wire N__43860;
    wire N__43859;
    wire N__43858;
    wire N__43857;
    wire N__43856;
    wire N__43855;
    wire N__43854;
    wire N__43853;
    wire N__43852;
    wire N__43851;
    wire N__43850;
    wire N__43849;
    wire N__43848;
    wire N__43847;
    wire N__43846;
    wire N__43845;
    wire N__43844;
    wire N__43841;
    wire N__43836;
    wire N__43833;
    wire N__43828;
    wire N__43827;
    wire N__43824;
    wire N__43821;
    wire N__43804;
    wire N__43795;
    wire N__43792;
    wire N__43777;
    wire N__43772;
    wire N__43767;
    wire N__43764;
    wire N__43761;
    wire N__43754;
    wire N__43749;
    wire N__43746;
    wire N__43741;
    wire N__43730;
    wire N__43727;
    wire N__43724;
    wire N__43721;
    wire N__43718;
    wire N__43715;
    wire N__43712;
    wire N__43711;
    wire N__43708;
    wire N__43707;
    wire N__43704;
    wire N__43701;
    wire N__43700;
    wire N__43697;
    wire N__43694;
    wire N__43691;
    wire N__43688;
    wire N__43687;
    wire N__43684;
    wire N__43681;
    wire N__43676;
    wire N__43673;
    wire N__43670;
    wire N__43667;
    wire N__43662;
    wire N__43659;
    wire N__43654;
    wire N__43649;
    wire N__43648;
    wire N__43647;
    wire N__43646;
    wire N__43645;
    wire N__43642;
    wire N__43639;
    wire N__43638;
    wire N__43635;
    wire N__43632;
    wire N__43623;
    wire N__43620;
    wire N__43619;
    wire N__43612;
    wire N__43609;
    wire N__43604;
    wire N__43603;
    wire N__43602;
    wire N__43601;
    wire N__43598;
    wire N__43595;
    wire N__43594;
    wire N__43593;
    wire N__43592;
    wire N__43591;
    wire N__43588;
    wire N__43585;
    wire N__43582;
    wire N__43577;
    wire N__43566;
    wire N__43563;
    wire N__43560;
    wire N__43553;
    wire N__43550;
    wire N__43547;
    wire N__43546;
    wire N__43545;
    wire N__43544;
    wire N__43543;
    wire N__43542;
    wire N__43541;
    wire N__43538;
    wire N__43527;
    wire N__43524;
    wire N__43523;
    wire N__43520;
    wire N__43517;
    wire N__43514;
    wire N__43511;
    wire N__43502;
    wire N__43501;
    wire N__43498;
    wire N__43497;
    wire N__43494;
    wire N__43491;
    wire N__43488;
    wire N__43485;
    wire N__43480;
    wire N__43477;
    wire N__43474;
    wire N__43471;
    wire N__43468;
    wire N__43463;
    wire N__43462;
    wire N__43461;
    wire N__43458;
    wire N__43455;
    wire N__43452;
    wire N__43451;
    wire N__43448;
    wire N__43445;
    wire N__43442;
    wire N__43439;
    wire N__43434;
    wire N__43429;
    wire N__43424;
    wire N__43423;
    wire N__43420;
    wire N__43419;
    wire N__43416;
    wire N__43413;
    wire N__43410;
    wire N__43403;
    wire N__43402;
    wire N__43401;
    wire N__43398;
    wire N__43395;
    wire N__43392;
    wire N__43389;
    wire N__43386;
    wire N__43383;
    wire N__43380;
    wire N__43377;
    wire N__43370;
    wire N__43367;
    wire N__43366;
    wire N__43363;
    wire N__43362;
    wire N__43359;
    wire N__43356;
    wire N__43353;
    wire N__43346;
    wire N__43345;
    wire N__43344;
    wire N__43343;
    wire N__43338;
    wire N__43335;
    wire N__43334;
    wire N__43333;
    wire N__43330;
    wire N__43327;
    wire N__43320;
    wire N__43317;
    wire N__43314;
    wire N__43311;
    wire N__43304;
    wire N__43301;
    wire N__43298;
    wire N__43297;
    wire N__43296;
    wire N__43293;
    wire N__43290;
    wire N__43289;
    wire N__43286;
    wire N__43283;
    wire N__43280;
    wire N__43275;
    wire N__43272;
    wire N__43267;
    wire N__43264;
    wire N__43261;
    wire N__43256;
    wire N__43255;
    wire N__43254;
    wire N__43253;
    wire N__43246;
    wire N__43243;
    wire N__43242;
    wire N__43241;
    wire N__43240;
    wire N__43239;
    wire N__43236;
    wire N__43233;
    wire N__43230;
    wire N__43225;
    wire N__43222;
    wire N__43211;
    wire N__43210;
    wire N__43207;
    wire N__43206;
    wire N__43205;
    wire N__43202;
    wire N__43199;
    wire N__43194;
    wire N__43191;
    wire N__43186;
    wire N__43183;
    wire N__43180;
    wire N__43175;
    wire N__43172;
    wire N__43169;
    wire N__43166;
    wire N__43163;
    wire N__43160;
    wire N__43157;
    wire N__43154;
    wire N__43153;
    wire N__43152;
    wire N__43151;
    wire N__43150;
    wire N__43147;
    wire N__43144;
    wire N__43141;
    wire N__43136;
    wire N__43127;
    wire N__43124;
    wire N__43121;
    wire N__43118;
    wire N__43117;
    wire N__43114;
    wire N__43111;
    wire N__43106;
    wire N__43103;
    wire N__43100;
    wire N__43097;
    wire N__43096;
    wire N__43093;
    wire N__43090;
    wire N__43087;
    wire N__43084;
    wire N__43081;
    wire N__43078;
    wire N__43077;
    wire N__43076;
    wire N__43071;
    wire N__43068;
    wire N__43065;
    wire N__43060;
    wire N__43055;
    wire N__43054;
    wire N__43051;
    wire N__43050;
    wire N__43043;
    wire N__43040;
    wire N__43037;
    wire N__43034;
    wire N__43033;
    wire N__43030;
    wire N__43027;
    wire N__43024;
    wire N__43023;
    wire N__43020;
    wire N__43017;
    wire N__43014;
    wire N__43011;
    wire N__43004;
    wire N__43003;
    wire N__42998;
    wire N__42995;
    wire N__42992;
    wire N__42989;
    wire N__42986;
    wire N__42983;
    wire N__42982;
    wire N__42981;
    wire N__42980;
    wire N__42971;
    wire N__42970;
    wire N__42969;
    wire N__42968;
    wire N__42967;
    wire N__42966;
    wire N__42965;
    wire N__42964;
    wire N__42963;
    wire N__42962;
    wire N__42961;
    wire N__42960;
    wire N__42959;
    wire N__42958;
    wire N__42957;
    wire N__42956;
    wire N__42955;
    wire N__42954;
    wire N__42953;
    wire N__42952;
    wire N__42951;
    wire N__42950;
    wire N__42949;
    wire N__42948;
    wire N__42947;
    wire N__42946;
    wire N__42945;
    wire N__42942;
    wire N__42937;
    wire N__42928;
    wire N__42919;
    wire N__42910;
    wire N__42901;
    wire N__42892;
    wire N__42883;
    wire N__42878;
    wire N__42873;
    wire N__42860;
    wire N__42857;
    wire N__42856;
    wire N__42853;
    wire N__42850;
    wire N__42849;
    wire N__42846;
    wire N__42843;
    wire N__42840;
    wire N__42839;
    wire N__42832;
    wire N__42829;
    wire N__42826;
    wire N__42823;
    wire N__42818;
    wire N__42815;
    wire N__42812;
    wire N__42809;
    wire N__42806;
    wire N__42803;
    wire N__42800;
    wire N__42797;
    wire N__42796;
    wire N__42793;
    wire N__42790;
    wire N__42789;
    wire N__42786;
    wire N__42783;
    wire N__42780;
    wire N__42775;
    wire N__42770;
    wire N__42769;
    wire N__42768;
    wire N__42765;
    wire N__42764;
    wire N__42761;
    wire N__42758;
    wire N__42755;
    wire N__42752;
    wire N__42749;
    wire N__42744;
    wire N__42737;
    wire N__42734;
    wire N__42731;
    wire N__42728;
    wire N__42725;
    wire N__42722;
    wire N__42719;
    wire N__42716;
    wire N__42713;
    wire N__42710;
    wire N__42707;
    wire N__42704;
    wire N__42701;
    wire N__42698;
    wire N__42695;
    wire N__42692;
    wire N__42689;
    wire N__42686;
    wire N__42683;
    wire N__42682;
    wire N__42679;
    wire N__42676;
    wire N__42671;
    wire N__42668;
    wire N__42667;
    wire N__42664;
    wire N__42661;
    wire N__42658;
    wire N__42653;
    wire N__42652;
    wire N__42651;
    wire N__42650;
    wire N__42649;
    wire N__42648;
    wire N__42647;
    wire N__42646;
    wire N__42645;
    wire N__42644;
    wire N__42641;
    wire N__42640;
    wire N__42637;
    wire N__42636;
    wire N__42633;
    wire N__42632;
    wire N__42631;
    wire N__42630;
    wire N__42629;
    wire N__42628;
    wire N__42627;
    wire N__42626;
    wire N__42625;
    wire N__42624;
    wire N__42623;
    wire N__42622;
    wire N__42621;
    wire N__42620;
    wire N__42615;
    wire N__42612;
    wire N__42605;
    wire N__42594;
    wire N__42583;
    wire N__42574;
    wire N__42571;
    wire N__42564;
    wire N__42561;
    wire N__42560;
    wire N__42559;
    wire N__42558;
    wire N__42555;
    wire N__42552;
    wire N__42551;
    wire N__42544;
    wire N__42535;
    wire N__42528;
    wire N__42527;
    wire N__42526;
    wire N__42525;
    wire N__42522;
    wire N__42519;
    wire N__42516;
    wire N__42509;
    wire N__42502;
    wire N__42491;
    wire N__42488;
    wire N__42485;
    wire N__42482;
    wire N__42481;
    wire N__42480;
    wire N__42477;
    wire N__42472;
    wire N__42467;
    wire N__42466;
    wire N__42465;
    wire N__42464;
    wire N__42463;
    wire N__42462;
    wire N__42461;
    wire N__42454;
    wire N__42447;
    wire N__42446;
    wire N__42445;
    wire N__42444;
    wire N__42443;
    wire N__42442;
    wire N__42441;
    wire N__42440;
    wire N__42439;
    wire N__42438;
    wire N__42435;
    wire N__42432;
    wire N__42429;
    wire N__42422;
    wire N__42421;
    wire N__42420;
    wire N__42419;
    wire N__42418;
    wire N__42417;
    wire N__42412;
    wire N__42403;
    wire N__42400;
    wire N__42393;
    wire N__42384;
    wire N__42381;
    wire N__42380;
    wire N__42379;
    wire N__42378;
    wire N__42375;
    wire N__42372;
    wire N__42363;
    wire N__42356;
    wire N__42347;
    wire N__42346;
    wire N__42343;
    wire N__42340;
    wire N__42339;
    wire N__42336;
    wire N__42333;
    wire N__42330;
    wire N__42329;
    wire N__42326;
    wire N__42323;
    wire N__42320;
    wire N__42319;
    wire N__42316;
    wire N__42311;
    wire N__42308;
    wire N__42305;
    wire N__42296;
    wire N__42293;
    wire N__42290;
    wire N__42287;
    wire N__42284;
    wire N__42281;
    wire N__42278;
    wire N__42275;
    wire N__42274;
    wire N__42271;
    wire N__42268;
    wire N__42265;
    wire N__42260;
    wire N__42259;
    wire N__42256;
    wire N__42253;
    wire N__42250;
    wire N__42247;
    wire N__42244;
    wire N__42243;
    wire N__42240;
    wire N__42237;
    wire N__42234;
    wire N__42233;
    wire N__42230;
    wire N__42225;
    wire N__42222;
    wire N__42219;
    wire N__42216;
    wire N__42209;
    wire N__42206;
    wire N__42205;
    wire N__42204;
    wire N__42201;
    wire N__42196;
    wire N__42191;
    wire N__42190;
    wire N__42187;
    wire N__42184;
    wire N__42183;
    wire N__42182;
    wire N__42181;
    wire N__42178;
    wire N__42175;
    wire N__42172;
    wire N__42169;
    wire N__42166;
    wire N__42163;
    wire N__42160;
    wire N__42157;
    wire N__42154;
    wire N__42151;
    wire N__42148;
    wire N__42141;
    wire N__42134;
    wire N__42131;
    wire N__42130;
    wire N__42129;
    wire N__42126;
    wire N__42123;
    wire N__42120;
    wire N__42117;
    wire N__42114;
    wire N__42111;
    wire N__42104;
    wire N__42103;
    wire N__42102;
    wire N__42101;
    wire N__42100;
    wire N__42099;
    wire N__42094;
    wire N__42093;
    wire N__42092;
    wire N__42089;
    wire N__42082;
    wire N__42079;
    wire N__42076;
    wire N__42073;
    wire N__42070;
    wire N__42067;
    wire N__42062;
    wire N__42053;
    wire N__42050;
    wire N__42049;
    wire N__42048;
    wire N__42045;
    wire N__42042;
    wire N__42039;
    wire N__42036;
    wire N__42033;
    wire N__42028;
    wire N__42025;
    wire N__42020;
    wire N__42019;
    wire N__42014;
    wire N__42013;
    wire N__42010;
    wire N__42007;
    wire N__42004;
    wire N__41999;
    wire N__41998;
    wire N__41995;
    wire N__41992;
    wire N__41991;
    wire N__41988;
    wire N__41985;
    wire N__41982;
    wire N__41979;
    wire N__41976;
    wire N__41973;
    wire N__41966;
    wire N__41963;
    wire N__41960;
    wire N__41957;
    wire N__41954;
    wire N__41951;
    wire N__41948;
    wire N__41945;
    wire N__41942;
    wire N__41939;
    wire N__41936;
    wire N__41933;
    wire N__41932;
    wire N__41931;
    wire N__41930;
    wire N__41927;
    wire N__41922;
    wire N__41919;
    wire N__41916;
    wire N__41913;
    wire N__41910;
    wire N__41907;
    wire N__41904;
    wire N__41901;
    wire N__41894;
    wire N__41891;
    wire N__41888;
    wire N__41887;
    wire N__41886;
    wire N__41883;
    wire N__41880;
    wire N__41877;
    wire N__41876;
    wire N__41873;
    wire N__41870;
    wire N__41867;
    wire N__41864;
    wire N__41861;
    wire N__41856;
    wire N__41853;
    wire N__41850;
    wire N__41847;
    wire N__41844;
    wire N__41837;
    wire N__41836;
    wire N__41833;
    wire N__41830;
    wire N__41825;
    wire N__41824;
    wire N__41821;
    wire N__41818;
    wire N__41813;
    wire N__41810;
    wire N__41809;
    wire N__41804;
    wire N__41801;
    wire N__41798;
    wire N__41797;
    wire N__41794;
    wire N__41793;
    wire N__41792;
    wire N__41789;
    wire N__41786;
    wire N__41783;
    wire N__41780;
    wire N__41777;
    wire N__41768;
    wire N__41767;
    wire N__41764;
    wire N__41763;
    wire N__41760;
    wire N__41757;
    wire N__41756;
    wire N__41753;
    wire N__41750;
    wire N__41747;
    wire N__41744;
    wire N__41741;
    wire N__41740;
    wire N__41737;
    wire N__41734;
    wire N__41731;
    wire N__41728;
    wire N__41725;
    wire N__41722;
    wire N__41715;
    wire N__41708;
    wire N__41705;
    wire N__41702;
    wire N__41699;
    wire N__41698;
    wire N__41697;
    wire N__41696;
    wire N__41693;
    wire N__41690;
    wire N__41687;
    wire N__41684;
    wire N__41675;
    wire N__41672;
    wire N__41671;
    wire N__41670;
    wire N__41667;
    wire N__41664;
    wire N__41661;
    wire N__41660;
    wire N__41655;
    wire N__41652;
    wire N__41649;
    wire N__41648;
    wire N__41645;
    wire N__41640;
    wire N__41637;
    wire N__41634;
    wire N__41631;
    wire N__41624;
    wire N__41621;
    wire N__41618;
    wire N__41615;
    wire N__41612;
    wire N__41609;
    wire N__41606;
    wire N__41603;
    wire N__41600;
    wire N__41597;
    wire N__41594;
    wire N__41591;
    wire N__41588;
    wire N__41585;
    wire N__41582;
    wire N__41579;
    wire N__41576;
    wire N__41575;
    wire N__41572;
    wire N__41569;
    wire N__41568;
    wire N__41567;
    wire N__41564;
    wire N__41559;
    wire N__41556;
    wire N__41551;
    wire N__41548;
    wire N__41545;
    wire N__41540;
    wire N__41537;
    wire N__41534;
    wire N__41531;
    wire N__41528;
    wire N__41527;
    wire N__41524;
    wire N__41521;
    wire N__41520;
    wire N__41517;
    wire N__41514;
    wire N__41511;
    wire N__41504;
    wire N__41501;
    wire N__41498;
    wire N__41495;
    wire N__41492;
    wire N__41491;
    wire N__41490;
    wire N__41489;
    wire N__41486;
    wire N__41485;
    wire N__41484;
    wire N__41483;
    wire N__41482;
    wire N__41481;
    wire N__41480;
    wire N__41479;
    wire N__41476;
    wire N__41473;
    wire N__41470;
    wire N__41457;
    wire N__41454;
    wire N__41453;
    wire N__41452;
    wire N__41451;
    wire N__41448;
    wire N__41447;
    wire N__41444;
    wire N__41441;
    wire N__41438;
    wire N__41437;
    wire N__41434;
    wire N__41425;
    wire N__41420;
    wire N__41415;
    wire N__41412;
    wire N__41409;
    wire N__41406;
    wire N__41393;
    wire N__41390;
    wire N__41387;
    wire N__41384;
    wire N__41381;
    wire N__41378;
    wire N__41375;
    wire N__41372;
    wire N__41369;
    wire N__41366;
    wire N__41363;
    wire N__41360;
    wire N__41357;
    wire N__41354;
    wire N__41351;
    wire N__41348;
    wire N__41345;
    wire N__41342;
    wire N__41339;
    wire N__41336;
    wire N__41333;
    wire N__41330;
    wire N__41327;
    wire N__41324;
    wire N__41321;
    wire N__41318;
    wire N__41315;
    wire N__41312;
    wire N__41309;
    wire N__41306;
    wire N__41303;
    wire N__41300;
    wire N__41297;
    wire N__41294;
    wire N__41291;
    wire N__41288;
    wire N__41285;
    wire N__41282;
    wire N__41279;
    wire N__41276;
    wire N__41275;
    wire N__41272;
    wire N__41269;
    wire N__41266;
    wire N__41263;
    wire N__41260;
    wire N__41257;
    wire N__41254;
    wire N__41253;
    wire N__41252;
    wire N__41249;
    wire N__41248;
    wire N__41245;
    wire N__41242;
    wire N__41239;
    wire N__41236;
    wire N__41233;
    wire N__41228;
    wire N__41225;
    wire N__41220;
    wire N__41217;
    wire N__41210;
    wire N__41207;
    wire N__41204;
    wire N__41201;
    wire N__41198;
    wire N__41195;
    wire N__41192;
    wire N__41189;
    wire N__41186;
    wire N__41183;
    wire N__41180;
    wire N__41177;
    wire N__41174;
    wire N__41171;
    wire N__41168;
    wire N__41165;
    wire N__41162;
    wire N__41159;
    wire N__41156;
    wire N__41153;
    wire N__41150;
    wire N__41147;
    wire N__41144;
    wire N__41141;
    wire N__41138;
    wire N__41135;
    wire N__41132;
    wire N__41129;
    wire N__41126;
    wire N__41123;
    wire N__41120;
    wire N__41117;
    wire N__41114;
    wire N__41111;
    wire N__41108;
    wire N__41105;
    wire N__41102;
    wire N__41099;
    wire N__41096;
    wire N__41093;
    wire N__41090;
    wire N__41087;
    wire N__41084;
    wire N__41081;
    wire N__41078;
    wire N__41075;
    wire N__41072;
    wire N__41069;
    wire N__41068;
    wire N__41067;
    wire N__41066;
    wire N__41065;
    wire N__41064;
    wire N__41063;
    wire N__41062;
    wire N__41061;
    wire N__41060;
    wire N__41059;
    wire N__41058;
    wire N__41055;
    wire N__41054;
    wire N__41053;
    wire N__41046;
    wire N__41037;
    wire N__41030;
    wire N__41029;
    wire N__41028;
    wire N__41027;
    wire N__41026;
    wire N__41023;
    wire N__41022;
    wire N__41021;
    wire N__41018;
    wire N__41015;
    wire N__41012;
    wire N__41009;
    wire N__41004;
    wire N__41001;
    wire N__41000;
    wire N__40999;
    wire N__40998;
    wire N__40991;
    wire N__40988;
    wire N__40985;
    wire N__40982;
    wire N__40981;
    wire N__40970;
    wire N__40961;
    wire N__40956;
    wire N__40953;
    wire N__40950;
    wire N__40947;
    wire N__40942;
    wire N__40937;
    wire N__40934;
    wire N__40929;
    wire N__40926;
    wire N__40919;
    wire N__40918;
    wire N__40917;
    wire N__40916;
    wire N__40915;
    wire N__40914;
    wire N__40911;
    wire N__40910;
    wire N__40909;
    wire N__40906;
    wire N__40903;
    wire N__40902;
    wire N__40901;
    wire N__40900;
    wire N__40899;
    wire N__40896;
    wire N__40895;
    wire N__40894;
    wire N__40891;
    wire N__40888;
    wire N__40885;
    wire N__40882;
    wire N__40879;
    wire N__40876;
    wire N__40873;
    wire N__40872;
    wire N__40869;
    wire N__40866;
    wire N__40863;
    wire N__40862;
    wire N__40861;
    wire N__40860;
    wire N__40859;
    wire N__40858;
    wire N__40857;
    wire N__40854;
    wire N__40853;
    wire N__40852;
    wire N__40849;
    wire N__40842;
    wire N__40839;
    wire N__40836;
    wire N__40831;
    wire N__40826;
    wire N__40821;
    wire N__40812;
    wire N__40803;
    wire N__40802;
    wire N__40795;
    wire N__40792;
    wire N__40789;
    wire N__40784;
    wire N__40775;
    wire N__40772;
    wire N__40769;
    wire N__40766;
    wire N__40763;
    wire N__40760;
    wire N__40755;
    wire N__40752;
    wire N__40739;
    wire N__40738;
    wire N__40735;
    wire N__40732;
    wire N__40729;
    wire N__40728;
    wire N__40725;
    wire N__40722;
    wire N__40719;
    wire N__40718;
    wire N__40717;
    wire N__40716;
    wire N__40713;
    wire N__40708;
    wire N__40705;
    wire N__40700;
    wire N__40691;
    wire N__40690;
    wire N__40687;
    wire N__40684;
    wire N__40683;
    wire N__40682;
    wire N__40681;
    wire N__40680;
    wire N__40679;
    wire N__40674;
    wire N__40671;
    wire N__40668;
    wire N__40667;
    wire N__40666;
    wire N__40665;
    wire N__40664;
    wire N__40663;
    wire N__40656;
    wire N__40655;
    wire N__40650;
    wire N__40647;
    wire N__40644;
    wire N__40641;
    wire N__40640;
    wire N__40637;
    wire N__40636;
    wire N__40635;
    wire N__40634;
    wire N__40633;
    wire N__40632;
    wire N__40631;
    wire N__40630;
    wire N__40629;
    wire N__40628;
    wire N__40625;
    wire N__40622;
    wire N__40619;
    wire N__40616;
    wire N__40611;
    wire N__40604;
    wire N__40595;
    wire N__40588;
    wire N__40583;
    wire N__40580;
    wire N__40579;
    wire N__40572;
    wire N__40569;
    wire N__40564;
    wire N__40557;
    wire N__40554;
    wire N__40551;
    wire N__40548;
    wire N__40543;
    wire N__40538;
    wire N__40529;
    wire N__40526;
    wire N__40523;
    wire N__40522;
    wire N__40519;
    wire N__40518;
    wire N__40515;
    wire N__40514;
    wire N__40511;
    wire N__40508;
    wire N__40505;
    wire N__40502;
    wire N__40499;
    wire N__40496;
    wire N__40491;
    wire N__40488;
    wire N__40485;
    wire N__40482;
    wire N__40475;
    wire N__40472;
    wire N__40469;
    wire N__40466;
    wire N__40463;
    wire N__40460;
    wire N__40457;
    wire N__40454;
    wire N__40453;
    wire N__40450;
    wire N__40447;
    wire N__40444;
    wire N__40441;
    wire N__40440;
    wire N__40439;
    wire N__40436;
    wire N__40433;
    wire N__40430;
    wire N__40429;
    wire N__40426;
    wire N__40419;
    wire N__40414;
    wire N__40409;
    wire N__40406;
    wire N__40403;
    wire N__40400;
    wire N__40397;
    wire N__40394;
    wire N__40393;
    wire N__40390;
    wire N__40389;
    wire N__40386;
    wire N__40383;
    wire N__40380;
    wire N__40377;
    wire N__40374;
    wire N__40371;
    wire N__40368;
    wire N__40365;
    wire N__40360;
    wire N__40355;
    wire N__40352;
    wire N__40349;
    wire N__40346;
    wire N__40345;
    wire N__40344;
    wire N__40343;
    wire N__40342;
    wire N__40337;
    wire N__40336;
    wire N__40335;
    wire N__40332;
    wire N__40329;
    wire N__40328;
    wire N__40327;
    wire N__40326;
    wire N__40323;
    wire N__40320;
    wire N__40319;
    wire N__40318;
    wire N__40317;
    wire N__40316;
    wire N__40311;
    wire N__40308;
    wire N__40299;
    wire N__40296;
    wire N__40293;
    wire N__40284;
    wire N__40281;
    wire N__40278;
    wire N__40275;
    wire N__40272;
    wire N__40269;
    wire N__40262;
    wire N__40259;
    wire N__40250;
    wire N__40249;
    wire N__40248;
    wire N__40245;
    wire N__40242;
    wire N__40239;
    wire N__40236;
    wire N__40233;
    wire N__40230;
    wire N__40225;
    wire N__40222;
    wire N__40217;
    wire N__40216;
    wire N__40215;
    wire N__40210;
    wire N__40207;
    wire N__40206;
    wire N__40205;
    wire N__40202;
    wire N__40195;
    wire N__40192;
    wire N__40189;
    wire N__40186;
    wire N__40183;
    wire N__40178;
    wire N__40177;
    wire N__40174;
    wire N__40171;
    wire N__40168;
    wire N__40165;
    wire N__40164;
    wire N__40161;
    wire N__40158;
    wire N__40155;
    wire N__40150;
    wire N__40147;
    wire N__40142;
    wire N__40139;
    wire N__40138;
    wire N__40135;
    wire N__40132;
    wire N__40129;
    wire N__40126;
    wire N__40121;
    wire N__40118;
    wire N__40117;
    wire N__40114;
    wire N__40111;
    wire N__40108;
    wire N__40105;
    wire N__40102;
    wire N__40099;
    wire N__40094;
    wire N__40093;
    wire N__40092;
    wire N__40089;
    wire N__40084;
    wire N__40081;
    wire N__40078;
    wire N__40075;
    wire N__40072;
    wire N__40067;
    wire N__40066;
    wire N__40065;
    wire N__40064;
    wire N__40061;
    wire N__40056;
    wire N__40053;
    wire N__40050;
    wire N__40047;
    wire N__40044;
    wire N__40041;
    wire N__40040;
    wire N__40039;
    wire N__40036;
    wire N__40031;
    wire N__40026;
    wire N__40019;
    wire N__40018;
    wire N__40017;
    wire N__40016;
    wire N__40015;
    wire N__40014;
    wire N__40013;
    wire N__40012;
    wire N__40011;
    wire N__40008;
    wire N__40007;
    wire N__40006;
    wire N__40003;
    wire N__40002;
    wire N__40001;
    wire N__39998;
    wire N__39995;
    wire N__39994;
    wire N__39991;
    wire N__39990;
    wire N__39989;
    wire N__39988;
    wire N__39985;
    wire N__39982;
    wire N__39979;
    wire N__39978;
    wire N__39977;
    wire N__39972;
    wire N__39969;
    wire N__39966;
    wire N__39963;
    wire N__39962;
    wire N__39961;
    wire N__39946;
    wire N__39933;
    wire N__39932;
    wire N__39929;
    wire N__39928;
    wire N__39925;
    wire N__39920;
    wire N__39917;
    wire N__39914;
    wire N__39911;
    wire N__39910;
    wire N__39907;
    wire N__39904;
    wire N__39899;
    wire N__39896;
    wire N__39893;
    wire N__39890;
    wire N__39883;
    wire N__39880;
    wire N__39873;
    wire N__39870;
    wire N__39863;
    wire N__39854;
    wire N__39853;
    wire N__39852;
    wire N__39851;
    wire N__39850;
    wire N__39849;
    wire N__39848;
    wire N__39847;
    wire N__39846;
    wire N__39845;
    wire N__39842;
    wire N__39839;
    wire N__39836;
    wire N__39833;
    wire N__39830;
    wire N__39827;
    wire N__39824;
    wire N__39823;
    wire N__39822;
    wire N__39821;
    wire N__39820;
    wire N__39819;
    wire N__39818;
    wire N__39813;
    wire N__39812;
    wire N__39811;
    wire N__39808;
    wire N__39799;
    wire N__39792;
    wire N__39785;
    wire N__39778;
    wire N__39775;
    wire N__39770;
    wire N__39769;
    wire N__39768;
    wire N__39767;
    wire N__39766;
    wire N__39755;
    wire N__39750;
    wire N__39747;
    wire N__39744;
    wire N__39739;
    wire N__39738;
    wire N__39735;
    wire N__39732;
    wire N__39729;
    wire N__39726;
    wire N__39723;
    wire N__39720;
    wire N__39719;
    wire N__39716;
    wire N__39713;
    wire N__39710;
    wire N__39705;
    wire N__39700;
    wire N__39697;
    wire N__39694;
    wire N__39689;
    wire N__39680;
    wire N__39679;
    wire N__39678;
    wire N__39675;
    wire N__39670;
    wire N__39669;
    wire N__39668;
    wire N__39667;
    wire N__39666;
    wire N__39665;
    wire N__39664;
    wire N__39663;
    wire N__39662;
    wire N__39661;
    wire N__39660;
    wire N__39659;
    wire N__39658;
    wire N__39657;
    wire N__39656;
    wire N__39655;
    wire N__39654;
    wire N__39651;
    wire N__39648;
    wire N__39645;
    wire N__39642;
    wire N__39629;
    wire N__39614;
    wire N__39611;
    wire N__39610;
    wire N__39609;
    wire N__39608;
    wire N__39601;
    wire N__39594;
    wire N__39591;
    wire N__39588;
    wire N__39583;
    wire N__39580;
    wire N__39577;
    wire N__39570;
    wire N__39569;
    wire N__39568;
    wire N__39565;
    wire N__39562;
    wire N__39559;
    wire N__39554;
    wire N__39551;
    wire N__39548;
    wire N__39545;
    wire N__39536;
    wire N__39535;
    wire N__39532;
    wire N__39529;
    wire N__39524;
    wire N__39521;
    wire N__39518;
    wire N__39515;
    wire N__39514;
    wire N__39513;
    wire N__39512;
    wire N__39503;
    wire N__39500;
    wire N__39497;
    wire N__39496;
    wire N__39493;
    wire N__39490;
    wire N__39489;
    wire N__39486;
    wire N__39483;
    wire N__39480;
    wire N__39473;
    wire N__39470;
    wire N__39469;
    wire N__39466;
    wire N__39463;
    wire N__39462;
    wire N__39459;
    wire N__39456;
    wire N__39453;
    wire N__39446;
    wire N__39443;
    wire N__39440;
    wire N__39437;
    wire N__39434;
    wire N__39431;
    wire N__39428;
    wire N__39425;
    wire N__39422;
    wire N__39419;
    wire N__39416;
    wire N__39413;
    wire N__39410;
    wire N__39407;
    wire N__39406;
    wire N__39405;
    wire N__39402;
    wire N__39401;
    wire N__39398;
    wire N__39395;
    wire N__39392;
    wire N__39389;
    wire N__39386;
    wire N__39383;
    wire N__39380;
    wire N__39379;
    wire N__39376;
    wire N__39373;
    wire N__39368;
    wire N__39365;
    wire N__39362;
    wire N__39353;
    wire N__39352;
    wire N__39351;
    wire N__39350;
    wire N__39347;
    wire N__39344;
    wire N__39341;
    wire N__39338;
    wire N__39335;
    wire N__39332;
    wire N__39331;
    wire N__39328;
    wire N__39325;
    wire N__39322;
    wire N__39319;
    wire N__39316;
    wire N__39313;
    wire N__39302;
    wire N__39299;
    wire N__39296;
    wire N__39293;
    wire N__39290;
    wire N__39287;
    wire N__39284;
    wire N__39281;
    wire N__39278;
    wire N__39275;
    wire N__39272;
    wire N__39269;
    wire N__39266;
    wire N__39263;
    wire N__39260;
    wire N__39259;
    wire N__39256;
    wire N__39255;
    wire N__39254;
    wire N__39251;
    wire N__39248;
    wire N__39243;
    wire N__39240;
    wire N__39233;
    wire N__39232;
    wire N__39231;
    wire N__39228;
    wire N__39225;
    wire N__39222;
    wire N__39217;
    wire N__39212;
    wire N__39209;
    wire N__39208;
    wire N__39207;
    wire N__39204;
    wire N__39201;
    wire N__39198;
    wire N__39193;
    wire N__39188;
    wire N__39185;
    wire N__39184;
    wire N__39183;
    wire N__39180;
    wire N__39177;
    wire N__39174;
    wire N__39171;
    wire N__39164;
    wire N__39161;
    wire N__39160;
    wire N__39159;
    wire N__39156;
    wire N__39153;
    wire N__39150;
    wire N__39147;
    wire N__39140;
    wire N__39137;
    wire N__39136;
    wire N__39135;
    wire N__39132;
    wire N__39129;
    wire N__39126;
    wire N__39121;
    wire N__39116;
    wire N__39113;
    wire N__39112;
    wire N__39111;
    wire N__39108;
    wire N__39105;
    wire N__39102;
    wire N__39097;
    wire N__39092;
    wire N__39089;
    wire N__39088;
    wire N__39085;
    wire N__39082;
    wire N__39077;
    wire N__39074;
    wire N__39073;
    wire N__39072;
    wire N__39071;
    wire N__39070;
    wire N__39069;
    wire N__39068;
    wire N__39067;
    wire N__39066;
    wire N__39065;
    wire N__39064;
    wire N__39063;
    wire N__39062;
    wire N__39061;
    wire N__39060;
    wire N__39059;
    wire N__39058;
    wire N__39057;
    wire N__39056;
    wire N__39055;
    wire N__39054;
    wire N__39053;
    wire N__39052;
    wire N__39051;
    wire N__39050;
    wire N__39049;
    wire N__39044;
    wire N__39035;
    wire N__39034;
    wire N__39033;
    wire N__39032;
    wire N__39031;
    wire N__39022;
    wire N__39013;
    wire N__39004;
    wire N__38995;
    wire N__38986;
    wire N__38983;
    wire N__38980;
    wire N__38971;
    wire N__38962;
    wire N__38959;
    wire N__38956;
    wire N__38953;
    wire N__38948;
    wire N__38939;
    wire N__38936;
    wire N__38935;
    wire N__38932;
    wire N__38929;
    wire N__38924;
    wire N__38921;
    wire N__38918;
    wire N__38917;
    wire N__38916;
    wire N__38913;
    wire N__38910;
    wire N__38909;
    wire N__38906;
    wire N__38901;
    wire N__38898;
    wire N__38895;
    wire N__38890;
    wire N__38887;
    wire N__38884;
    wire N__38879;
    wire N__38878;
    wire N__38877;
    wire N__38874;
    wire N__38871;
    wire N__38868;
    wire N__38863;
    wire N__38858;
    wire N__38855;
    wire N__38854;
    wire N__38853;
    wire N__38850;
    wire N__38847;
    wire N__38844;
    wire N__38839;
    wire N__38834;
    wire N__38831;
    wire N__38830;
    wire N__38829;
    wire N__38826;
    wire N__38823;
    wire N__38820;
    wire N__38817;
    wire N__38810;
    wire N__38807;
    wire N__38806;
    wire N__38805;
    wire N__38802;
    wire N__38799;
    wire N__38796;
    wire N__38793;
    wire N__38786;
    wire N__38783;
    wire N__38782;
    wire N__38781;
    wire N__38778;
    wire N__38775;
    wire N__38772;
    wire N__38767;
    wire N__38762;
    wire N__38759;
    wire N__38758;
    wire N__38757;
    wire N__38754;
    wire N__38751;
    wire N__38748;
    wire N__38743;
    wire N__38738;
    wire N__38735;
    wire N__38734;
    wire N__38733;
    wire N__38730;
    wire N__38725;
    wire N__38720;
    wire N__38717;
    wire N__38716;
    wire N__38715;
    wire N__38712;
    wire N__38707;
    wire N__38702;
    wire N__38699;
    wire N__38698;
    wire N__38697;
    wire N__38694;
    wire N__38691;
    wire N__38688;
    wire N__38683;
    wire N__38678;
    wire N__38675;
    wire N__38674;
    wire N__38673;
    wire N__38670;
    wire N__38667;
    wire N__38664;
    wire N__38659;
    wire N__38654;
    wire N__38651;
    wire N__38650;
    wire N__38649;
    wire N__38646;
    wire N__38643;
    wire N__38640;
    wire N__38637;
    wire N__38630;
    wire N__38627;
    wire N__38626;
    wire N__38625;
    wire N__38622;
    wire N__38619;
    wire N__38616;
    wire N__38613;
    wire N__38606;
    wire N__38603;
    wire N__38602;
    wire N__38601;
    wire N__38598;
    wire N__38595;
    wire N__38592;
    wire N__38587;
    wire N__38582;
    wire N__38579;
    wire N__38578;
    wire N__38577;
    wire N__38574;
    wire N__38571;
    wire N__38568;
    wire N__38563;
    wire N__38558;
    wire N__38555;
    wire N__38554;
    wire N__38553;
    wire N__38550;
    wire N__38545;
    wire N__38540;
    wire N__38537;
    wire N__38536;
    wire N__38535;
    wire N__38532;
    wire N__38527;
    wire N__38522;
    wire N__38519;
    wire N__38516;
    wire N__38513;
    wire N__38510;
    wire N__38509;
    wire N__38506;
    wire N__38503;
    wire N__38500;
    wire N__38497;
    wire N__38494;
    wire N__38489;
    wire N__38486;
    wire N__38483;
    wire N__38480;
    wire N__38477;
    wire N__38476;
    wire N__38473;
    wire N__38470;
    wire N__38467;
    wire N__38464;
    wire N__38461;
    wire N__38456;
    wire N__38455;
    wire N__38454;
    wire N__38451;
    wire N__38448;
    wire N__38445;
    wire N__38438;
    wire N__38435;
    wire N__38434;
    wire N__38433;
    wire N__38430;
    wire N__38427;
    wire N__38424;
    wire N__38417;
    wire N__38414;
    wire N__38413;
    wire N__38412;
    wire N__38409;
    wire N__38406;
    wire N__38403;
    wire N__38398;
    wire N__38393;
    wire N__38390;
    wire N__38389;
    wire N__38388;
    wire N__38385;
    wire N__38382;
    wire N__38379;
    wire N__38374;
    wire N__38369;
    wire N__38366;
    wire N__38365;
    wire N__38364;
    wire N__38361;
    wire N__38356;
    wire N__38351;
    wire N__38348;
    wire N__38347;
    wire N__38346;
    wire N__38343;
    wire N__38338;
    wire N__38333;
    wire N__38330;
    wire N__38327;
    wire N__38324;
    wire N__38321;
    wire N__38320;
    wire N__38317;
    wire N__38314;
    wire N__38311;
    wire N__38306;
    wire N__38303;
    wire N__38300;
    wire N__38297;
    wire N__38294;
    wire N__38291;
    wire N__38288;
    wire N__38287;
    wire N__38286;
    wire N__38283;
    wire N__38280;
    wire N__38277;
    wire N__38274;
    wire N__38269;
    wire N__38264;
    wire N__38261;
    wire N__38258;
    wire N__38255;
    wire N__38252;
    wire N__38251;
    wire N__38248;
    wire N__38245;
    wire N__38242;
    wire N__38239;
    wire N__38234;
    wire N__38231;
    wire N__38228;
    wire N__38225;
    wire N__38222;
    wire N__38219;
    wire N__38218;
    wire N__38215;
    wire N__38212;
    wire N__38209;
    wire N__38204;
    wire N__38201;
    wire N__38198;
    wire N__38195;
    wire N__38194;
    wire N__38191;
    wire N__38188;
    wire N__38185;
    wire N__38180;
    wire N__38179;
    wire N__38178;
    wire N__38177;
    wire N__38176;
    wire N__38175;
    wire N__38174;
    wire N__38173;
    wire N__38170;
    wire N__38167;
    wire N__38166;
    wire N__38165;
    wire N__38164;
    wire N__38163;
    wire N__38162;
    wire N__38161;
    wire N__38160;
    wire N__38159;
    wire N__38148;
    wire N__38147;
    wire N__38146;
    wire N__38145;
    wire N__38144;
    wire N__38143;
    wire N__38142;
    wire N__38127;
    wire N__38118;
    wire N__38117;
    wire N__38114;
    wire N__38107;
    wire N__38104;
    wire N__38103;
    wire N__38098;
    wire N__38093;
    wire N__38090;
    wire N__38085;
    wire N__38080;
    wire N__38075;
    wire N__38072;
    wire N__38069;
    wire N__38064;
    wire N__38061;
    wire N__38058;
    wire N__38051;
    wire N__38050;
    wire N__38049;
    wire N__38048;
    wire N__38047;
    wire N__38046;
    wire N__38045;
    wire N__38044;
    wire N__38043;
    wire N__38040;
    wire N__38039;
    wire N__38038;
    wire N__38037;
    wire N__38034;
    wire N__38031;
    wire N__38028;
    wire N__38025;
    wire N__38024;
    wire N__38023;
    wire N__38022;
    wire N__38019;
    wire N__38018;
    wire N__38017;
    wire N__38016;
    wire N__38015;
    wire N__38012;
    wire N__38009;
    wire N__38006;
    wire N__38005;
    wire N__38004;
    wire N__37999;
    wire N__37998;
    wire N__37987;
    wire N__37982;
    wire N__37967;
    wire N__37964;
    wire N__37955;
    wire N__37952;
    wire N__37951;
    wire N__37948;
    wire N__37947;
    wire N__37944;
    wire N__37937;
    wire N__37934;
    wire N__37931;
    wire N__37924;
    wire N__37919;
    wire N__37910;
    wire N__37907;
    wire N__37904;
    wire N__37901;
    wire N__37900;
    wire N__37899;
    wire N__37898;
    wire N__37897;
    wire N__37896;
    wire N__37895;
    wire N__37894;
    wire N__37893;
    wire N__37892;
    wire N__37889;
    wire N__37886;
    wire N__37885;
    wire N__37884;
    wire N__37881;
    wire N__37878;
    wire N__37877;
    wire N__37876;
    wire N__37875;
    wire N__37874;
    wire N__37873;
    wire N__37862;
    wire N__37861;
    wire N__37860;
    wire N__37859;
    wire N__37858;
    wire N__37855;
    wire N__37850;
    wire N__37845;
    wire N__37830;
    wire N__37827;
    wire N__37826;
    wire N__37823;
    wire N__37818;
    wire N__37815;
    wire N__37812;
    wire N__37803;
    wire N__37800;
    wire N__37795;
    wire N__37794;
    wire N__37793;
    wire N__37786;
    wire N__37783;
    wire N__37780;
    wire N__37775;
    wire N__37770;
    wire N__37767;
    wire N__37760;
    wire N__37757;
    wire N__37756;
    wire N__37753;
    wire N__37750;
    wire N__37747;
    wire N__37742;
    wire N__37739;
    wire N__37736;
    wire N__37733;
    wire N__37732;
    wire N__37729;
    wire N__37726;
    wire N__37723;
    wire N__37720;
    wire N__37715;
    wire N__37712;
    wire N__37709;
    wire N__37706;
    wire N__37705;
    wire N__37702;
    wire N__37699;
    wire N__37696;
    wire N__37693;
    wire N__37690;
    wire N__37685;
    wire N__37682;
    wire N__37679;
    wire N__37676;
    wire N__37675;
    wire N__37672;
    wire N__37669;
    wire N__37666;
    wire N__37661;
    wire N__37658;
    wire N__37655;
    wire N__37652;
    wire N__37651;
    wire N__37648;
    wire N__37645;
    wire N__37642;
    wire N__37637;
    wire N__37634;
    wire N__37631;
    wire N__37628;
    wire N__37627;
    wire N__37624;
    wire N__37621;
    wire N__37618;
    wire N__37613;
    wire N__37610;
    wire N__37607;
    wire N__37604;
    wire N__37601;
    wire N__37598;
    wire N__37597;
    wire N__37594;
    wire N__37591;
    wire N__37588;
    wire N__37585;
    wire N__37580;
    wire N__37577;
    wire N__37574;
    wire N__37571;
    wire N__37568;
    wire N__37565;
    wire N__37564;
    wire N__37561;
    wire N__37558;
    wire N__37555;
    wire N__37552;
    wire N__37547;
    wire N__37544;
    wire N__37541;
    wire N__37538;
    wire N__37537;
    wire N__37534;
    wire N__37531;
    wire N__37528;
    wire N__37523;
    wire N__37520;
    wire N__37517;
    wire N__37514;
    wire N__37513;
    wire N__37510;
    wire N__37507;
    wire N__37504;
    wire N__37499;
    wire N__37496;
    wire N__37493;
    wire N__37490;
    wire N__37487;
    wire N__37486;
    wire N__37483;
    wire N__37480;
    wire N__37477;
    wire N__37474;
    wire N__37469;
    wire N__37466;
    wire N__37465;
    wire N__37464;
    wire N__37457;
    wire N__37456;
    wire N__37455;
    wire N__37454;
    wire N__37451;
    wire N__37444;
    wire N__37439;
    wire N__37438;
    wire N__37437;
    wire N__37434;
    wire N__37429;
    wire N__37424;
    wire N__37423;
    wire N__37422;
    wire N__37419;
    wire N__37414;
    wire N__37409;
    wire N__37406;
    wire N__37405;
    wire N__37402;
    wire N__37399;
    wire N__37398;
    wire N__37395;
    wire N__37390;
    wire N__37385;
    wire N__37382;
    wire N__37379;
    wire N__37378;
    wire N__37375;
    wire N__37372;
    wire N__37369;
    wire N__37364;
    wire N__37363;
    wire N__37362;
    wire N__37361;
    wire N__37354;
    wire N__37351;
    wire N__37350;
    wire N__37349;
    wire N__37346;
    wire N__37343;
    wire N__37338;
    wire N__37333;
    wire N__37328;
    wire N__37327;
    wire N__37326;
    wire N__37323;
    wire N__37320;
    wire N__37317;
    wire N__37314;
    wire N__37313;
    wire N__37310;
    wire N__37307;
    wire N__37304;
    wire N__37301;
    wire N__37296;
    wire N__37293;
    wire N__37290;
    wire N__37287;
    wire N__37280;
    wire N__37279;
    wire N__37278;
    wire N__37277;
    wire N__37276;
    wire N__37275;
    wire N__37264;
    wire N__37261;
    wire N__37260;
    wire N__37257;
    wire N__37256;
    wire N__37255;
    wire N__37254;
    wire N__37251;
    wire N__37248;
    wire N__37245;
    wire N__37238;
    wire N__37235;
    wire N__37226;
    wire N__37225;
    wire N__37224;
    wire N__37221;
    wire N__37218;
    wire N__37215;
    wire N__37212;
    wire N__37209;
    wire N__37206;
    wire N__37203;
    wire N__37202;
    wire N__37197;
    wire N__37194;
    wire N__37191;
    wire N__37188;
    wire N__37181;
    wire N__37178;
    wire N__37175;
    wire N__37174;
    wire N__37171;
    wire N__37168;
    wire N__37165;
    wire N__37160;
    wire N__37157;
    wire N__37154;
    wire N__37151;
    wire N__37150;
    wire N__37147;
    wire N__37144;
    wire N__37141;
    wire N__37136;
    wire N__37133;
    wire N__37130;
    wire N__37127;
    wire N__37126;
    wire N__37123;
    wire N__37120;
    wire N__37117;
    wire N__37112;
    wire N__37109;
    wire N__37106;
    wire N__37103;
    wire N__37100;
    wire N__37099;
    wire N__37096;
    wire N__37093;
    wire N__37090;
    wire N__37085;
    wire N__37082;
    wire N__37079;
    wire N__37076;
    wire N__37075;
    wire N__37072;
    wire N__37069;
    wire N__37066;
    wire N__37063;
    wire N__37062;
    wire N__37059;
    wire N__37056;
    wire N__37053;
    wire N__37046;
    wire N__37043;
    wire N__37040;
    wire N__37037;
    wire N__37034;
    wire N__37031;
    wire N__37028;
    wire N__37025;
    wire N__37022;
    wire N__37019;
    wire N__37016;
    wire N__37013;
    wire N__37010;
    wire N__37007;
    wire N__37004;
    wire N__37001;
    wire N__36998;
    wire N__36995;
    wire N__36992;
    wire N__36989;
    wire N__36986;
    wire N__36983;
    wire N__36980;
    wire N__36977;
    wire N__36974;
    wire N__36971;
    wire N__36968;
    wire N__36965;
    wire N__36962;
    wire N__36961;
    wire N__36958;
    wire N__36955;
    wire N__36952;
    wire N__36947;
    wire N__36944;
    wire N__36941;
    wire N__36938;
    wire N__36935;
    wire N__36934;
    wire N__36931;
    wire N__36928;
    wire N__36925;
    wire N__36920;
    wire N__36917;
    wire N__36914;
    wire N__36911;
    wire N__36908;
    wire N__36905;
    wire N__36902;
    wire N__36899;
    wire N__36896;
    wire N__36895;
    wire N__36892;
    wire N__36889;
    wire N__36886;
    wire N__36881;
    wire N__36878;
    wire N__36875;
    wire N__36872;
    wire N__36869;
    wire N__36866;
    wire N__36863;
    wire N__36860;
    wire N__36857;
    wire N__36854;
    wire N__36851;
    wire N__36848;
    wire N__36845;
    wire N__36842;
    wire N__36839;
    wire N__36836;
    wire N__36833;
    wire N__36830;
    wire N__36827;
    wire N__36826;
    wire N__36823;
    wire N__36820;
    wire N__36817;
    wire N__36814;
    wire N__36809;
    wire N__36806;
    wire N__36803;
    wire N__36800;
    wire N__36797;
    wire N__36794;
    wire N__36791;
    wire N__36788;
    wire N__36785;
    wire N__36782;
    wire N__36779;
    wire N__36776;
    wire N__36773;
    wire N__36770;
    wire N__36767;
    wire N__36764;
    wire N__36761;
    wire N__36758;
    wire N__36755;
    wire N__36752;
    wire N__36749;
    wire N__36746;
    wire N__36743;
    wire N__36742;
    wire N__36739;
    wire N__36736;
    wire N__36731;
    wire N__36728;
    wire N__36725;
    wire N__36722;
    wire N__36719;
    wire N__36718;
    wire N__36715;
    wire N__36712;
    wire N__36707;
    wire N__36704;
    wire N__36701;
    wire N__36700;
    wire N__36697;
    wire N__36694;
    wire N__36693;
    wire N__36688;
    wire N__36685;
    wire N__36682;
    wire N__36677;
    wire N__36674;
    wire N__36673;
    wire N__36670;
    wire N__36669;
    wire N__36666;
    wire N__36663;
    wire N__36660;
    wire N__36655;
    wire N__36650;
    wire N__36647;
    wire N__36646;
    wire N__36643;
    wire N__36642;
    wire N__36639;
    wire N__36636;
    wire N__36633;
    wire N__36628;
    wire N__36623;
    wire N__36620;
    wire N__36619;
    wire N__36616;
    wire N__36613;
    wire N__36612;
    wire N__36607;
    wire N__36604;
    wire N__36601;
    wire N__36596;
    wire N__36593;
    wire N__36592;
    wire N__36589;
    wire N__36586;
    wire N__36585;
    wire N__36580;
    wire N__36577;
    wire N__36574;
    wire N__36569;
    wire N__36566;
    wire N__36565;
    wire N__36562;
    wire N__36559;
    wire N__36556;
    wire N__36551;
    wire N__36548;
    wire N__36547;
    wire N__36546;
    wire N__36545;
    wire N__36544;
    wire N__36543;
    wire N__36542;
    wire N__36541;
    wire N__36540;
    wire N__36539;
    wire N__36538;
    wire N__36537;
    wire N__36536;
    wire N__36535;
    wire N__36534;
    wire N__36533;
    wire N__36532;
    wire N__36531;
    wire N__36530;
    wire N__36529;
    wire N__36528;
    wire N__36527;
    wire N__36526;
    wire N__36525;
    wire N__36524;
    wire N__36523;
    wire N__36522;
    wire N__36521;
    wire N__36520;
    wire N__36519;
    wire N__36510;
    wire N__36501;
    wire N__36492;
    wire N__36483;
    wire N__36478;
    wire N__36469;
    wire N__36460;
    wire N__36451;
    wire N__36448;
    wire N__36433;
    wire N__36428;
    wire N__36425;
    wire N__36424;
    wire N__36421;
    wire N__36418;
    wire N__36415;
    wire N__36410;
    wire N__36409;
    wire N__36408;
    wire N__36407;
    wire N__36404;
    wire N__36401;
    wire N__36398;
    wire N__36395;
    wire N__36390;
    wire N__36385;
    wire N__36382;
    wire N__36377;
    wire N__36374;
    wire N__36371;
    wire N__36368;
    wire N__36365;
    wire N__36364;
    wire N__36361;
    wire N__36358;
    wire N__36357;
    wire N__36352;
    wire N__36349;
    wire N__36346;
    wire N__36341;
    wire N__36338;
    wire N__36337;
    wire N__36334;
    wire N__36331;
    wire N__36330;
    wire N__36325;
    wire N__36322;
    wire N__36319;
    wire N__36314;
    wire N__36311;
    wire N__36310;
    wire N__36307;
    wire N__36304;
    wire N__36303;
    wire N__36300;
    wire N__36297;
    wire N__36294;
    wire N__36289;
    wire N__36284;
    wire N__36281;
    wire N__36280;
    wire N__36277;
    wire N__36276;
    wire N__36273;
    wire N__36270;
    wire N__36267;
    wire N__36262;
    wire N__36257;
    wire N__36254;
    wire N__36253;
    wire N__36250;
    wire N__36247;
    wire N__36246;
    wire N__36241;
    wire N__36238;
    wire N__36235;
    wire N__36230;
    wire N__36227;
    wire N__36226;
    wire N__36223;
    wire N__36220;
    wire N__36219;
    wire N__36214;
    wire N__36211;
    wire N__36208;
    wire N__36203;
    wire N__36200;
    wire N__36199;
    wire N__36198;
    wire N__36193;
    wire N__36190;
    wire N__36187;
    wire N__36182;
    wire N__36179;
    wire N__36178;
    wire N__36177;
    wire N__36172;
    wire N__36169;
    wire N__36166;
    wire N__36161;
    wire N__36158;
    wire N__36157;
    wire N__36154;
    wire N__36151;
    wire N__36150;
    wire N__36145;
    wire N__36142;
    wire N__36139;
    wire N__36134;
    wire N__36131;
    wire N__36130;
    wire N__36129;
    wire N__36124;
    wire N__36121;
    wire N__36118;
    wire N__36113;
    wire N__36110;
    wire N__36109;
    wire N__36108;
    wire N__36103;
    wire N__36100;
    wire N__36097;
    wire N__36092;
    wire N__36089;
    wire N__36086;
    wire N__36083;
    wire N__36082;
    wire N__36079;
    wire N__36078;
    wire N__36075;
    wire N__36072;
    wire N__36069;
    wire N__36064;
    wire N__36059;
    wire N__36056;
    wire N__36055;
    wire N__36052;
    wire N__36049;
    wire N__36046;
    wire N__36045;
    wire N__36040;
    wire N__36037;
    wire N__36034;
    wire N__36029;
    wire N__36026;
    wire N__36025;
    wire N__36022;
    wire N__36019;
    wire N__36018;
    wire N__36013;
    wire N__36010;
    wire N__36007;
    wire N__36002;
    wire N__35999;
    wire N__35998;
    wire N__35995;
    wire N__35992;
    wire N__35991;
    wire N__35986;
    wire N__35983;
    wire N__35980;
    wire N__35975;
    wire N__35972;
    wire N__35971;
    wire N__35970;
    wire N__35965;
    wire N__35962;
    wire N__35959;
    wire N__35954;
    wire N__35951;
    wire N__35950;
    wire N__35949;
    wire N__35944;
    wire N__35941;
    wire N__35938;
    wire N__35933;
    wire N__35930;
    wire N__35929;
    wire N__35926;
    wire N__35923;
    wire N__35920;
    wire N__35917;
    wire N__35916;
    wire N__35911;
    wire N__35908;
    wire N__35903;
    wire N__35900;
    wire N__35899;
    wire N__35896;
    wire N__35893;
    wire N__35888;
    wire N__35885;
    wire N__35882;
    wire N__35881;
    wire N__35878;
    wire N__35875;
    wire N__35872;
    wire N__35869;
    wire N__35868;
    wire N__35863;
    wire N__35860;
    wire N__35855;
    wire N__35854;
    wire N__35851;
    wire N__35850;
    wire N__35847;
    wire N__35844;
    wire N__35841;
    wire N__35836;
    wire N__35831;
    wire N__35828;
    wire N__35827;
    wire N__35824;
    wire N__35821;
    wire N__35820;
    wire N__35817;
    wire N__35814;
    wire N__35811;
    wire N__35808;
    wire N__35801;
    wire N__35798;
    wire N__35797;
    wire N__35796;
    wire N__35791;
    wire N__35788;
    wire N__35785;
    wire N__35780;
    wire N__35777;
    wire N__35776;
    wire N__35775;
    wire N__35770;
    wire N__35767;
    wire N__35764;
    wire N__35759;
    wire N__35756;
    wire N__35755;
    wire N__35752;
    wire N__35749;
    wire N__35744;
    wire N__35743;
    wire N__35740;
    wire N__35737;
    wire N__35734;
    wire N__35729;
    wire N__35726;
    wire N__35725;
    wire N__35722;
    wire N__35719;
    wire N__35718;
    wire N__35713;
    wire N__35710;
    wire N__35707;
    wire N__35702;
    wire N__35699;
    wire N__35698;
    wire N__35697;
    wire N__35696;
    wire N__35695;
    wire N__35684;
    wire N__35681;
    wire N__35678;
    wire N__35677;
    wire N__35674;
    wire N__35671;
    wire N__35670;
    wire N__35667;
    wire N__35664;
    wire N__35661;
    wire N__35658;
    wire N__35657;
    wire N__35656;
    wire N__35651;
    wire N__35648;
    wire N__35645;
    wire N__35642;
    wire N__35633;
    wire N__35630;
    wire N__35627;
    wire N__35624;
    wire N__35621;
    wire N__35618;
    wire N__35615;
    wire N__35612;
    wire N__35609;
    wire N__35606;
    wire N__35603;
    wire N__35600;
    wire N__35597;
    wire N__35594;
    wire N__35593;
    wire N__35592;
    wire N__35589;
    wire N__35584;
    wire N__35579;
    wire N__35576;
    wire N__35573;
    wire N__35570;
    wire N__35569;
    wire N__35566;
    wire N__35563;
    wire N__35560;
    wire N__35559;
    wire N__35558;
    wire N__35553;
    wire N__35548;
    wire N__35543;
    wire N__35540;
    wire N__35539;
    wire N__35538;
    wire N__35535;
    wire N__35532;
    wire N__35529;
    wire N__35522;
    wire N__35519;
    wire N__35518;
    wire N__35517;
    wire N__35514;
    wire N__35513;
    wire N__35510;
    wire N__35507;
    wire N__35504;
    wire N__35501;
    wire N__35500;
    wire N__35497;
    wire N__35494;
    wire N__35491;
    wire N__35488;
    wire N__35485;
    wire N__35482;
    wire N__35479;
    wire N__35474;
    wire N__35471;
    wire N__35468;
    wire N__35465;
    wire N__35462;
    wire N__35453;
    wire N__35450;
    wire N__35449;
    wire N__35448;
    wire N__35445;
    wire N__35442;
    wire N__35439;
    wire N__35432;
    wire N__35431;
    wire N__35428;
    wire N__35427;
    wire N__35426;
    wire N__35423;
    wire N__35422;
    wire N__35419;
    wire N__35416;
    wire N__35413;
    wire N__35410;
    wire N__35407;
    wire N__35404;
    wire N__35401;
    wire N__35398;
    wire N__35395;
    wire N__35392;
    wire N__35389;
    wire N__35386;
    wire N__35383;
    wire N__35380;
    wire N__35369;
    wire N__35366;
    wire N__35363;
    wire N__35360;
    wire N__35357;
    wire N__35354;
    wire N__35351;
    wire N__35348;
    wire N__35345;
    wire N__35342;
    wire N__35339;
    wire N__35336;
    wire N__35333;
    wire N__35330;
    wire N__35327;
    wire N__35324;
    wire N__35321;
    wire N__35318;
    wire N__35315;
    wire N__35314;
    wire N__35313;
    wire N__35306;
    wire N__35303;
    wire N__35302;
    wire N__35299;
    wire N__35298;
    wire N__35295;
    wire N__35292;
    wire N__35289;
    wire N__35288;
    wire N__35285;
    wire N__35280;
    wire N__35277;
    wire N__35270;
    wire N__35267;
    wire N__35264;
    wire N__35261;
    wire N__35260;
    wire N__35259;
    wire N__35258;
    wire N__35257;
    wire N__35256;
    wire N__35253;
    wire N__35250;
    wire N__35249;
    wire N__35246;
    wire N__35243;
    wire N__35240;
    wire N__35237;
    wire N__35232;
    wire N__35229;
    wire N__35224;
    wire N__35213;
    wire N__35210;
    wire N__35207;
    wire N__35206;
    wire N__35203;
    wire N__35200;
    wire N__35195;
    wire N__35194;
    wire N__35191;
    wire N__35188;
    wire N__35183;
    wire N__35180;
    wire N__35177;
    wire N__35174;
    wire N__35171;
    wire N__35170;
    wire N__35167;
    wire N__35162;
    wire N__35159;
    wire N__35156;
    wire N__35155;
    wire N__35150;
    wire N__35147;
    wire N__35144;
    wire N__35143;
    wire N__35140;
    wire N__35137;
    wire N__35132;
    wire N__35129;
    wire N__35128;
    wire N__35125;
    wire N__35124;
    wire N__35121;
    wire N__35118;
    wire N__35117;
    wire N__35114;
    wire N__35111;
    wire N__35108;
    wire N__35105;
    wire N__35102;
    wire N__35099;
    wire N__35090;
    wire N__35087;
    wire N__35084;
    wire N__35081;
    wire N__35080;
    wire N__35077;
    wire N__35076;
    wire N__35075;
    wire N__35072;
    wire N__35069;
    wire N__35066;
    wire N__35063;
    wire N__35060;
    wire N__35057;
    wire N__35054;
    wire N__35049;
    wire N__35042;
    wire N__35039;
    wire N__35038;
    wire N__35035;
    wire N__35032;
    wire N__35031;
    wire N__35028;
    wire N__35025;
    wire N__35022;
    wire N__35015;
    wire N__35012;
    wire N__35011;
    wire N__35008;
    wire N__35003;
    wire N__35002;
    wire N__34999;
    wire N__34996;
    wire N__34991;
    wire N__34988;
    wire N__34985;
    wire N__34984;
    wire N__34983;
    wire N__34978;
    wire N__34975;
    wire N__34972;
    wire N__34969;
    wire N__34964;
    wire N__34961;
    wire N__34960;
    wire N__34957;
    wire N__34954;
    wire N__34951;
    wire N__34948;
    wire N__34947;
    wire N__34944;
    wire N__34941;
    wire N__34938;
    wire N__34935;
    wire N__34928;
    wire N__34925;
    wire N__34922;
    wire N__34919;
    wire N__34916;
    wire N__34913;
    wire N__34910;
    wire N__34907;
    wire N__34906;
    wire N__34905;
    wire N__34904;
    wire N__34901;
    wire N__34894;
    wire N__34891;
    wire N__34888;
    wire N__34885;
    wire N__34882;
    wire N__34879;
    wire N__34876;
    wire N__34871;
    wire N__34868;
    wire N__34865;
    wire N__34862;
    wire N__34859;
    wire N__34858;
    wire N__34855;
    wire N__34852;
    wire N__34847;
    wire N__34844;
    wire N__34841;
    wire N__34840;
    wire N__34839;
    wire N__34836;
    wire N__34833;
    wire N__34830;
    wire N__34823;
    wire N__34820;
    wire N__34817;
    wire N__34814;
    wire N__34813;
    wire N__34810;
    wire N__34807;
    wire N__34804;
    wire N__34803;
    wire N__34800;
    wire N__34797;
    wire N__34794;
    wire N__34791;
    wire N__34784;
    wire N__34781;
    wire N__34778;
    wire N__34775;
    wire N__34772;
    wire N__34769;
    wire N__34766;
    wire N__34763;
    wire N__34760;
    wire N__34757;
    wire N__34754;
    wire N__34751;
    wire N__34748;
    wire N__34745;
    wire N__34742;
    wire N__34739;
    wire N__34736;
    wire N__34733;
    wire N__34730;
    wire N__34727;
    wire N__34726;
    wire N__34723;
    wire N__34720;
    wire N__34715;
    wire N__34712;
    wire N__34709;
    wire N__34706;
    wire N__34703;
    wire N__34700;
    wire N__34699;
    wire N__34696;
    wire N__34693;
    wire N__34688;
    wire N__34685;
    wire N__34682;
    wire N__34679;
    wire N__34676;
    wire N__34673;
    wire N__34670;
    wire N__34667;
    wire N__34666;
    wire N__34663;
    wire N__34660;
    wire N__34655;
    wire N__34652;
    wire N__34649;
    wire N__34646;
    wire N__34643;
    wire N__34640;
    wire N__34637;
    wire N__34636;
    wire N__34633;
    wire N__34630;
    wire N__34627;
    wire N__34624;
    wire N__34619;
    wire N__34616;
    wire N__34613;
    wire N__34610;
    wire N__34607;
    wire N__34606;
    wire N__34603;
    wire N__34600;
    wire N__34597;
    wire N__34592;
    wire N__34589;
    wire N__34586;
    wire N__34583;
    wire N__34580;
    wire N__34577;
    wire N__34574;
    wire N__34571;
    wire N__34568;
    wire N__34565;
    wire N__34564;
    wire N__34561;
    wire N__34558;
    wire N__34557;
    wire N__34552;
    wire N__34549;
    wire N__34546;
    wire N__34545;
    wire N__34544;
    wire N__34541;
    wire N__34538;
    wire N__34537;
    wire N__34536;
    wire N__34531;
    wire N__34528;
    wire N__34525;
    wire N__34522;
    wire N__34519;
    wire N__34516;
    wire N__34513;
    wire N__34510;
    wire N__34507;
    wire N__34504;
    wire N__34501;
    wire N__34498;
    wire N__34491;
    wire N__34488;
    wire N__34483;
    wire N__34480;
    wire N__34475;
    wire N__34474;
    wire N__34471;
    wire N__34468;
    wire N__34465;
    wire N__34462;
    wire N__34459;
    wire N__34454;
    wire N__34453;
    wire N__34448;
    wire N__34445;
    wire N__34442;
    wire N__34439;
    wire N__34436;
    wire N__34433;
    wire N__34432;
    wire N__34431;
    wire N__34428;
    wire N__34423;
    wire N__34418;
    wire N__34417;
    wire N__34412;
    wire N__34411;
    wire N__34410;
    wire N__34407;
    wire N__34404;
    wire N__34403;
    wire N__34402;
    wire N__34399;
    wire N__34396;
    wire N__34393;
    wire N__34388;
    wire N__34379;
    wire N__34376;
    wire N__34373;
    wire N__34370;
    wire N__34369;
    wire N__34366;
    wire N__34365;
    wire N__34362;
    wire N__34359;
    wire N__34356;
    wire N__34349;
    wire N__34346;
    wire N__34345;
    wire N__34342;
    wire N__34339;
    wire N__34334;
    wire N__34331;
    wire N__34328;
    wire N__34325;
    wire N__34322;
    wire N__34319;
    wire N__34316;
    wire N__34313;
    wire N__34310;
    wire N__34309;
    wire N__34306;
    wire N__34303;
    wire N__34298;
    wire N__34295;
    wire N__34292;
    wire N__34289;
    wire N__34286;
    wire N__34283;
    wire N__34280;
    wire N__34279;
    wire N__34276;
    wire N__34273;
    wire N__34268;
    wire N__34265;
    wire N__34262;
    wire N__34259;
    wire N__34256;
    wire N__34253;
    wire N__34250;
    wire N__34249;
    wire N__34246;
    wire N__34243;
    wire N__34238;
    wire N__34235;
    wire N__34232;
    wire N__34229;
    wire N__34226;
    wire N__34223;
    wire N__34220;
    wire N__34217;
    wire N__34214;
    wire N__34211;
    wire N__34208;
    wire N__34205;
    wire N__34202;
    wire N__34199;
    wire N__34196;
    wire N__34193;
    wire N__34190;
    wire N__34187;
    wire N__34184;
    wire N__34181;
    wire N__34178;
    wire N__34175;
    wire N__34172;
    wire N__34169;
    wire N__34166;
    wire N__34165;
    wire N__34162;
    wire N__34159;
    wire N__34158;
    wire N__34155;
    wire N__34152;
    wire N__34151;
    wire N__34150;
    wire N__34147;
    wire N__34144;
    wire N__34141;
    wire N__34138;
    wire N__34135;
    wire N__34132;
    wire N__34125;
    wire N__34122;
    wire N__34115;
    wire N__34114;
    wire N__34111;
    wire N__34108;
    wire N__34107;
    wire N__34106;
    wire N__34103;
    wire N__34100;
    wire N__34099;
    wire N__34096;
    wire N__34093;
    wire N__34090;
    wire N__34087;
    wire N__34084;
    wire N__34081;
    wire N__34078;
    wire N__34075;
    wire N__34072;
    wire N__34069;
    wire N__34066;
    wire N__34055;
    wire N__34052;
    wire N__34049;
    wire N__34048;
    wire N__34047;
    wire N__34046;
    wire N__34043;
    wire N__34040;
    wire N__34037;
    wire N__34034;
    wire N__34031;
    wire N__34030;
    wire N__34029;
    wire N__34024;
    wire N__34021;
    wire N__34018;
    wire N__34015;
    wire N__34012;
    wire N__34009;
    wire N__33998;
    wire N__33995;
    wire N__33992;
    wire N__33989;
    wire N__33986;
    wire N__33983;
    wire N__33980;
    wire N__33977;
    wire N__33974;
    wire N__33971;
    wire N__33968;
    wire N__33965;
    wire N__33962;
    wire N__33959;
    wire N__33956;
    wire N__33953;
    wire N__33950;
    wire N__33947;
    wire N__33944;
    wire N__33941;
    wire N__33938;
    wire N__33935;
    wire N__33932;
    wire N__33929;
    wire N__33926;
    wire N__33923;
    wire N__33920;
    wire N__33917;
    wire N__33916;
    wire N__33913;
    wire N__33910;
    wire N__33907;
    wire N__33904;
    wire N__33903;
    wire N__33902;
    wire N__33901;
    wire N__33898;
    wire N__33895;
    wire N__33892;
    wire N__33887;
    wire N__33878;
    wire N__33877;
    wire N__33876;
    wire N__33873;
    wire N__33870;
    wire N__33867;
    wire N__33866;
    wire N__33863;
    wire N__33860;
    wire N__33857;
    wire N__33854;
    wire N__33853;
    wire N__33850;
    wire N__33845;
    wire N__33840;
    wire N__33833;
    wire N__33832;
    wire N__33827;
    wire N__33826;
    wire N__33823;
    wire N__33820;
    wire N__33817;
    wire N__33812;
    wire N__33809;
    wire N__33806;
    wire N__33805;
    wire N__33804;
    wire N__33801;
    wire N__33796;
    wire N__33791;
    wire N__33788;
    wire N__33787;
    wire N__33784;
    wire N__33783;
    wire N__33780;
    wire N__33777;
    wire N__33774;
    wire N__33773;
    wire N__33770;
    wire N__33767;
    wire N__33762;
    wire N__33755;
    wire N__33752;
    wire N__33749;
    wire N__33746;
    wire N__33743;
    wire N__33740;
    wire N__33737;
    wire N__33734;
    wire N__33731;
    wire N__33728;
    wire N__33725;
    wire N__33722;
    wire N__33719;
    wire N__33716;
    wire N__33713;
    wire N__33712;
    wire N__33711;
    wire N__33704;
    wire N__33701;
    wire N__33698;
    wire N__33695;
    wire N__33692;
    wire N__33691;
    wire N__33688;
    wire N__33685;
    wire N__33680;
    wire N__33677;
    wire N__33674;
    wire N__33671;
    wire N__33668;
    wire N__33665;
    wire N__33662;
    wire N__33659;
    wire N__33656;
    wire N__33653;
    wire N__33650;
    wire N__33647;
    wire N__33646;
    wire N__33641;
    wire N__33638;
    wire N__33635;
    wire N__33632;
    wire N__33629;
    wire N__33628;
    wire N__33623;
    wire N__33620;
    wire N__33617;
    wire N__33614;
    wire N__33611;
    wire N__33608;
    wire N__33605;
    wire N__33602;
    wire N__33599;
    wire N__33596;
    wire N__33593;
    wire N__33592;
    wire N__33591;
    wire N__33586;
    wire N__33585;
    wire N__33582;
    wire N__33579;
    wire N__33576;
    wire N__33569;
    wire N__33566;
    wire N__33563;
    wire N__33560;
    wire N__33557;
    wire N__33554;
    wire N__33553;
    wire N__33550;
    wire N__33547;
    wire N__33542;
    wire N__33541;
    wire N__33538;
    wire N__33535;
    wire N__33530;
    wire N__33529;
    wire N__33526;
    wire N__33523;
    wire N__33520;
    wire N__33515;
    wire N__33514;
    wire N__33513;
    wire N__33512;
    wire N__33509;
    wire N__33506;
    wire N__33503;
    wire N__33500;
    wire N__33491;
    wire N__33490;
    wire N__33489;
    wire N__33486;
    wire N__33483;
    wire N__33482;
    wire N__33479;
    wire N__33476;
    wire N__33473;
    wire N__33470;
    wire N__33463;
    wire N__33460;
    wire N__33457;
    wire N__33452;
    wire N__33449;
    wire N__33446;
    wire N__33443;
    wire N__33440;
    wire N__33437;
    wire N__33434;
    wire N__33431;
    wire N__33428;
    wire N__33427;
    wire N__33426;
    wire N__33423;
    wire N__33420;
    wire N__33417;
    wire N__33412;
    wire N__33409;
    wire N__33404;
    wire N__33401;
    wire N__33398;
    wire N__33395;
    wire N__33392;
    wire N__33389;
    wire N__33386;
    wire N__33383;
    wire N__33380;
    wire N__33377;
    wire N__33374;
    wire N__33371;
    wire N__33368;
    wire N__33365;
    wire N__33362;
    wire N__33359;
    wire N__33356;
    wire N__33353;
    wire N__33350;
    wire N__33347;
    wire N__33344;
    wire N__33341;
    wire N__33338;
    wire N__33335;
    wire N__33332;
    wire N__33329;
    wire N__33326;
    wire N__33323;
    wire N__33320;
    wire N__33317;
    wire N__33314;
    wire N__33311;
    wire N__33308;
    wire N__33305;
    wire N__33304;
    wire N__33303;
    wire N__33298;
    wire N__33295;
    wire N__33290;
    wire N__33289;
    wire N__33288;
    wire N__33287;
    wire N__33284;
    wire N__33281;
    wire N__33278;
    wire N__33273;
    wire N__33266;
    wire N__33263;
    wire N__33260;
    wire N__33257;
    wire N__33254;
    wire N__33251;
    wire N__33248;
    wire N__33247;
    wire N__33244;
    wire N__33243;
    wire N__33242;
    wire N__33239;
    wire N__33236;
    wire N__33231;
    wire N__33224;
    wire N__33221;
    wire N__33218;
    wire N__33215;
    wire N__33212;
    wire N__33209;
    wire N__33206;
    wire N__33203;
    wire N__33200;
    wire N__33197;
    wire N__33194;
    wire N__33191;
    wire N__33188;
    wire N__33185;
    wire N__33182;
    wire N__33179;
    wire N__33176;
    wire N__33173;
    wire N__33170;
    wire N__33167;
    wire N__33164;
    wire N__33161;
    wire N__33158;
    wire N__33155;
    wire N__33152;
    wire N__33149;
    wire N__33146;
    wire N__33143;
    wire N__33140;
    wire N__33137;
    wire N__33134;
    wire N__33131;
    wire N__33128;
    wire N__33125;
    wire N__33122;
    wire N__33119;
    wire N__33116;
    wire N__33113;
    wire N__33110;
    wire N__33107;
    wire N__33104;
    wire N__33101;
    wire N__33098;
    wire N__33095;
    wire N__33092;
    wire N__33089;
    wire N__33086;
    wire N__33083;
    wire N__33080;
    wire N__33077;
    wire N__33074;
    wire N__33071;
    wire N__33068;
    wire N__33065;
    wire N__33062;
    wire N__33059;
    wire N__33056;
    wire N__33053;
    wire N__33050;
    wire N__33047;
    wire N__33044;
    wire N__33041;
    wire N__33038;
    wire N__33035;
    wire N__33032;
    wire N__33029;
    wire N__33026;
    wire N__33023;
    wire N__33020;
    wire N__33017;
    wire N__33014;
    wire N__33011;
    wire N__33008;
    wire N__33005;
    wire N__33002;
    wire N__32999;
    wire N__32996;
    wire N__32993;
    wire N__32990;
    wire N__32987;
    wire N__32984;
    wire N__32981;
    wire N__32978;
    wire N__32975;
    wire N__32972;
    wire N__32969;
    wire N__32966;
    wire N__32963;
    wire N__32960;
    wire N__32957;
    wire N__32954;
    wire N__32951;
    wire N__32948;
    wire N__32945;
    wire N__32942;
    wire N__32939;
    wire N__32936;
    wire N__32933;
    wire N__32930;
    wire N__32927;
    wire N__32924;
    wire N__32921;
    wire N__32918;
    wire N__32915;
    wire N__32912;
    wire N__32909;
    wire N__32906;
    wire N__32903;
    wire N__32900;
    wire N__32897;
    wire N__32894;
    wire N__32891;
    wire N__32888;
    wire N__32885;
    wire N__32882;
    wire N__32879;
    wire N__32876;
    wire N__32875;
    wire N__32872;
    wire N__32869;
    wire N__32866;
    wire N__32863;
    wire N__32858;
    wire N__32855;
    wire N__32852;
    wire N__32849;
    wire N__32846;
    wire N__32843;
    wire N__32842;
    wire N__32839;
    wire N__32838;
    wire N__32835;
    wire N__32832;
    wire N__32827;
    wire N__32822;
    wire N__32819;
    wire N__32816;
    wire N__32815;
    wire N__32810;
    wire N__32807;
    wire N__32804;
    wire N__32801;
    wire N__32798;
    wire N__32795;
    wire N__32794;
    wire N__32789;
    wire N__32786;
    wire N__32783;
    wire N__32780;
    wire N__32777;
    wire N__32774;
    wire N__32771;
    wire N__32768;
    wire N__32765;
    wire N__32762;
    wire N__32759;
    wire N__32756;
    wire N__32753;
    wire N__32750;
    wire N__32747;
    wire N__32744;
    wire N__32741;
    wire N__32740;
    wire N__32739;
    wire N__32738;
    wire N__32737;
    wire N__32726;
    wire N__32723;
    wire N__32720;
    wire N__32717;
    wire N__32716;
    wire N__32711;
    wire N__32708;
    wire N__32705;
    wire N__32702;
    wire N__32701;
    wire N__32700;
    wire N__32699;
    wire N__32698;
    wire N__32697;
    wire N__32696;
    wire N__32691;
    wire N__32680;
    wire N__32675;
    wire N__32672;
    wire N__32669;
    wire N__32666;
    wire N__32663;
    wire N__32660;
    wire N__32657;
    wire N__32654;
    wire N__32651;
    wire N__32648;
    wire N__32645;
    wire N__32642;
    wire N__32639;
    wire N__32636;
    wire N__32633;
    wire N__32630;
    wire N__32627;
    wire N__32624;
    wire N__32621;
    wire N__32618;
    wire N__32615;
    wire N__32612;
    wire N__32609;
    wire N__32606;
    wire N__32603;
    wire N__32600;
    wire N__32597;
    wire N__32594;
    wire N__32591;
    wire N__32588;
    wire N__32585;
    wire N__32582;
    wire N__32579;
    wire N__32576;
    wire N__32573;
    wire N__32570;
    wire N__32567;
    wire N__32564;
    wire N__32561;
    wire N__32558;
    wire N__32555;
    wire N__32552;
    wire N__32549;
    wire N__32546;
    wire N__32543;
    wire N__32540;
    wire N__32539;
    wire N__32538;
    wire N__32535;
    wire N__32532;
    wire N__32529;
    wire N__32526;
    wire N__32521;
    wire N__32518;
    wire N__32515;
    wire N__32510;
    wire N__32507;
    wire N__32506;
    wire N__32505;
    wire N__32504;
    wire N__32499;
    wire N__32496;
    wire N__32493;
    wire N__32486;
    wire N__32483;
    wire N__32480;
    wire N__32477;
    wire N__32474;
    wire N__32471;
    wire N__32468;
    wire N__32465;
    wire N__32462;
    wire N__32459;
    wire N__32456;
    wire N__32453;
    wire N__32450;
    wire N__32447;
    wire N__32444;
    wire N__32441;
    wire N__32438;
    wire N__32435;
    wire N__32432;
    wire N__32429;
    wire N__32426;
    wire N__32423;
    wire N__32420;
    wire N__32417;
    wire N__32414;
    wire N__32411;
    wire N__32408;
    wire N__32405;
    wire N__32402;
    wire N__32399;
    wire N__32396;
    wire N__32393;
    wire N__32392;
    wire N__32389;
    wire N__32386;
    wire N__32385;
    wire N__32382;
    wire N__32381;
    wire N__32380;
    wire N__32375;
    wire N__32372;
    wire N__32367;
    wire N__32362;
    wire N__32357;
    wire N__32356;
    wire N__32353;
    wire N__32352;
    wire N__32351;
    wire N__32350;
    wire N__32347;
    wire N__32342;
    wire N__32335;
    wire N__32330;
    wire N__32329;
    wire N__32328;
    wire N__32327;
    wire N__32324;
    wire N__32321;
    wire N__32316;
    wire N__32309;
    wire N__32308;
    wire N__32307;
    wire N__32306;
    wire N__32305;
    wire N__32304;
    wire N__32301;
    wire N__32300;
    wire N__32293;
    wire N__32288;
    wire N__32283;
    wire N__32276;
    wire N__32273;
    wire N__32270;
    wire N__32267;
    wire N__32264;
    wire N__32261;
    wire N__32258;
    wire N__32255;
    wire N__32252;
    wire N__32251;
    wire N__32250;
    wire N__32247;
    wire N__32246;
    wire N__32243;
    wire N__32240;
    wire N__32237;
    wire N__32234;
    wire N__32231;
    wire N__32228;
    wire N__32219;
    wire N__32218;
    wire N__32217;
    wire N__32214;
    wire N__32211;
    wire N__32208;
    wire N__32203;
    wire N__32200;
    wire N__32197;
    wire N__32194;
    wire N__32191;
    wire N__32188;
    wire N__32185;
    wire N__32182;
    wire N__32179;
    wire N__32176;
    wire N__32171;
    wire N__32168;
    wire N__32167;
    wire N__32166;
    wire N__32163;
    wire N__32158;
    wire N__32153;
    wire N__32152;
    wire N__32151;
    wire N__32150;
    wire N__32145;
    wire N__32140;
    wire N__32135;
    wire N__32134;
    wire N__32133;
    wire N__32130;
    wire N__32127;
    wire N__32126;
    wire N__32123;
    wire N__32120;
    wire N__32117;
    wire N__32114;
    wire N__32111;
    wire N__32106;
    wire N__32103;
    wire N__32098;
    wire N__32095;
    wire N__32090;
    wire N__32089;
    wire N__32088;
    wire N__32087;
    wire N__32086;
    wire N__32085;
    wire N__32084;
    wire N__32083;
    wire N__32082;
    wire N__32081;
    wire N__32080;
    wire N__32079;
    wire N__32078;
    wire N__32077;
    wire N__32076;
    wire N__32075;
    wire N__32074;
    wire N__32073;
    wire N__32072;
    wire N__32071;
    wire N__32070;
    wire N__32069;
    wire N__32068;
    wire N__32067;
    wire N__32066;
    wire N__32065;
    wire N__32064;
    wire N__32063;
    wire N__32062;
    wire N__32061;
    wire N__32056;
    wire N__32047;
    wire N__32038;
    wire N__32029;
    wire N__32020;
    wire N__32011;
    wire N__32002;
    wire N__31993;
    wire N__31988;
    wire N__31983;
    wire N__31978;
    wire N__31973;
    wire N__31970;
    wire N__31967;
    wire N__31964;
    wire N__31955;
    wire N__31952;
    wire N__31949;
    wire N__31946;
    wire N__31943;
    wire N__31940;
    wire N__31937;
    wire N__31934;
    wire N__31931;
    wire N__31928;
    wire N__31925;
    wire N__31922;
    wire N__31919;
    wire N__31916;
    wire N__31913;
    wire N__31910;
    wire N__31907;
    wire N__31904;
    wire N__31903;
    wire N__31900;
    wire N__31897;
    wire N__31894;
    wire N__31891;
    wire N__31886;
    wire N__31883;
    wire N__31880;
    wire N__31877;
    wire N__31874;
    wire N__31871;
    wire N__31868;
    wire N__31867;
    wire N__31866;
    wire N__31863;
    wire N__31860;
    wire N__31859;
    wire N__31856;
    wire N__31853;
    wire N__31850;
    wire N__31847;
    wire N__31842;
    wire N__31837;
    wire N__31832;
    wire N__31829;
    wire N__31826;
    wire N__31825;
    wire N__31824;
    wire N__31823;
    wire N__31820;
    wire N__31817;
    wire N__31814;
    wire N__31811;
    wire N__31806;
    wire N__31803;
    wire N__31796;
    wire N__31793;
    wire N__31790;
    wire N__31787;
    wire N__31784;
    wire N__31783;
    wire N__31782;
    wire N__31779;
    wire N__31774;
    wire N__31769;
    wire N__31768;
    wire N__31765;
    wire N__31762;
    wire N__31759;
    wire N__31756;
    wire N__31751;
    wire N__31750;
    wire N__31749;
    wire N__31748;
    wire N__31743;
    wire N__31740;
    wire N__31737;
    wire N__31730;
    wire N__31727;
    wire N__31724;
    wire N__31721;
    wire N__31718;
    wire N__31715;
    wire N__31712;
    wire N__31709;
    wire N__31706;
    wire N__31705;
    wire N__31704;
    wire N__31701;
    wire N__31698;
    wire N__31695;
    wire N__31692;
    wire N__31689;
    wire N__31686;
    wire N__31679;
    wire N__31676;
    wire N__31675;
    wire N__31672;
    wire N__31671;
    wire N__31668;
    wire N__31665;
    wire N__31662;
    wire N__31655;
    wire N__31654;
    wire N__31651;
    wire N__31648;
    wire N__31645;
    wire N__31642;
    wire N__31639;
    wire N__31636;
    wire N__31631;
    wire N__31628;
    wire N__31627;
    wire N__31626;
    wire N__31623;
    wire N__31622;
    wire N__31617;
    wire N__31614;
    wire N__31611;
    wire N__31608;
    wire N__31603;
    wire N__31600;
    wire N__31597;
    wire N__31592;
    wire N__31589;
    wire N__31588;
    wire N__31587;
    wire N__31584;
    wire N__31581;
    wire N__31578;
    wire N__31573;
    wire N__31572;
    wire N__31569;
    wire N__31566;
    wire N__31563;
    wire N__31556;
    wire N__31553;
    wire N__31550;
    wire N__31549;
    wire N__31548;
    wire N__31545;
    wire N__31544;
    wire N__31541;
    wire N__31538;
    wire N__31535;
    wire N__31532;
    wire N__31529;
    wire N__31526;
    wire N__31521;
    wire N__31518;
    wire N__31515;
    wire N__31508;
    wire N__31507;
    wire N__31504;
    wire N__31503;
    wire N__31502;
    wire N__31499;
    wire N__31496;
    wire N__31491;
    wire N__31488;
    wire N__31481;
    wire N__31478;
    wire N__31475;
    wire N__31472;
    wire N__31469;
    wire N__31466;
    wire N__31463;
    wire N__31460;
    wire N__31457;
    wire N__31454;
    wire N__31451;
    wire N__31448;
    wire N__31445;
    wire N__31442;
    wire N__31439;
    wire N__31436;
    wire N__31435;
    wire N__31432;
    wire N__31429;
    wire N__31426;
    wire N__31423;
    wire N__31418;
    wire N__31417;
    wire N__31414;
    wire N__31411;
    wire N__31408;
    wire N__31405;
    wire N__31400;
    wire N__31397;
    wire N__31394;
    wire N__31391;
    wire N__31388;
    wire N__31385;
    wire N__31382;
    wire N__31379;
    wire N__31376;
    wire N__31373;
    wire N__31370;
    wire N__31367;
    wire N__31364;
    wire N__31361;
    wire N__31358;
    wire N__31355;
    wire N__31352;
    wire N__31349;
    wire N__31346;
    wire N__31343;
    wire N__31340;
    wire N__31337;
    wire N__31334;
    wire N__31331;
    wire N__31328;
    wire N__31325;
    wire N__31322;
    wire N__31319;
    wire N__31316;
    wire N__31313;
    wire N__31310;
    wire N__31307;
    wire N__31304;
    wire N__31301;
    wire N__31298;
    wire N__31295;
    wire N__31292;
    wire N__31289;
    wire N__31286;
    wire N__31283;
    wire N__31280;
    wire N__31277;
    wire N__31274;
    wire N__31271;
    wire N__31268;
    wire N__31265;
    wire N__31262;
    wire N__31259;
    wire N__31256;
    wire N__31253;
    wire N__31250;
    wire N__31247;
    wire N__31244;
    wire N__31241;
    wire N__31238;
    wire N__31235;
    wire N__31232;
    wire N__31229;
    wire N__31228;
    wire N__31227;
    wire N__31226;
    wire N__31225;
    wire N__31224;
    wire N__31221;
    wire N__31218;
    wire N__31215;
    wire N__31212;
    wire N__31209;
    wire N__31206;
    wire N__31203;
    wire N__31200;
    wire N__31197;
    wire N__31194;
    wire N__31191;
    wire N__31188;
    wire N__31185;
    wire N__31180;
    wire N__31177;
    wire N__31174;
    wire N__31163;
    wire N__31160;
    wire N__31157;
    wire N__31154;
    wire N__31151;
    wire N__31148;
    wire N__31145;
    wire N__31142;
    wire N__31139;
    wire N__31138;
    wire N__31135;
    wire N__31132;
    wire N__31129;
    wire N__31124;
    wire N__31121;
    wire N__31118;
    wire N__31115;
    wire N__31112;
    wire N__31111;
    wire N__31110;
    wire N__31107;
    wire N__31106;
    wire N__31101;
    wire N__31098;
    wire N__31095;
    wire N__31092;
    wire N__31085;
    wire N__31082;
    wire N__31079;
    wire N__31076;
    wire N__31073;
    wire N__31072;
    wire N__31071;
    wire N__31070;
    wire N__31067;
    wire N__31062;
    wire N__31059;
    wire N__31054;
    wire N__31051;
    wire N__31046;
    wire N__31045;
    wire N__31042;
    wire N__31041;
    wire N__31034;
    wire N__31033;
    wire N__31030;
    wire N__31027;
    wire N__31022;
    wire N__31019;
    wire N__31016;
    wire N__31013;
    wire N__31010;
    wire N__31007;
    wire N__31004;
    wire N__31003;
    wire N__31002;
    wire N__30999;
    wire N__30996;
    wire N__30993;
    wire N__30992;
    wire N__30989;
    wire N__30984;
    wire N__30981;
    wire N__30978;
    wire N__30973;
    wire N__30968;
    wire N__30965;
    wire N__30964;
    wire N__30963;
    wire N__30960;
    wire N__30955;
    wire N__30954;
    wire N__30951;
    wire N__30948;
    wire N__30945;
    wire N__30938;
    wire N__30935;
    wire N__30932;
    wire N__30929;
    wire N__30926;
    wire N__30923;
    wire N__30920;
    wire N__30917;
    wire N__30914;
    wire N__30911;
    wire N__30908;
    wire N__30905;
    wire N__30902;
    wire N__30899;
    wire N__30896;
    wire N__30893;
    wire N__30890;
    wire N__30887;
    wire N__30884;
    wire N__30883;
    wire N__30880;
    wire N__30879;
    wire N__30876;
    wire N__30873;
    wire N__30870;
    wire N__30869;
    wire N__30864;
    wire N__30861;
    wire N__30858;
    wire N__30855;
    wire N__30852;
    wire N__30849;
    wire N__30842;
    wire N__30839;
    wire N__30838;
    wire N__30835;
    wire N__30832;
    wire N__30831;
    wire N__30828;
    wire N__30827;
    wire N__30824;
    wire N__30821;
    wire N__30818;
    wire N__30815;
    wire N__30812;
    wire N__30809;
    wire N__30800;
    wire N__30797;
    wire N__30794;
    wire N__30791;
    wire N__30788;
    wire N__30785;
    wire N__30782;
    wire N__30779;
    wire N__30776;
    wire N__30773;
    wire N__30772;
    wire N__30771;
    wire N__30768;
    wire N__30763;
    wire N__30762;
    wire N__30759;
    wire N__30756;
    wire N__30753;
    wire N__30750;
    wire N__30745;
    wire N__30740;
    wire N__30739;
    wire N__30738;
    wire N__30737;
    wire N__30730;
    wire N__30727;
    wire N__30724;
    wire N__30721;
    wire N__30716;
    wire N__30715;
    wire N__30712;
    wire N__30709;
    wire N__30708;
    wire N__30707;
    wire N__30704;
    wire N__30701;
    wire N__30698;
    wire N__30695;
    wire N__30688;
    wire N__30685;
    wire N__30680;
    wire N__30679;
    wire N__30676;
    wire N__30673;
    wire N__30672;
    wire N__30669;
    wire N__30664;
    wire N__30663;
    wire N__30658;
    wire N__30655;
    wire N__30650;
    wire N__30647;
    wire N__30644;
    wire N__30641;
    wire N__30638;
    wire N__30635;
    wire N__30632;
    wire N__30631;
    wire N__30630;
    wire N__30627;
    wire N__30624;
    wire N__30621;
    wire N__30618;
    wire N__30615;
    wire N__30612;
    wire N__30605;
    wire N__30604;
    wire N__30603;
    wire N__30600;
    wire N__30599;
    wire N__30598;
    wire N__30595;
    wire N__30594;
    wire N__30591;
    wire N__30590;
    wire N__30587;
    wire N__30584;
    wire N__30575;
    wire N__30574;
    wire N__30571;
    wire N__30564;
    wire N__30561;
    wire N__30560;
    wire N__30557;
    wire N__30554;
    wire N__30551;
    wire N__30548;
    wire N__30539;
    wire N__30536;
    wire N__30533;
    wire N__30530;
    wire N__30529;
    wire N__30526;
    wire N__30523;
    wire N__30520;
    wire N__30517;
    wire N__30514;
    wire N__30511;
    wire N__30508;
    wire N__30505;
    wire N__30500;
    wire N__30499;
    wire N__30496;
    wire N__30493;
    wire N__30490;
    wire N__30489;
    wire N__30484;
    wire N__30481;
    wire N__30476;
    wire N__30473;
    wire N__30470;
    wire N__30467;
    wire N__30464;
    wire N__30463;
    wire N__30462;
    wire N__30459;
    wire N__30456;
    wire N__30453;
    wire N__30452;
    wire N__30449;
    wire N__30446;
    wire N__30443;
    wire N__30440;
    wire N__30435;
    wire N__30430;
    wire N__30425;
    wire N__30424;
    wire N__30421;
    wire N__30418;
    wire N__30417;
    wire N__30416;
    wire N__30413;
    wire N__30410;
    wire N__30407;
    wire N__30404;
    wire N__30401;
    wire N__30398;
    wire N__30395;
    wire N__30392;
    wire N__30383;
    wire N__30380;
    wire N__30377;
    wire N__30374;
    wire N__30371;
    wire N__30368;
    wire N__30365;
    wire N__30362;
    wire N__30359;
    wire N__30358;
    wire N__30357;
    wire N__30354;
    wire N__30351;
    wire N__30350;
    wire N__30347;
    wire N__30344;
    wire N__30341;
    wire N__30338;
    wire N__30335;
    wire N__30332;
    wire N__30325;
    wire N__30320;
    wire N__30319;
    wire N__30316;
    wire N__30313;
    wire N__30312;
    wire N__30307;
    wire N__30304;
    wire N__30303;
    wire N__30300;
    wire N__30297;
    wire N__30294;
    wire N__30287;
    wire N__30284;
    wire N__30281;
    wire N__30278;
    wire N__30275;
    wire N__30272;
    wire N__30271;
    wire N__30270;
    wire N__30269;
    wire N__30266;
    wire N__30263;
    wire N__30260;
    wire N__30257;
    wire N__30254;
    wire N__30251;
    wire N__30246;
    wire N__30239;
    wire N__30236;
    wire N__30235;
    wire N__30234;
    wire N__30233;
    wire N__30226;
    wire N__30223;
    wire N__30220;
    wire N__30217;
    wire N__30212;
    wire N__30211;
    wire N__30208;
    wire N__30207;
    wire N__30204;
    wire N__30201;
    wire N__30198;
    wire N__30197;
    wire N__30194;
    wire N__30191;
    wire N__30188;
    wire N__30185;
    wire N__30182;
    wire N__30177;
    wire N__30174;
    wire N__30167;
    wire N__30166;
    wire N__30165;
    wire N__30164;
    wire N__30157;
    wire N__30154;
    wire N__30151;
    wire N__30148;
    wire N__30145;
    wire N__30142;
    wire N__30137;
    wire N__30134;
    wire N__30131;
    wire N__30128;
    wire N__30125;
    wire N__30122;
    wire N__30121;
    wire N__30120;
    wire N__30117;
    wire N__30112;
    wire N__30111;
    wire N__30108;
    wire N__30105;
    wire N__30102;
    wire N__30099;
    wire N__30096;
    wire N__30093;
    wire N__30086;
    wire N__30083;
    wire N__30080;
    wire N__30077;
    wire N__30074;
    wire N__30073;
    wire N__30070;
    wire N__30069;
    wire N__30066;
    wire N__30065;
    wire N__30062;
    wire N__30059;
    wire N__30056;
    wire N__30053;
    wire N__30044;
    wire N__30041;
    wire N__30038;
    wire N__30037;
    wire N__30034;
    wire N__30031;
    wire N__30030;
    wire N__30029;
    wire N__30024;
    wire N__30021;
    wire N__30018;
    wire N__30015;
    wire N__30012;
    wire N__30009;
    wire N__30002;
    wire N__29999;
    wire N__29996;
    wire N__29993;
    wire N__29990;
    wire N__29987;
    wire N__29984;
    wire N__29981;
    wire N__29978;
    wire N__29975;
    wire N__29972;
    wire N__29969;
    wire N__29968;
    wire N__29967;
    wire N__29964;
    wire N__29961;
    wire N__29958;
    wire N__29957;
    wire N__29952;
    wire N__29949;
    wire N__29946;
    wire N__29943;
    wire N__29938;
    wire N__29933;
    wire N__29930;
    wire N__29929;
    wire N__29926;
    wire N__29925;
    wire N__29922;
    wire N__29921;
    wire N__29918;
    wire N__29915;
    wire N__29912;
    wire N__29909;
    wire N__29904;
    wire N__29901;
    wire N__29898;
    wire N__29891;
    wire N__29888;
    wire N__29885;
    wire N__29882;
    wire N__29881;
    wire N__29880;
    wire N__29877;
    wire N__29874;
    wire N__29873;
    wire N__29870;
    wire N__29865;
    wire N__29862;
    wire N__29859;
    wire N__29856;
    wire N__29853;
    wire N__29846;
    wire N__29845;
    wire N__29842;
    wire N__29839;
    wire N__29838;
    wire N__29837;
    wire N__29834;
    wire N__29831;
    wire N__29828;
    wire N__29825;
    wire N__29822;
    wire N__29817;
    wire N__29814;
    wire N__29807;
    wire N__29804;
    wire N__29801;
    wire N__29798;
    wire N__29795;
    wire N__29792;
    wire N__29789;
    wire N__29786;
    wire N__29783;
    wire N__29780;
    wire N__29779;
    wire N__29778;
    wire N__29771;
    wire N__29770;
    wire N__29767;
    wire N__29764;
    wire N__29761;
    wire N__29758;
    wire N__29753;
    wire N__29750;
    wire N__29747;
    wire N__29744;
    wire N__29741;
    wire N__29738;
    wire N__29737;
    wire N__29736;
    wire N__29733;
    wire N__29728;
    wire N__29725;
    wire N__29722;
    wire N__29721;
    wire N__29718;
    wire N__29715;
    wire N__29712;
    wire N__29705;
    wire N__29702;
    wire N__29699;
    wire N__29696;
    wire N__29693;
    wire N__29690;
    wire N__29687;
    wire N__29684;
    wire N__29681;
    wire N__29680;
    wire N__29679;
    wire N__29676;
    wire N__29671;
    wire N__29670;
    wire N__29667;
    wire N__29664;
    wire N__29661;
    wire N__29656;
    wire N__29653;
    wire N__29648;
    wire N__29645;
    wire N__29642;
    wire N__29641;
    wire N__29640;
    wire N__29637;
    wire N__29632;
    wire N__29631;
    wire N__29628;
    wire N__29625;
    wire N__29622;
    wire N__29615;
    wire N__29614;
    wire N__29611;
    wire N__29608;
    wire N__29605;
    wire N__29604;
    wire N__29599;
    wire N__29596;
    wire N__29593;
    wire N__29590;
    wire N__29585;
    wire N__29582;
    wire N__29581;
    wire N__29578;
    wire N__29575;
    wire N__29570;
    wire N__29569;
    wire N__29566;
    wire N__29563;
    wire N__29558;
    wire N__29555;
    wire N__29552;
    wire N__29549;
    wire N__29548;
    wire N__29545;
    wire N__29542;
    wire N__29537;
    wire N__29534;
    wire N__29531;
    wire N__29530;
    wire N__29529;
    wire N__29526;
    wire N__29523;
    wire N__29520;
    wire N__29519;
    wire N__29514;
    wire N__29511;
    wire N__29508;
    wire N__29505;
    wire N__29502;
    wire N__29499;
    wire N__29492;
    wire N__29489;
    wire N__29488;
    wire N__29487;
    wire N__29484;
    wire N__29479;
    wire N__29476;
    wire N__29473;
    wire N__29472;
    wire N__29469;
    wire N__29466;
    wire N__29463;
    wire N__29456;
    wire N__29453;
    wire N__29452;
    wire N__29451;
    wire N__29448;
    wire N__29443;
    wire N__29442;
    wire N__29439;
    wire N__29436;
    wire N__29433;
    wire N__29430;
    wire N__29427;
    wire N__29424;
    wire N__29417;
    wire N__29414;
    wire N__29411;
    wire N__29408;
    wire N__29407;
    wire N__29404;
    wire N__29403;
    wire N__29400;
    wire N__29397;
    wire N__29392;
    wire N__29391;
    wire N__29388;
    wire N__29385;
    wire N__29382;
    wire N__29379;
    wire N__29376;
    wire N__29373;
    wire N__29366;
    wire N__29363;
    wire N__29360;
    wire N__29357;
    wire N__29354;
    wire N__29351;
    wire N__29348;
    wire N__29345;
    wire N__29342;
    wire N__29339;
    wire N__29336;
    wire N__29333;
    wire N__29330;
    wire N__29327;
    wire N__29326;
    wire N__29325;
    wire N__29322;
    wire N__29319;
    wire N__29316;
    wire N__29313;
    wire N__29306;
    wire N__29303;
    wire N__29300;
    wire N__29297;
    wire N__29294;
    wire N__29293;
    wire N__29290;
    wire N__29287;
    wire N__29282;
    wire N__29279;
    wire N__29278;
    wire N__29275;
    wire N__29272;
    wire N__29269;
    wire N__29264;
    wire N__29261;
    wire N__29258;
    wire N__29255;
    wire N__29254;
    wire N__29251;
    wire N__29248;
    wire N__29245;
    wire N__29242;
    wire N__29237;
    wire N__29234;
    wire N__29231;
    wire N__29228;
    wire N__29225;
    wire N__29222;
    wire N__29221;
    wire N__29218;
    wire N__29215;
    wire N__29212;
    wire N__29207;
    wire N__29204;
    wire N__29201;
    wire N__29198;
    wire N__29195;
    wire N__29194;
    wire N__29191;
    wire N__29188;
    wire N__29185;
    wire N__29180;
    wire N__29177;
    wire N__29174;
    wire N__29171;
    wire N__29168;
    wire N__29167;
    wire N__29164;
    wire N__29161;
    wire N__29158;
    wire N__29153;
    wire N__29150;
    wire N__29147;
    wire N__29144;
    wire N__29141;
    wire N__29140;
    wire N__29137;
    wire N__29134;
    wire N__29131;
    wire N__29126;
    wire N__29123;
    wire N__29120;
    wire N__29117;
    wire N__29114;
    wire N__29113;
    wire N__29110;
    wire N__29107;
    wire N__29104;
    wire N__29099;
    wire N__29096;
    wire N__29093;
    wire N__29090;
    wire N__29087;
    wire N__29084;
    wire N__29081;
    wire N__29078;
    wire N__29075;
    wire N__29074;
    wire N__29071;
    wire N__29068;
    wire N__29063;
    wire N__29060;
    wire N__29057;
    wire N__29054;
    wire N__29051;
    wire N__29048;
    wire N__29045;
    wire N__29042;
    wire N__29041;
    wire N__29038;
    wire N__29035;
    wire N__29030;
    wire N__29027;
    wire N__29024;
    wire N__29021;
    wire N__29018;
    wire N__29015;
    wire N__29012;
    wire N__29009;
    wire N__29008;
    wire N__29005;
    wire N__29002;
    wire N__28997;
    wire N__28994;
    wire N__28991;
    wire N__28988;
    wire N__28985;
    wire N__28982;
    wire N__28979;
    wire N__28978;
    wire N__28975;
    wire N__28972;
    wire N__28967;
    wire N__28964;
    wire N__28961;
    wire N__28958;
    wire N__28955;
    wire N__28952;
    wire N__28949;
    wire N__28946;
    wire N__28945;
    wire N__28942;
    wire N__28939;
    wire N__28936;
    wire N__28933;
    wire N__28928;
    wire N__28925;
    wire N__28922;
    wire N__28919;
    wire N__28916;
    wire N__28915;
    wire N__28912;
    wire N__28909;
    wire N__28906;
    wire N__28903;
    wire N__28900;
    wire N__28895;
    wire N__28892;
    wire N__28889;
    wire N__28886;
    wire N__28885;
    wire N__28882;
    wire N__28879;
    wire N__28876;
    wire N__28873;
    wire N__28870;
    wire N__28865;
    wire N__28862;
    wire N__28859;
    wire N__28856;
    wire N__28855;
    wire N__28854;
    wire N__28853;
    wire N__28852;
    wire N__28851;
    wire N__28850;
    wire N__28849;
    wire N__28848;
    wire N__28847;
    wire N__28846;
    wire N__28845;
    wire N__28844;
    wire N__28843;
    wire N__28842;
    wire N__28841;
    wire N__28840;
    wire N__28839;
    wire N__28838;
    wire N__28837;
    wire N__28836;
    wire N__28835;
    wire N__28834;
    wire N__28833;
    wire N__28832;
    wire N__28831;
    wire N__28830;
    wire N__28829;
    wire N__28828;
    wire N__28827;
    wire N__28824;
    wire N__28823;
    wire N__28822;
    wire N__28821;
    wire N__28820;
    wire N__28819;
    wire N__28818;
    wire N__28817;
    wire N__28810;
    wire N__28801;
    wire N__28800;
    wire N__28797;
    wire N__28796;
    wire N__28793;
    wire N__28792;
    wire N__28789;
    wire N__28786;
    wire N__28783;
    wire N__28780;
    wire N__28777;
    wire N__28774;
    wire N__28771;
    wire N__28768;
    wire N__28765;
    wire N__28762;
    wire N__28759;
    wire N__28756;
    wire N__28753;
    wire N__28750;
    wire N__28747;
    wire N__28744;
    wire N__28741;
    wire N__28738;
    wire N__28735;
    wire N__28732;
    wire N__28731;
    wire N__28728;
    wire N__28721;
    wire N__28712;
    wire N__28707;
    wire N__28700;
    wire N__28699;
    wire N__28698;
    wire N__28697;
    wire N__28696;
    wire N__28695;
    wire N__28694;
    wire N__28693;
    wire N__28682;
    wire N__28675;
    wire N__28666;
    wire N__28657;
    wire N__28656;
    wire N__28649;
    wire N__28642;
    wire N__28639;
    wire N__28632;
    wire N__28627;
    wire N__28624;
    wire N__28621;
    wire N__28618;
    wire N__28615;
    wire N__28612;
    wire N__28609;
    wire N__28606;
    wire N__28603;
    wire N__28600;
    wire N__28595;
    wire N__28592;
    wire N__28587;
    wire N__28582;
    wire N__28579;
    wire N__28572;
    wire N__28563;
    wire N__28558;
    wire N__28555;
    wire N__28552;
    wire N__28549;
    wire N__28548;
    wire N__28547;
    wire N__28544;
    wire N__28537;
    wire N__28532;
    wire N__28529;
    wire N__28528;
    wire N__28525;
    wire N__28522;
    wire N__28519;
    wire N__28516;
    wire N__28513;
    wire N__28510;
    wire N__28507;
    wire N__28504;
    wire N__28501;
    wire N__28496;
    wire N__28493;
    wire N__28486;
    wire N__28483;
    wire N__28478;
    wire N__28469;
    wire N__28466;
    wire N__28463;
    wire N__28460;
    wire N__28457;
    wire N__28454;
    wire N__28451;
    wire N__28448;
    wire N__28445;
    wire N__28442;
    wire N__28439;
    wire N__28436;
    wire N__28433;
    wire N__28430;
    wire N__28427;
    wire N__28424;
    wire N__28421;
    wire N__28418;
    wire N__28415;
    wire N__28412;
    wire N__28409;
    wire N__28406;
    wire N__28403;
    wire N__28400;
    wire N__28397;
    wire N__28394;
    wire N__28391;
    wire N__28388;
    wire N__28387;
    wire N__28384;
    wire N__28381;
    wire N__28378;
    wire N__28377;
    wire N__28374;
    wire N__28371;
    wire N__28368;
    wire N__28361;
    wire N__28358;
    wire N__28355;
    wire N__28354;
    wire N__28351;
    wire N__28348;
    wire N__28343;
    wire N__28340;
    wire N__28337;
    wire N__28334;
    wire N__28331;
    wire N__28328;
    wire N__28325;
    wire N__28322;
    wire N__28319;
    wire N__28316;
    wire N__28313;
    wire N__28312;
    wire N__28309;
    wire N__28306;
    wire N__28301;
    wire N__28298;
    wire N__28295;
    wire N__28292;
    wire N__28289;
    wire N__28286;
    wire N__28283;
    wire N__28280;
    wire N__28279;
    wire N__28276;
    wire N__28273;
    wire N__28268;
    wire N__28265;
    wire N__28262;
    wire N__28259;
    wire N__28256;
    wire N__28253;
    wire N__28250;
    wire N__28249;
    wire N__28248;
    wire N__28247;
    wire N__28240;
    wire N__28237;
    wire N__28234;
    wire N__28231;
    wire N__28226;
    wire N__28223;
    wire N__28220;
    wire N__28217;
    wire N__28214;
    wire N__28211;
    wire N__28208;
    wire N__28205;
    wire N__28202;
    wire N__28199;
    wire N__28196;
    wire N__28193;
    wire N__28190;
    wire N__28187;
    wire N__28184;
    wire N__28181;
    wire N__28178;
    wire N__28175;
    wire N__28172;
    wire N__28169;
    wire N__28166;
    wire N__28163;
    wire N__28160;
    wire N__28157;
    wire N__28154;
    wire N__28151;
    wire N__28148;
    wire N__28145;
    wire N__28144;
    wire N__28141;
    wire N__28140;
    wire N__28139;
    wire N__28136;
    wire N__28131;
    wire N__28128;
    wire N__28123;
    wire N__28120;
    wire N__28115;
    wire N__28112;
    wire N__28109;
    wire N__28106;
    wire N__28103;
    wire N__28100;
    wire N__28097;
    wire N__28094;
    wire N__28091;
    wire N__28088;
    wire N__28085;
    wire N__28082;
    wire N__28079;
    wire N__28076;
    wire N__28073;
    wire N__28070;
    wire N__28067;
    wire N__28064;
    wire N__28061;
    wire N__28058;
    wire N__28055;
    wire N__28052;
    wire N__28049;
    wire N__28046;
    wire N__28043;
    wire N__28040;
    wire N__28037;
    wire N__28034;
    wire N__28031;
    wire N__28028;
    wire N__28025;
    wire N__28022;
    wire N__28019;
    wire N__28016;
    wire N__28013;
    wire N__28010;
    wire N__28007;
    wire N__28004;
    wire N__28001;
    wire N__28000;
    wire N__27997;
    wire N__27994;
    wire N__27993;
    wire N__27992;
    wire N__27989;
    wire N__27984;
    wire N__27981;
    wire N__27976;
    wire N__27973;
    wire N__27968;
    wire N__27965;
    wire N__27962;
    wire N__27959;
    wire N__27956;
    wire N__27953;
    wire N__27950;
    wire N__27949;
    wire N__27948;
    wire N__27945;
    wire N__27940;
    wire N__27939;
    wire N__27934;
    wire N__27931;
    wire N__27928;
    wire N__27925;
    wire N__27920;
    wire N__27917;
    wire N__27914;
    wire N__27911;
    wire N__27908;
    wire N__27905;
    wire N__27902;
    wire N__27899;
    wire N__27896;
    wire N__27893;
    wire N__27890;
    wire N__27887;
    wire N__27884;
    wire N__27881;
    wire N__27878;
    wire N__27875;
    wire N__27872;
    wire N__27869;
    wire N__27866;
    wire N__27863;
    wire N__27860;
    wire N__27857;
    wire N__27854;
    wire N__27853;
    wire N__27852;
    wire N__27849;
    wire N__27846;
    wire N__27843;
    wire N__27842;
    wire N__27835;
    wire N__27832;
    wire N__27829;
    wire N__27826;
    wire N__27821;
    wire N__27818;
    wire N__27815;
    wire N__27812;
    wire N__27809;
    wire N__27806;
    wire N__27803;
    wire N__27800;
    wire N__27799;
    wire N__27798;
    wire N__27797;
    wire N__27794;
    wire N__27789;
    wire N__27786;
    wire N__27783;
    wire N__27778;
    wire N__27773;
    wire N__27770;
    wire N__27767;
    wire N__27764;
    wire N__27761;
    wire N__27758;
    wire N__27757;
    wire N__27756;
    wire N__27753;
    wire N__27752;
    wire N__27749;
    wire N__27746;
    wire N__27741;
    wire N__27738;
    wire N__27735;
    wire N__27732;
    wire N__27729;
    wire N__27722;
    wire N__27719;
    wire N__27716;
    wire N__27713;
    wire N__27710;
    wire N__27707;
    wire N__27704;
    wire N__27701;
    wire N__27698;
    wire N__27695;
    wire N__27692;
    wire N__27689;
    wire N__27686;
    wire N__27683;
    wire N__27680;
    wire N__27677;
    wire N__27676;
    wire N__27675;
    wire N__27674;
    wire N__27669;
    wire N__27666;
    wire N__27663;
    wire N__27660;
    wire N__27655;
    wire N__27650;
    wire N__27647;
    wire N__27644;
    wire N__27641;
    wire N__27638;
    wire N__27635;
    wire N__27632;
    wire N__27629;
    wire N__27626;
    wire N__27623;
    wire N__27620;
    wire N__27617;
    wire N__27614;
    wire N__27611;
    wire N__27608;
    wire N__27605;
    wire N__27602;
    wire N__27599;
    wire N__27598;
    wire N__27597;
    wire N__27596;
    wire N__27595;
    wire N__27592;
    wire N__27591;
    wire N__27582;
    wire N__27579;
    wire N__27576;
    wire N__27569;
    wire N__27568;
    wire N__27565;
    wire N__27564;
    wire N__27563;
    wire N__27560;
    wire N__27555;
    wire N__27552;
    wire N__27545;
    wire N__27542;
    wire N__27539;
    wire N__27536;
    wire N__27533;
    wire N__27530;
    wire N__27527;
    wire N__27526;
    wire N__27521;
    wire N__27520;
    wire N__27517;
    wire N__27514;
    wire N__27509;
    wire N__27506;
    wire N__27503;
    wire N__27500;
    wire N__27497;
    wire N__27494;
    wire N__27491;
    wire N__27488;
    wire N__27487;
    wire N__27486;
    wire N__27485;
    wire N__27480;
    wire N__27477;
    wire N__27474;
    wire N__27469;
    wire N__27466;
    wire N__27461;
    wire N__27458;
    wire N__27455;
    wire N__27452;
    wire N__27449;
    wire N__27446;
    wire N__27443;
    wire N__27440;
    wire N__27437;
    wire N__27434;
    wire N__27431;
    wire N__27428;
    wire N__27425;
    wire N__27422;
    wire N__27419;
    wire N__27416;
    wire N__27413;
    wire N__27410;
    wire N__27407;
    wire N__27404;
    wire N__27401;
    wire N__27398;
    wire N__27397;
    wire N__27394;
    wire N__27393;
    wire N__27390;
    wire N__27389;
    wire N__27386;
    wire N__27383;
    wire N__27380;
    wire N__27377;
    wire N__27368;
    wire N__27365;
    wire N__27362;
    wire N__27359;
    wire N__27356;
    wire N__27353;
    wire N__27350;
    wire N__27347;
    wire N__27346;
    wire N__27345;
    wire N__27342;
    wire N__27339;
    wire N__27336;
    wire N__27329;
    wire N__27326;
    wire N__27325;
    wire N__27324;
    wire N__27321;
    wire N__27318;
    wire N__27315;
    wire N__27308;
    wire N__27305;
    wire N__27304;
    wire N__27303;
    wire N__27300;
    wire N__27297;
    wire N__27294;
    wire N__27291;
    wire N__27284;
    wire N__27281;
    wire N__27280;
    wire N__27279;
    wire N__27278;
    wire N__27277;
    wire N__27276;
    wire N__27275;
    wire N__27274;
    wire N__27273;
    wire N__27272;
    wire N__27269;
    wire N__27266;
    wire N__27257;
    wire N__27248;
    wire N__27245;
    wire N__27242;
    wire N__27233;
    wire N__27230;
    wire N__27229;
    wire N__27228;
    wire N__27225;
    wire N__27222;
    wire N__27219;
    wire N__27216;
    wire N__27209;
    wire N__27206;
    wire N__27203;
    wire N__27200;
    wire N__27197;
    wire N__27196;
    wire N__27195;
    wire N__27192;
    wire N__27189;
    wire N__27186;
    wire N__27179;
    wire N__27176;
    wire N__27175;
    wire N__27174;
    wire N__27171;
    wire N__27168;
    wire N__27165;
    wire N__27158;
    wire N__27155;
    wire N__27154;
    wire N__27153;
    wire N__27150;
    wire N__27147;
    wire N__27144;
    wire N__27137;
    wire N__27134;
    wire N__27133;
    wire N__27132;
    wire N__27129;
    wire N__27126;
    wire N__27123;
    wire N__27116;
    wire N__27113;
    wire N__27112;
    wire N__27111;
    wire N__27108;
    wire N__27105;
    wire N__27102;
    wire N__27095;
    wire N__27092;
    wire N__27091;
    wire N__27090;
    wire N__27087;
    wire N__27084;
    wire N__27081;
    wire N__27074;
    wire N__27071;
    wire N__27070;
    wire N__27067;
    wire N__27064;
    wire N__27063;
    wire N__27058;
    wire N__27055;
    wire N__27052;
    wire N__27047;
    wire N__27044;
    wire N__27043;
    wire N__27040;
    wire N__27037;
    wire N__27036;
    wire N__27031;
    wire N__27028;
    wire N__27025;
    wire N__27020;
    wire N__27017;
    wire N__27016;
    wire N__27013;
    wire N__27010;
    wire N__27005;
    wire N__27004;
    wire N__27001;
    wire N__26998;
    wire N__26995;
    wire N__26990;
    wire N__26987;
    wire N__26986;
    wire N__26983;
    wire N__26980;
    wire N__26979;
    wire N__26974;
    wire N__26971;
    wire N__26968;
    wire N__26963;
    wire N__26960;
    wire N__26957;
    wire N__26956;
    wire N__26953;
    wire N__26950;
    wire N__26947;
    wire N__26942;
    wire N__26939;
    wire N__26936;
    wire N__26935;
    wire N__26932;
    wire N__26929;
    wire N__26926;
    wire N__26921;
    wire N__26918;
    wire N__26915;
    wire N__26914;
    wire N__26911;
    wire N__26908;
    wire N__26907;
    wire N__26902;
    wire N__26899;
    wire N__26896;
    wire N__26891;
    wire N__26888;
    wire N__26887;
    wire N__26884;
    wire N__26881;
    wire N__26880;
    wire N__26875;
    wire N__26872;
    wire N__26869;
    wire N__26864;
    wire N__26861;
    wire N__26860;
    wire N__26857;
    wire N__26854;
    wire N__26849;
    wire N__26848;
    wire N__26845;
    wire N__26842;
    wire N__26839;
    wire N__26834;
    wire N__26831;
    wire N__26830;
    wire N__26827;
    wire N__26824;
    wire N__26819;
    wire N__26818;
    wire N__26815;
    wire N__26812;
    wire N__26809;
    wire N__26804;
    wire N__26801;
    wire N__26800;
    wire N__26795;
    wire N__26794;
    wire N__26791;
    wire N__26788;
    wire N__26785;
    wire N__26780;
    wire N__26777;
    wire N__26776;
    wire N__26771;
    wire N__26770;
    wire N__26767;
    wire N__26764;
    wire N__26761;
    wire N__26756;
    wire N__26753;
    wire N__26752;
    wire N__26749;
    wire N__26746;
    wire N__26741;
    wire N__26740;
    wire N__26737;
    wire N__26734;
    wire N__26731;
    wire N__26726;
    wire N__26723;
    wire N__26722;
    wire N__26719;
    wire N__26716;
    wire N__26715;
    wire N__26710;
    wire N__26707;
    wire N__26704;
    wire N__26699;
    wire N__26696;
    wire N__26695;
    wire N__26692;
    wire N__26689;
    wire N__26686;
    wire N__26685;
    wire N__26680;
    wire N__26677;
    wire N__26674;
    wire N__26669;
    wire N__26666;
    wire N__26665;
    wire N__26662;
    wire N__26659;
    wire N__26658;
    wire N__26653;
    wire N__26650;
    wire N__26647;
    wire N__26642;
    wire N__26639;
    wire N__26638;
    wire N__26635;
    wire N__26632;
    wire N__26627;
    wire N__26626;
    wire N__26623;
    wire N__26620;
    wire N__26617;
    wire N__26612;
    wire N__26609;
    wire N__26608;
    wire N__26605;
    wire N__26602;
    wire N__26601;
    wire N__26596;
    wire N__26593;
    wire N__26590;
    wire N__26585;
    wire N__26582;
    wire N__26581;
    wire N__26580;
    wire N__26575;
    wire N__26572;
    wire N__26569;
    wire N__26564;
    wire N__26561;
    wire N__26560;
    wire N__26555;
    wire N__26554;
    wire N__26551;
    wire N__26548;
    wire N__26545;
    wire N__26540;
    wire N__26537;
    wire N__26536;
    wire N__26533;
    wire N__26530;
    wire N__26529;
    wire N__26524;
    wire N__26521;
    wire N__26518;
    wire N__26513;
    wire N__26510;
    wire N__26509;
    wire N__26506;
    wire N__26503;
    wire N__26498;
    wire N__26497;
    wire N__26494;
    wire N__26491;
    wire N__26488;
    wire N__26483;
    wire N__26480;
    wire N__26477;
    wire N__26476;
    wire N__26475;
    wire N__26474;
    wire N__26473;
    wire N__26462;
    wire N__26459;
    wire N__26456;
    wire N__26455;
    wire N__26452;
    wire N__26449;
    wire N__26446;
    wire N__26443;
    wire N__26442;
    wire N__26439;
    wire N__26436;
    wire N__26433;
    wire N__26426;
    wire N__26423;
    wire N__26422;
    wire N__26419;
    wire N__26416;
    wire N__26415;
    wire N__26410;
    wire N__26407;
    wire N__26402;
    wire N__26399;
    wire N__26398;
    wire N__26395;
    wire N__26392;
    wire N__26391;
    wire N__26386;
    wire N__26383;
    wire N__26380;
    wire N__26375;
    wire N__26372;
    wire N__26371;
    wire N__26368;
    wire N__26365;
    wire N__26360;
    wire N__26359;
    wire N__26356;
    wire N__26353;
    wire N__26350;
    wire N__26345;
    wire N__26342;
    wire N__26341;
    wire N__26340;
    wire N__26335;
    wire N__26332;
    wire N__26329;
    wire N__26324;
    wire N__26321;
    wire N__26320;
    wire N__26315;
    wire N__26314;
    wire N__26311;
    wire N__26308;
    wire N__26305;
    wire N__26300;
    wire N__26297;
    wire N__26296;
    wire N__26293;
    wire N__26290;
    wire N__26287;
    wire N__26286;
    wire N__26283;
    wire N__26280;
    wire N__26277;
    wire N__26272;
    wire N__26267;
    wire N__26264;
    wire N__26263;
    wire N__26260;
    wire N__26257;
    wire N__26256;
    wire N__26251;
    wire N__26248;
    wire N__26245;
    wire N__26240;
    wire N__26237;
    wire N__26234;
    wire N__26231;
    wire N__26228;
    wire N__26225;
    wire N__26222;
    wire N__26219;
    wire N__26216;
    wire N__26213;
    wire N__26210;
    wire N__26207;
    wire N__26204;
    wire N__26201;
    wire N__26198;
    wire N__26195;
    wire N__26192;
    wire N__26189;
    wire N__26186;
    wire N__26183;
    wire N__26180;
    wire N__26177;
    wire N__26174;
    wire N__26171;
    wire N__26168;
    wire N__26165;
    wire N__26162;
    wire N__26159;
    wire N__26156;
    wire N__26153;
    wire N__26150;
    wire N__26147;
    wire N__26144;
    wire N__26141;
    wire N__26138;
    wire N__26135;
    wire N__26132;
    wire N__26129;
    wire N__26126;
    wire N__26123;
    wire N__26120;
    wire N__26117;
    wire N__26114;
    wire N__26111;
    wire N__26108;
    wire N__26105;
    wire N__26102;
    wire N__26099;
    wire N__26096;
    wire N__26093;
    wire N__26090;
    wire N__26087;
    wire N__26084;
    wire N__26081;
    wire N__26078;
    wire N__26075;
    wire N__26072;
    wire N__26069;
    wire N__26066;
    wire N__26063;
    wire N__26060;
    wire N__26057;
    wire N__26054;
    wire N__26051;
    wire N__26048;
    wire N__26045;
    wire N__26042;
    wire N__26039;
    wire N__26036;
    wire N__26033;
    wire N__26030;
    wire N__26027;
    wire N__26024;
    wire N__26021;
    wire N__26018;
    wire N__26015;
    wire N__26012;
    wire N__26009;
    wire N__26006;
    wire N__26003;
    wire N__26000;
    wire N__25997;
    wire N__25994;
    wire N__25991;
    wire N__25988;
    wire N__25985;
    wire N__25982;
    wire N__25979;
    wire N__25976;
    wire N__25973;
    wire N__25970;
    wire N__25967;
    wire N__25964;
    wire N__25961;
    wire N__25958;
    wire N__25955;
    wire N__25954;
    wire N__25951;
    wire N__25950;
    wire N__25947;
    wire N__25946;
    wire N__25943;
    wire N__25940;
    wire N__25937;
    wire N__25934;
    wire N__25927;
    wire N__25922;
    wire N__25919;
    wire N__25916;
    wire N__25913;
    wire N__25910;
    wire N__25907;
    wire N__25906;
    wire N__25905;
    wire N__25902;
    wire N__25899;
    wire N__25896;
    wire N__25893;
    wire N__25890;
    wire N__25887;
    wire N__25886;
    wire N__25883;
    wire N__25878;
    wire N__25875;
    wire N__25872;
    wire N__25865;
    wire N__25862;
    wire N__25859;
    wire N__25856;
    wire N__25853;
    wire N__25852;
    wire N__25849;
    wire N__25848;
    wire N__25847;
    wire N__25844;
    wire N__25841;
    wire N__25838;
    wire N__25835;
    wire N__25832;
    wire N__25829;
    wire N__25826;
    wire N__25823;
    wire N__25820;
    wire N__25817;
    wire N__25808;
    wire N__25805;
    wire N__25802;
    wire N__25799;
    wire N__25796;
    wire N__25795;
    wire N__25792;
    wire N__25791;
    wire N__25788;
    wire N__25787;
    wire N__25784;
    wire N__25781;
    wire N__25778;
    wire N__25775;
    wire N__25772;
    wire N__25769;
    wire N__25766;
    wire N__25763;
    wire N__25760;
    wire N__25755;
    wire N__25752;
    wire N__25745;
    wire N__25742;
    wire N__25739;
    wire N__25736;
    wire N__25733;
    wire N__25732;
    wire N__25731;
    wire N__25730;
    wire N__25729;
    wire N__25728;
    wire N__25725;
    wire N__25724;
    wire N__25721;
    wire N__25720;
    wire N__25717;
    wire N__25714;
    wire N__25699;
    wire N__25696;
    wire N__25693;
    wire N__25690;
    wire N__25687;
    wire N__25682;
    wire N__25679;
    wire N__25678;
    wire N__25677;
    wire N__25676;
    wire N__25675;
    wire N__25674;
    wire N__25673;
    wire N__25672;
    wire N__25671;
    wire N__25670;
    wire N__25669;
    wire N__25668;
    wire N__25667;
    wire N__25666;
    wire N__25665;
    wire N__25664;
    wire N__25659;
    wire N__25658;
    wire N__25655;
    wire N__25654;
    wire N__25653;
    wire N__25650;
    wire N__25649;
    wire N__25646;
    wire N__25645;
    wire N__25642;
    wire N__25639;
    wire N__25636;
    wire N__25635;
    wire N__25634;
    wire N__25633;
    wire N__25632;
    wire N__25629;
    wire N__25626;
    wire N__25623;
    wire N__25620;
    wire N__25619;
    wire N__25618;
    wire N__25615;
    wire N__25614;
    wire N__25613;
    wire N__25610;
    wire N__25607;
    wire N__25604;
    wire N__25603;
    wire N__25602;
    wire N__25601;
    wire N__25598;
    wire N__25595;
    wire N__25590;
    wire N__25587;
    wire N__25582;
    wire N__25579;
    wire N__25564;
    wire N__25561;
    wire N__25548;
    wire N__25543;
    wire N__25528;
    wire N__25525;
    wire N__25518;
    wire N__25513;
    wire N__25508;
    wire N__25493;
    wire N__25490;
    wire N__25487;
    wire N__25484;
    wire N__25481;
    wire N__25478;
    wire N__25475;
    wire N__25472;
    wire N__25469;
    wire N__25466;
    wire N__25463;
    wire N__25462;
    wire N__25461;
    wire N__25460;
    wire N__25457;
    wire N__25454;
    wire N__25449;
    wire N__25442;
    wire N__25441;
    wire N__25438;
    wire N__25435;
    wire N__25432;
    wire N__25429;
    wire N__25426;
    wire N__25423;
    wire N__25420;
    wire N__25417;
    wire N__25412;
    wire N__25409;
    wire N__25406;
    wire N__25403;
    wire N__25400;
    wire N__25397;
    wire N__25396;
    wire N__25393;
    wire N__25390;
    wire N__25387;
    wire N__25386;
    wire N__25385;
    wire N__25382;
    wire N__25379;
    wire N__25376;
    wire N__25373;
    wire N__25370;
    wire N__25361;
    wire N__25360;
    wire N__25357;
    wire N__25354;
    wire N__25351;
    wire N__25348;
    wire N__25345;
    wire N__25342;
    wire N__25339;
    wire N__25336;
    wire N__25331;
    wire N__25328;
    wire N__25325;
    wire N__25322;
    wire N__25321;
    wire N__25320;
    wire N__25317;
    wire N__25316;
    wire N__25313;
    wire N__25310;
    wire N__25307;
    wire N__25304;
    wire N__25299;
    wire N__25292;
    wire N__25289;
    wire N__25288;
    wire N__25285;
    wire N__25282;
    wire N__25279;
    wire N__25274;
    wire N__25271;
    wire N__25268;
    wire N__25265;
    wire N__25262;
    wire N__25259;
    wire N__25258;
    wire N__25257;
    wire N__25254;
    wire N__25251;
    wire N__25250;
    wire N__25247;
    wire N__25244;
    wire N__25241;
    wire N__25238;
    wire N__25235;
    wire N__25226;
    wire N__25223;
    wire N__25222;
    wire N__25219;
    wire N__25216;
    wire N__25213;
    wire N__25208;
    wire N__25205;
    wire N__25202;
    wire N__25199;
    wire N__25196;
    wire N__25193;
    wire N__25190;
    wire N__25187;
    wire N__25184;
    wire N__25181;
    wire N__25180;
    wire N__25177;
    wire N__25176;
    wire N__25173;
    wire N__25170;
    wire N__25167;
    wire N__25166;
    wire N__25163;
    wire N__25158;
    wire N__25155;
    wire N__25152;
    wire N__25145;
    wire N__25144;
    wire N__25141;
    wire N__25138;
    wire N__25135;
    wire N__25132;
    wire N__25129;
    wire N__25126;
    wire N__25123;
    wire N__25118;
    wire N__25115;
    wire N__25112;
    wire N__25109;
    wire N__25106;
    wire N__25105;
    wire N__25102;
    wire N__25101;
    wire N__25098;
    wire N__25095;
    wire N__25092;
    wire N__25091;
    wire N__25088;
    wire N__25083;
    wire N__25080;
    wire N__25077;
    wire N__25070;
    wire N__25067;
    wire N__25064;
    wire N__25061;
    wire N__25058;
    wire N__25055;
    wire N__25054;
    wire N__25051;
    wire N__25050;
    wire N__25047;
    wire N__25044;
    wire N__25041;
    wire N__25040;
    wire N__25037;
    wire N__25034;
    wire N__25031;
    wire N__25028;
    wire N__25025;
    wire N__25020;
    wire N__25017;
    wire N__25014;
    wire N__25007;
    wire N__25004;
    wire N__25001;
    wire N__24998;
    wire N__24995;
    wire N__24992;
    wire N__24989;
    wire N__24986;
    wire N__24983;
    wire N__24982;
    wire N__24979;
    wire N__24976;
    wire N__24973;
    wire N__24972;
    wire N__24971;
    wire N__24968;
    wire N__24965;
    wire N__24962;
    wire N__24959;
    wire N__24956;
    wire N__24947;
    wire N__24946;
    wire N__24943;
    wire N__24940;
    wire N__24937;
    wire N__24934;
    wire N__24931;
    wire N__24926;
    wire N__24923;
    wire N__24920;
    wire N__24917;
    wire N__24914;
    wire N__24911;
    wire N__24910;
    wire N__24907;
    wire N__24904;
    wire N__24901;
    wire N__24898;
    wire N__24895;
    wire N__24892;
    wire N__24887;
    wire N__24884;
    wire N__24881;
    wire N__24880;
    wire N__24879;
    wire N__24876;
    wire N__24875;
    wire N__24872;
    wire N__24869;
    wire N__24866;
    wire N__24863;
    wire N__24860;
    wire N__24857;
    wire N__24852;
    wire N__24845;
    wire N__24842;
    wire N__24839;
    wire N__24836;
    wire N__24833;
    wire N__24832;
    wire N__24829;
    wire N__24826;
    wire N__24825;
    wire N__24822;
    wire N__24821;
    wire N__24818;
    wire N__24815;
    wire N__24812;
    wire N__24809;
    wire N__24804;
    wire N__24797;
    wire N__24796;
    wire N__24793;
    wire N__24790;
    wire N__24787;
    wire N__24784;
    wire N__24779;
    wire N__24776;
    wire N__24773;
    wire N__24770;
    wire N__24767;
    wire N__24764;
    wire N__24761;
    wire N__24758;
    wire N__24755;
    wire N__24754;
    wire N__24753;
    wire N__24750;
    wire N__24747;
    wire N__24746;
    wire N__24743;
    wire N__24740;
    wire N__24737;
    wire N__24734;
    wire N__24731;
    wire N__24728;
    wire N__24719;
    wire N__24718;
    wire N__24715;
    wire N__24712;
    wire N__24709;
    wire N__24706;
    wire N__24703;
    wire N__24700;
    wire N__24697;
    wire N__24692;
    wire N__24689;
    wire N__24686;
    wire N__24683;
    wire N__24680;
    wire N__24679;
    wire N__24678;
    wire N__24677;
    wire N__24674;
    wire N__24671;
    wire N__24666;
    wire N__24659;
    wire N__24658;
    wire N__24655;
    wire N__24652;
    wire N__24649;
    wire N__24646;
    wire N__24643;
    wire N__24640;
    wire N__24637;
    wire N__24634;
    wire N__24629;
    wire N__24626;
    wire N__24623;
    wire N__24620;
    wire N__24617;
    wire N__24614;
    wire N__24613;
    wire N__24612;
    wire N__24611;
    wire N__24610;
    wire N__24607;
    wire N__24600;
    wire N__24599;
    wire N__24596;
    wire N__24593;
    wire N__24590;
    wire N__24587;
    wire N__24578;
    wire N__24577;
    wire N__24574;
    wire N__24571;
    wire N__24568;
    wire N__24565;
    wire N__24562;
    wire N__24559;
    wire N__24556;
    wire N__24551;
    wire N__24548;
    wire N__24545;
    wire N__24542;
    wire N__24539;
    wire N__24536;
    wire N__24535;
    wire N__24534;
    wire N__24533;
    wire N__24530;
    wire N__24527;
    wire N__24522;
    wire N__24515;
    wire N__24514;
    wire N__24511;
    wire N__24508;
    wire N__24505;
    wire N__24502;
    wire N__24499;
    wire N__24496;
    wire N__24493;
    wire N__24490;
    wire N__24485;
    wire N__24482;
    wire N__24479;
    wire N__24476;
    wire N__24473;
    wire N__24472;
    wire N__24469;
    wire N__24466;
    wire N__24465;
    wire N__24460;
    wire N__24459;
    wire N__24456;
    wire N__24453;
    wire N__24448;
    wire N__24443;
    wire N__24442;
    wire N__24439;
    wire N__24436;
    wire N__24433;
    wire N__24430;
    wire N__24427;
    wire N__24424;
    wire N__24421;
    wire N__24418;
    wire N__24413;
    wire N__24410;
    wire N__24407;
    wire N__24404;
    wire N__24401;
    wire N__24398;
    wire N__24395;
    wire N__24394;
    wire N__24391;
    wire N__24388;
    wire N__24387;
    wire N__24386;
    wire N__24381;
    wire N__24376;
    wire N__24373;
    wire N__24370;
    wire N__24365;
    wire N__24364;
    wire N__24361;
    wire N__24358;
    wire N__24355;
    wire N__24352;
    wire N__24349;
    wire N__24344;
    wire N__24341;
    wire N__24338;
    wire N__24335;
    wire N__24332;
    wire N__24329;
    wire N__24326;
    wire N__24323;
    wire N__24320;
    wire N__24317;
    wire N__24316;
    wire N__24313;
    wire N__24310;
    wire N__24307;
    wire N__24302;
    wire N__24299;
    wire N__24298;
    wire N__24295;
    wire N__24292;
    wire N__24291;
    wire N__24290;
    wire N__24287;
    wire N__24284;
    wire N__24279;
    wire N__24272;
    wire N__24269;
    wire N__24266;
    wire N__24263;
    wire N__24260;
    wire N__24257;
    wire N__24256;
    wire N__24255;
    wire N__24254;
    wire N__24251;
    wire N__24248;
    wire N__24243;
    wire N__24236;
    wire N__24235;
    wire N__24232;
    wire N__24229;
    wire N__24226;
    wire N__24223;
    wire N__24220;
    wire N__24217;
    wire N__24214;
    wire N__24211;
    wire N__24206;
    wire N__24203;
    wire N__24200;
    wire N__24197;
    wire N__24194;
    wire N__24191;
    wire N__24190;
    wire N__24189;
    wire N__24188;
    wire N__24185;
    wire N__24180;
    wire N__24177;
    wire N__24170;
    wire N__24169;
    wire N__24166;
    wire N__24163;
    wire N__24160;
    wire N__24157;
    wire N__24154;
    wire N__24151;
    wire N__24148;
    wire N__24145;
    wire N__24140;
    wire N__24137;
    wire N__24134;
    wire N__24131;
    wire N__24128;
    wire N__24127;
    wire N__24126;
    wire N__24123;
    wire N__24120;
    wire N__24119;
    wire N__24116;
    wire N__24111;
    wire N__24108;
    wire N__24101;
    wire N__24100;
    wire N__24097;
    wire N__24094;
    wire N__24091;
    wire N__24088;
    wire N__24085;
    wire N__24080;
    wire N__24077;
    wire N__24074;
    wire N__24071;
    wire N__24068;
    wire N__24065;
    wire N__24064;
    wire N__24063;
    wire N__24060;
    wire N__24057;
    wire N__24054;
    wire N__24051;
    wire N__24050;
    wire N__24047;
    wire N__24042;
    wire N__24039;
    wire N__24032;
    wire N__24031;
    wire N__24028;
    wire N__24025;
    wire N__24022;
    wire N__24019;
    wire N__24016;
    wire N__24013;
    wire N__24010;
    wire N__24007;
    wire N__24002;
    wire N__23999;
    wire N__23996;
    wire N__23993;
    wire N__23990;
    wire N__23989;
    wire N__23988;
    wire N__23985;
    wire N__23982;
    wire N__23981;
    wire N__23978;
    wire N__23975;
    wire N__23972;
    wire N__23969;
    wire N__23964;
    wire N__23957;
    wire N__23956;
    wire N__23953;
    wire N__23950;
    wire N__23947;
    wire N__23944;
    wire N__23941;
    wire N__23938;
    wire N__23935;
    wire N__23930;
    wire N__23927;
    wire N__23924;
    wire N__23921;
    wire N__23918;
    wire N__23915;
    wire N__23912;
    wire N__23911;
    wire N__23908;
    wire N__23905;
    wire N__23902;
    wire N__23899;
    wire N__23896;
    wire N__23891;
    wire N__23888;
    wire N__23885;
    wire N__23882;
    wire N__23881;
    wire N__23880;
    wire N__23877;
    wire N__23874;
    wire N__23871;
    wire N__23864;
    wire N__23863;
    wire N__23860;
    wire N__23857;
    wire N__23854;
    wire N__23851;
    wire N__23848;
    wire N__23845;
    wire N__23842;
    wire N__23839;
    wire N__23834;
    wire N__23831;
    wire N__23830;
    wire N__23829;
    wire N__23826;
    wire N__23823;
    wire N__23820;
    wire N__23815;
    wire N__23810;
    wire N__23807;
    wire N__23806;
    wire N__23803;
    wire N__23800;
    wire N__23797;
    wire N__23794;
    wire N__23791;
    wire N__23786;
    wire N__23783;
    wire N__23780;
    wire N__23779;
    wire N__23778;
    wire N__23775;
    wire N__23772;
    wire N__23769;
    wire N__23762;
    wire N__23759;
    wire N__23756;
    wire N__23755;
    wire N__23754;
    wire N__23753;
    wire N__23750;
    wire N__23743;
    wire N__23738;
    wire N__23735;
    wire N__23734;
    wire N__23731;
    wire N__23728;
    wire N__23725;
    wire N__23722;
    wire N__23719;
    wire N__23714;
    wire N__23711;
    wire N__23710;
    wire N__23709;
    wire N__23708;
    wire N__23705;
    wire N__23700;
    wire N__23697;
    wire N__23692;
    wire N__23687;
    wire N__23684;
    wire N__23683;
    wire N__23680;
    wire N__23679;
    wire N__23678;
    wire N__23677;
    wire N__23676;
    wire N__23675;
    wire N__23674;
    wire N__23673;
    wire N__23672;
    wire N__23671;
    wire N__23668;
    wire N__23665;
    wire N__23662;
    wire N__23659;
    wire N__23656;
    wire N__23653;
    wire N__23650;
    wire N__23649;
    wire N__23648;
    wire N__23645;
    wire N__23642;
    wire N__23641;
    wire N__23638;
    wire N__23637;
    wire N__23636;
    wire N__23635;
    wire N__23632;
    wire N__23631;
    wire N__23628;
    wire N__23623;
    wire N__23616;
    wire N__23613;
    wire N__23610;
    wire N__23607;
    wire N__23604;
    wire N__23601;
    wire N__23598;
    wire N__23595;
    wire N__23592;
    wire N__23589;
    wire N__23586;
    wire N__23585;
    wire N__23582;
    wire N__23579;
    wire N__23578;
    wire N__23573;
    wire N__23566;
    wire N__23563;
    wire N__23560;
    wire N__23555;
    wire N__23552;
    wire N__23545;
    wire N__23542;
    wire N__23537;
    wire N__23534;
    wire N__23531;
    wire N__23526;
    wire N__23517;
    wire N__23514;
    wire N__23509;
    wire N__23498;
    wire N__23497;
    wire N__23494;
    wire N__23493;
    wire N__23490;
    wire N__23489;
    wire N__23486;
    wire N__23483;
    wire N__23480;
    wire N__23477;
    wire N__23468;
    wire N__23465;
    wire N__23462;
    wire N__23461;
    wire N__23458;
    wire N__23455;
    wire N__23452;
    wire N__23449;
    wire N__23446;
    wire N__23441;
    wire N__23438;
    wire N__23435;
    wire N__23432;
    wire N__23429;
    wire N__23426;
    wire N__23423;
    wire N__23420;
    wire N__23417;
    wire N__23414;
    wire N__23411;
    wire N__23408;
    wire N__23405;
    wire N__23402;
    wire N__23399;
    wire N__23396;
    wire N__23393;
    wire N__23390;
    wire N__23387;
    wire N__23384;
    wire N__23381;
    wire N__23378;
    wire N__23375;
    wire N__23372;
    wire N__23369;
    wire N__23366;
    wire N__23363;
    wire N__23360;
    wire N__23357;
    wire N__23354;
    wire N__23351;
    wire N__23348;
    wire N__23345;
    wire N__23342;
    wire N__23339;
    wire N__23336;
    wire N__23333;
    wire N__23330;
    wire N__23327;
    wire N__23324;
    wire N__23321;
    wire N__23318;
    wire N__23315;
    wire N__23312;
    wire N__23309;
    wire N__23306;
    wire N__23303;
    wire N__23300;
    wire N__23297;
    wire N__23294;
    wire N__23291;
    wire N__23288;
    wire N__23285;
    wire N__23282;
    wire N__23279;
    wire N__23276;
    wire N__23273;
    wire N__23270;
    wire N__23267;
    wire N__23264;
    wire N__23261;
    wire N__23258;
    wire N__23255;
    wire N__23252;
    wire N__23249;
    wire N__23246;
    wire N__23243;
    wire N__23240;
    wire N__23237;
    wire N__23234;
    wire N__23231;
    wire N__23228;
    wire N__23225;
    wire N__23222;
    wire N__23219;
    wire N__23216;
    wire N__23213;
    wire N__23210;
    wire N__23207;
    wire N__23204;
    wire N__23201;
    wire N__23198;
    wire N__23195;
    wire N__23192;
    wire N__23189;
    wire N__23186;
    wire N__23183;
    wire N__23180;
    wire N__23177;
    wire N__23174;
    wire N__23171;
    wire N__23168;
    wire N__23165;
    wire N__23162;
    wire N__23159;
    wire N__23156;
    wire N__23153;
    wire N__23150;
    wire N__23147;
    wire N__23144;
    wire N__23141;
    wire N__23138;
    wire N__23135;
    wire N__23132;
    wire N__23129;
    wire N__23126;
    wire N__23123;
    wire N__23120;
    wire N__23117;
    wire N__23114;
    wire N__23111;
    wire N__23108;
    wire N__23105;
    wire N__23102;
    wire N__23099;
    wire N__23096;
    wire N__23093;
    wire N__23090;
    wire N__23087;
    wire N__23084;
    wire N__23081;
    wire N__23078;
    wire N__23075;
    wire N__23072;
    wire N__23069;
    wire N__23066;
    wire N__23063;
    wire N__23060;
    wire N__23057;
    wire N__23054;
    wire N__23051;
    wire N__23048;
    wire N__23045;
    wire N__23042;
    wire N__23039;
    wire N__23038;
    wire N__23037;
    wire N__23034;
    wire N__23031;
    wire N__23028;
    wire N__23027;
    wire N__23026;
    wire N__23021;
    wire N__23018;
    wire N__23015;
    wire N__23012;
    wire N__23005;
    wire N__23002;
    wire N__22999;
    wire N__22996;
    wire N__22993;
    wire N__22988;
    wire N__22985;
    wire N__22982;
    wire N__22979;
    wire N__22976;
    wire N__22973;
    wire N__22970;
    wire N__22967;
    wire N__22964;
    wire N__22961;
    wire N__22958;
    wire N__22955;
    wire N__22952;
    wire N__22949;
    wire N__22946;
    wire N__22943;
    wire N__22940;
    wire N__22937;
    wire N__22934;
    wire N__22931;
    wire N__22928;
    wire N__22925;
    wire N__22922;
    wire N__22919;
    wire N__22916;
    wire N__22913;
    wire N__22910;
    wire N__22907;
    wire N__22904;
    wire N__22901;
    wire N__22898;
    wire N__22895;
    wire N__22892;
    wire N__22889;
    wire N__22886;
    wire N__22883;
    wire N__22880;
    wire N__22877;
    wire N__22874;
    wire N__22871;
    wire N__22868;
    wire N__22865;
    wire N__22862;
    wire N__22859;
    wire N__22856;
    wire N__22853;
    wire N__22850;
    wire N__22847;
    wire N__22844;
    wire N__22841;
    wire N__22838;
    wire N__22835;
    wire N__22832;
    wire N__22829;
    wire N__22826;
    wire N__22823;
    wire N__22820;
    wire N__22817;
    wire N__22814;
    wire N__22811;
    wire N__22808;
    wire N__22805;
    wire N__22802;
    wire N__22799;
    wire N__22796;
    wire N__22793;
    wire N__22790;
    wire N__22787;
    wire N__22784;
    wire N__22781;
    wire N__22778;
    wire N__22775;
    wire N__22772;
    wire N__22769;
    wire N__22766;
    wire N__22763;
    wire N__22760;
    wire N__22757;
    wire N__22754;
    wire N__22751;
    wire N__22748;
    wire N__22745;
    wire N__22742;
    wire N__22741;
    wire N__22740;
    wire N__22739;
    wire N__22738;
    wire N__22737;
    wire N__22736;
    wire N__22735;
    wire N__22734;
    wire N__22733;
    wire N__22732;
    wire N__22727;
    wire N__22726;
    wire N__22725;
    wire N__22724;
    wire N__22723;
    wire N__22722;
    wire N__22721;
    wire N__22720;
    wire N__22719;
    wire N__22714;
    wire N__22699;
    wire N__22696;
    wire N__22691;
    wire N__22690;
    wire N__22689;
    wire N__22688;
    wire N__22687;
    wire N__22686;
    wire N__22685;
    wire N__22684;
    wire N__22683;
    wire N__22682;
    wire N__22669;
    wire N__22666;
    wire N__22663;
    wire N__22658;
    wire N__22653;
    wire N__22638;
    wire N__22625;
    wire N__22624;
    wire N__22623;
    wire N__22622;
    wire N__22621;
    wire N__22620;
    wire N__22619;
    wire N__22616;
    wire N__22615;
    wire N__22614;
    wire N__22613;
    wire N__22612;
    wire N__22611;
    wire N__22610;
    wire N__22609;
    wire N__22608;
    wire N__22605;
    wire N__22604;
    wire N__22601;
    wire N__22598;
    wire N__22595;
    wire N__22592;
    wire N__22591;
    wire N__22590;
    wire N__22589;
    wire N__22584;
    wire N__22581;
    wire N__22578;
    wire N__22577;
    wire N__22576;
    wire N__22575;
    wire N__22574;
    wire N__22571;
    wire N__22568;
    wire N__22565;
    wire N__22562;
    wire N__22559;
    wire N__22556;
    wire N__22555;
    wire N__22554;
    wire N__22553;
    wire N__22552;
    wire N__22551;
    wire N__22546;
    wire N__22531;
    wire N__22528;
    wire N__22523;
    wire N__22510;
    wire N__22495;
    wire N__22490;
    wire N__22487;
    wire N__22484;
    wire N__22479;
    wire N__22466;
    wire N__22465;
    wire N__22462;
    wire N__22459;
    wire N__22456;
    wire N__22453;
    wire N__22448;
    wire N__22447;
    wire N__22444;
    wire N__22441;
    wire N__22436;
    wire N__22433;
    wire N__22430;
    wire N__22427;
    wire N__22424;
    wire N__22421;
    wire N__22418;
    wire N__22415;
    wire N__22412;
    wire N__22409;
    wire N__22406;
    wire N__22403;
    wire N__22400;
    wire N__22397;
    wire N__22394;
    wire N__22391;
    wire N__22388;
    wire N__22385;
    wire N__22382;
    wire N__22379;
    wire N__22376;
    wire N__22373;
    wire N__22370;
    wire N__22367;
    wire N__22364;
    wire N__22361;
    wire N__22358;
    wire N__22355;
    wire N__22352;
    wire N__22349;
    wire N__22346;
    wire N__22343;
    wire N__22340;
    wire N__22337;
    wire N__22334;
    wire N__22331;
    wire N__22328;
    wire N__22325;
    wire N__22322;
    wire N__22319;
    wire N__22316;
    wire N__22313;
    wire N__22310;
    wire N__22307;
    wire N__22304;
    wire N__22301;
    wire N__22298;
    wire N__22295;
    wire N__22292;
    wire N__22289;
    wire N__22286;
    wire N__22283;
    wire N__22280;
    wire N__22277;
    wire N__22274;
    wire N__22271;
    wire N__22268;
    wire N__22265;
    wire N__22262;
    wire N__22259;
    wire N__22256;
    wire N__22253;
    wire N__22250;
    wire N__22247;
    wire N__22244;
    wire N__22241;
    wire N__22238;
    wire N__22235;
    wire N__22232;
    wire N__22229;
    wire N__22226;
    wire N__22223;
    wire N__22220;
    wire N__22217;
    wire N__22214;
    wire N__22211;
    wire N__22208;
    wire N__22205;
    wire N__22202;
    wire N__22199;
    wire N__22196;
    wire N__22193;
    wire N__22190;
    wire N__22187;
    wire N__22184;
    wire N__22181;
    wire N__22178;
    wire N__22175;
    wire N__22172;
    wire N__22169;
    wire N__22166;
    wire N__22163;
    wire N__22160;
    wire N__22157;
    wire N__22154;
    wire N__22151;
    wire N__22148;
    wire N__22145;
    wire N__22142;
    wire N__22139;
    wire N__22136;
    wire N__22133;
    wire N__22130;
    wire N__22127;
    wire N__22124;
    wire N__22121;
    wire N__22118;
    wire N__22115;
    wire N__22112;
    wire N__22109;
    wire N__22106;
    wire N__22103;
    wire N__22100;
    wire N__22097;
    wire N__22094;
    wire N__22091;
    wire N__22088;
    wire N__22085;
    wire N__22082;
    wire N__22079;
    wire N__22076;
    wire N__22073;
    wire N__22070;
    wire N__22067;
    wire N__22064;
    wire N__22061;
    wire N__22058;
    wire N__22055;
    wire N__22052;
    wire N__22049;
    wire N__22046;
    wire N__22043;
    wire N__22040;
    wire N__22037;
    wire N__22034;
    wire N__22033;
    wire N__22028;
    wire N__22025;
    wire N__22022;
    wire N__22019;
    wire N__22018;
    wire N__22015;
    wire N__22012;
    wire N__22007;
    wire N__22004;
    wire N__22001;
    wire N__21998;
    wire N__21995;
    wire N__21992;
    wire N__21989;
    wire N__21988;
    wire N__21985;
    wire N__21982;
    wire N__21977;
    wire N__21974;
    wire N__21971;
    wire N__21968;
    wire N__21965;
    wire N__21962;
    wire N__21959;
    wire N__21956;
    wire N__21953;
    wire N__21950;
    wire N__21947;
    wire N__21944;
    wire N__21941;
    wire N__21938;
    wire N__21935;
    wire N__21932;
    wire N__21929;
    wire N__21926;
    wire N__21923;
    wire N__21920;
    wire N__21917;
    wire N__21914;
    wire N__21911;
    wire N__21908;
    wire N__21907;
    wire N__21906;
    wire N__21905;
    wire N__21904;
    wire N__21901;
    wire N__21900;
    wire N__21897;
    wire N__21896;
    wire N__21893;
    wire N__21878;
    wire N__21875;
    wire N__21872;
    wire N__21871;
    wire N__21870;
    wire N__21869;
    wire N__21866;
    wire N__21859;
    wire N__21854;
    wire N__21851;
    wire N__21848;
    wire N__21845;
    wire N__21842;
    wire N__21839;
    wire N__21836;
    wire N__21833;
    wire N__21830;
    wire N__21827;
    wire N__21824;
    wire N__21821;
    wire N__21818;
    wire N__21815;
    wire N__21812;
    wire N__21809;
    wire N__21806;
    wire N__21803;
    wire N__21800;
    wire N__21797;
    wire N__21794;
    wire N__21791;
    wire N__21788;
    wire N__21785;
    wire N__21782;
    wire N__21779;
    wire N__21776;
    wire N__21773;
    wire N__21770;
    wire N__21767;
    wire N__21764;
    wire N__21761;
    wire N__21758;
    wire N__21755;
    wire N__21752;
    wire N__21749;
    wire N__21746;
    wire N__21743;
    wire N__21740;
    wire N__21737;
    wire N__21734;
    wire N__21731;
    wire N__21728;
    wire N__21725;
    wire N__21722;
    wire N__21719;
    wire N__21716;
    wire N__21715;
    wire N__21714;
    wire N__21713;
    wire N__21712;
    wire N__21711;
    wire N__21708;
    wire N__21705;
    wire N__21702;
    wire N__21697;
    wire N__21694;
    wire N__21685;
    wire N__21680;
    wire N__21677;
    wire N__21674;
    wire N__21671;
    wire N__21668;
    wire N__21667;
    wire N__21666;
    wire N__21665;
    wire N__21662;
    wire N__21659;
    wire N__21656;
    wire N__21655;
    wire N__21652;
    wire N__21649;
    wire N__21646;
    wire N__21643;
    wire N__21638;
    wire N__21629;
    wire N__21628;
    wire N__21625;
    wire N__21622;
    wire N__21621;
    wire N__21620;
    wire N__21619;
    wire N__21616;
    wire N__21613;
    wire N__21608;
    wire N__21605;
    wire N__21598;
    wire N__21593;
    wire N__21592;
    wire N__21589;
    wire N__21586;
    wire N__21581;
    wire N__21578;
    wire N__21575;
    wire N__21572;
    wire N__21569;
    wire N__21566;
    wire N__21563;
    wire N__21560;
    wire N__21557;
    wire N__21554;
    wire N__21551;
    wire N__21548;
    wire N__21545;
    wire N__21542;
    wire N__21539;
    wire N__21536;
    wire N__21533;
    wire N__21530;
    wire N__21527;
    wire N__21524;
    wire N__21521;
    wire N__21518;
    wire N__21515;
    wire N__21512;
    wire N__21509;
    wire N__21506;
    wire N__21503;
    wire N__21500;
    wire N__21497;
    wire N__21494;
    wire N__21491;
    wire N__21488;
    wire N__21485;
    wire N__21482;
    wire N__21479;
    wire N__21478;
    wire N__21475;
    wire N__21472;
    wire N__21467;
    wire N__21466;
    wire N__21465;
    wire N__21462;
    wire N__21459;
    wire N__21456;
    wire N__21453;
    wire N__21448;
    wire N__21443;
    wire N__21442;
    wire N__21439;
    wire N__21436;
    wire N__21431;
    wire N__21428;
    wire N__21427;
    wire N__21426;
    wire N__21425;
    wire N__21422;
    wire N__21417;
    wire N__21414;
    wire N__21411;
    wire N__21404;
    wire N__21401;
    wire N__21398;
    wire N__21395;
    wire N__21392;
    wire N__21389;
    wire N__21388;
    wire N__21385;
    wire N__21382;
    wire N__21377;
    wire N__21374;
    wire N__21371;
    wire N__21370;
    wire N__21365;
    wire N__21362;
    wire N__21359;
    wire N__21358;
    wire N__21355;
    wire N__21352;
    wire N__21349;
    wire N__21346;
    wire N__21343;
    wire N__21338;
    wire N__21335;
    wire N__21334;
    wire N__21331;
    wire N__21328;
    wire N__21323;
    wire N__21320;
    wire N__21319;
    wire N__21316;
    wire N__21313;
    wire N__21308;
    wire N__21305;
    wire N__21304;
    wire N__21301;
    wire N__21298;
    wire N__21293;
    wire N__21290;
    wire N__21289;
    wire N__21286;
    wire N__21283;
    wire N__21280;
    wire N__21275;
    wire N__21272;
    wire N__21269;
    wire N__21268;
    wire N__21267;
    wire N__21266;
    wire N__21265;
    wire N__21262;
    wire N__21259;
    wire N__21258;
    wire N__21257;
    wire N__21254;
    wire N__21253;
    wire N__21250;
    wire N__21247;
    wire N__21246;
    wire N__21245;
    wire N__21242;
    wire N__21237;
    wire N__21226;
    wire N__21223;
    wire N__21220;
    wire N__21217;
    wire N__21214;
    wire N__21207;
    wire N__21204;
    wire N__21201;
    wire N__21198;
    wire N__21195;
    wire N__21192;
    wire N__21185;
    wire N__21182;
    wire N__21179;
    wire N__21178;
    wire N__21173;
    wire N__21170;
    wire N__21167;
    wire N__21166;
    wire N__21161;
    wire N__21158;
    wire N__21155;
    wire N__21154;
    wire N__21151;
    wire N__21146;
    wire N__21143;
    wire N__21140;
    wire N__21137;
    wire N__21136;
    wire N__21133;
    wire N__21130;
    wire N__21125;
    wire N__21122;
    wire N__21121;
    wire N__21118;
    wire N__21115;
    wire N__21110;
    wire N__21107;
    wire N__21106;
    wire N__21101;
    wire N__21098;
    wire N__21095;
    wire N__21094;
    wire N__21091;
    wire N__21088;
    wire N__21083;
    wire N__21080;
    wire N__21077;
    wire N__21074;
    wire N__21073;
    wire N__21068;
    wire N__21065;
    wire N__21062;
    wire N__21061;
    wire N__21058;
    wire N__21057;
    wire N__21054;
    wire N__21051;
    wire N__21048;
    wire N__21045;
    wire N__21042;
    wire N__21037;
    wire N__21032;
    wire N__21029;
    wire N__21026;
    wire N__21025;
    wire N__21024;
    wire N__21021;
    wire N__21018;
    wire N__21015;
    wire N__21012;
    wire N__21009;
    wire N__21006;
    wire N__21001;
    wire N__20998;
    wire N__20995;
    wire N__20990;
    wire N__20987;
    wire N__20984;
    wire N__20981;
    wire N__20980;
    wire N__20977;
    wire N__20976;
    wire N__20973;
    wire N__20970;
    wire N__20967;
    wire N__20964;
    wire N__20961;
    wire N__20956;
    wire N__20951;
    wire N__20948;
    wire N__20947;
    wire N__20942;
    wire N__20939;
    wire N__20936;
    wire N__20935;
    wire N__20930;
    wire N__20927;
    wire N__20924;
    wire N__20921;
    wire N__20920;
    wire N__20917;
    wire N__20914;
    wire N__20909;
    wire N__20906;
    wire N__20905;
    wire N__20900;
    wire N__20897;
    wire N__20894;
    wire N__20891;
    wire N__20888;
    wire N__20887;
    wire N__20884;
    wire N__20881;
    wire N__20876;
    wire N__20873;
    wire N__20872;
    wire N__20869;
    wire N__20866;
    wire N__20861;
    wire N__20860;
    wire N__20859;
    wire N__20858;
    wire N__20857;
    wire N__20856;
    wire N__20855;
    wire N__20854;
    wire N__20851;
    wire N__20848;
    wire N__20847;
    wire N__20846;
    wire N__20843;
    wire N__20840;
    wire N__20833;
    wire N__20830;
    wire N__20825;
    wire N__20820;
    wire N__20815;
    wire N__20812;
    wire N__20811;
    wire N__20808;
    wire N__20803;
    wire N__20798;
    wire N__20795;
    wire N__20792;
    wire N__20789;
    wire N__20784;
    wire N__20777;
    wire N__20776;
    wire N__20775;
    wire N__20774;
    wire N__20773;
    wire N__20772;
    wire N__20771;
    wire N__20770;
    wire N__20769;
    wire N__20768;
    wire N__20763;
    wire N__20754;
    wire N__20747;
    wire N__20744;
    wire N__20737;
    wire N__20734;
    wire N__20731;
    wire N__20726;
    wire N__20725;
    wire N__20724;
    wire N__20723;
    wire N__20722;
    wire N__20721;
    wire N__20720;
    wire N__20719;
    wire N__20716;
    wire N__20713;
    wire N__20712;
    wire N__20709;
    wire N__20706;
    wire N__20703;
    wire N__20702;
    wire N__20697;
    wire N__20688;
    wire N__20685;
    wire N__20680;
    wire N__20677;
    wire N__20668;
    wire N__20665;
    wire N__20662;
    wire N__20657;
    wire N__20654;
    wire N__20651;
    wire N__20648;
    wire N__20645;
    wire N__20642;
    wire N__20639;
    wire N__20636;
    wire N__20633;
    wire N__20630;
    wire N__20627;
    wire N__20624;
    wire N__20621;
    wire N__20618;
    wire N__20615;
    wire N__20612;
    wire N__20609;
    wire N__20606;
    wire N__20603;
    wire N__20600;
    wire N__20597;
    wire N__20594;
    wire N__20591;
    wire N__20590;
    wire N__20587;
    wire N__20584;
    wire N__20583;
    wire N__20580;
    wire N__20577;
    wire N__20574;
    wire N__20569;
    wire N__20566;
    wire N__20563;
    wire N__20560;
    wire N__20555;
    wire N__20552;
    wire N__20549;
    wire N__20548;
    wire N__20545;
    wire N__20542;
    wire N__20541;
    wire N__20540;
    wire N__20537;
    wire N__20534;
    wire N__20531;
    wire N__20528;
    wire N__20523;
    wire N__20520;
    wire N__20517;
    wire N__20514;
    wire N__20509;
    wire N__20504;
    wire N__20501;
    wire N__20498;
    wire N__20495;
    wire N__20494;
    wire N__20493;
    wire N__20490;
    wire N__20487;
    wire N__20484;
    wire N__20477;
    wire N__20474;
    wire N__20471;
    wire N__20468;
    wire N__20467;
    wire N__20464;
    wire N__20463;
    wire N__20460;
    wire N__20457;
    wire N__20454;
    wire N__20451;
    wire N__20448;
    wire N__20443;
    wire N__20438;
    wire N__20435;
    wire N__20432;
    wire N__20431;
    wire N__20428;
    wire N__20425;
    wire N__20420;
    wire N__20417;
    wire N__20416;
    wire N__20413;
    wire N__20410;
    wire N__20405;
    wire N__20402;
    wire N__20399;
    wire N__20396;
    wire N__20393;
    wire N__20390;
    wire N__20387;
    wire N__20384;
    wire N__20381;
    wire N__20378;
    wire N__20375;
    wire N__20372;
    wire N__20369;
    wire N__20366;
    wire N__20363;
    wire N__20360;
    wire N__20357;
    wire N__20356;
    wire N__20353;
    wire N__20350;
    wire N__20345;
    wire N__20342;
    wire N__20341;
    wire N__20338;
    wire N__20335;
    wire N__20330;
    wire N__20327;
    wire N__20326;
    wire N__20323;
    wire N__20320;
    wire N__20315;
    wire N__20312;
    wire N__20311;
    wire N__20308;
    wire N__20305;
    wire N__20302;
    wire N__20297;
    wire N__20294;
    wire N__20291;
    wire N__20290;
    wire N__20287;
    wire N__20284;
    wire N__20281;
    wire N__20276;
    wire N__20273;
    wire N__20272;
    wire N__20269;
    wire N__20266;
    wire N__20261;
    wire N__20258;
    wire N__20255;
    wire N__20252;
    wire N__20249;
    wire N__20246;
    wire N__20243;
    wire N__20240;
    wire N__20237;
    wire N__20234;
    wire N__20231;
    wire N__20228;
    wire N__20225;
    wire N__20222;
    wire N__20219;
    wire N__20216;
    wire N__20213;
    wire N__20210;
    wire N__20207;
    wire N__20204;
    wire N__20201;
    wire N__20198;
    wire N__20197;
    wire N__20194;
    wire N__20191;
    wire N__20186;
    wire N__20183;
    wire N__20182;
    wire N__20179;
    wire N__20178;
    wire N__20175;
    wire N__20172;
    wire N__20169;
    wire N__20162;
    wire N__20159;
    wire N__20156;
    wire N__20153;
    wire N__20150;
    wire N__20149;
    wire N__20146;
    wire N__20143;
    wire N__20140;
    wire N__20139;
    wire N__20138;
    wire N__20137;
    wire N__20136;
    wire N__20135;
    wire N__20134;
    wire N__20133;
    wire N__20132;
    wire N__20127;
    wire N__20122;
    wire N__20111;
    wire N__20108;
    wire N__20105;
    wire N__20102;
    wire N__20101;
    wire N__20098;
    wire N__20095;
    wire N__20094;
    wire N__20091;
    wire N__20088;
    wire N__20085;
    wire N__20080;
    wire N__20077;
    wire N__20066;
    wire N__20063;
    wire N__20060;
    wire N__20057;
    wire N__20056;
    wire N__20055;
    wire N__20052;
    wire N__20049;
    wire N__20046;
    wire N__20043;
    wire N__20038;
    wire N__20035;
    wire N__20032;
    wire N__20027;
    wire N__20024;
    wire N__20021;
    wire N__20018;
    wire N__20015;
    wire N__20012;
    wire N__20009;
    wire N__20006;
    wire N__20005;
    wire N__20004;
    wire N__20003;
    wire N__20002;
    wire N__20001;
    wire N__20000;
    wire N__19997;
    wire N__19986;
    wire N__19983;
    wire N__19978;
    wire N__19975;
    wire N__19972;
    wire N__19969;
    wire N__19964;
    wire N__19961;
    wire N__19958;
    wire N__19955;
    wire N__19952;
    wire N__19949;
    wire N__19946;
    wire N__19943;
    wire N__19940;
    wire N__19937;
    wire N__19934;
    wire N__19931;
    wire N__19928;
    wire N__19925;
    wire N__19922;
    wire N__19919;
    wire N__19916;
    wire N__19913;
    wire N__19910;
    wire N__19907;
    wire N__19904;
    wire N__19901;
    wire N__19898;
    wire N__19895;
    wire N__19892;
    wire N__19889;
    wire N__19886;
    wire N__19883;
    wire N__19882;
    wire N__19879;
    wire N__19876;
    wire N__19873;
    wire N__19870;
    wire N__19865;
    wire N__19862;
    wire N__19859;
    wire N__19856;
    wire N__19853;
    wire N__19850;
    wire N__19847;
    wire N__19844;
    wire N__19841;
    wire N__19838;
    wire N__19835;
    wire N__19832;
    wire N__19829;
    wire N__19826;
    wire N__19823;
    wire N__19820;
    wire N__19817;
    wire N__19814;
    wire N__19811;
    wire N__19808;
    wire N__19805;
    wire N__19802;
    wire N__19799;
    wire N__19796;
    wire N__19795;
    wire N__19792;
    wire N__19789;
    wire N__19784;
    wire N__19781;
    wire N__19780;
    wire N__19779;
    wire N__19776;
    wire N__19773;
    wire N__19770;
    wire N__19767;
    wire N__19764;
    wire N__19757;
    wire N__19754;
    wire N__19751;
    wire N__19748;
    wire N__19745;
    wire N__19742;
    wire N__19739;
    wire N__19738;
    wire N__19737;
    wire N__19736;
    wire N__19727;
    wire N__19726;
    wire N__19723;
    wire N__19720;
    wire N__19715;
    wire N__19714;
    wire N__19713;
    wire N__19712;
    wire N__19709;
    wire N__19708;
    wire N__19705;
    wire N__19704;
    wire N__19703;
    wire N__19700;
    wire N__19697;
    wire N__19686;
    wire N__19685;
    wire N__19682;
    wire N__19681;
    wire N__19676;
    wire N__19673;
    wire N__19670;
    wire N__19667;
    wire N__19662;
    wire N__19659;
    wire N__19654;
    wire N__19649;
    wire N__19646;
    wire N__19643;
    wire N__19640;
    wire N__19637;
    wire N__19634;
    wire N__19631;
    wire N__19628;
    wire N__19627;
    wire N__19624;
    wire N__19621;
    wire N__19618;
    wire N__19613;
    wire N__19610;
    wire N__19609;
    wire N__19606;
    wire N__19603;
    wire N__19598;
    wire N__19595;
    wire N__19592;
    wire N__19589;
    wire N__19588;
    wire N__19585;
    wire N__19582;
    wire N__19577;
    wire N__19574;
    wire N__19571;
    wire N__19568;
    wire N__19567;
    wire N__19566;
    wire N__19563;
    wire N__19558;
    wire N__19553;
    wire N__19552;
    wire N__19549;
    wire N__19546;
    wire N__19543;
    wire N__19538;
    wire N__19537;
    wire N__19536;
    wire N__19533;
    wire N__19530;
    wire N__19527;
    wire N__19522;
    wire N__19517;
    wire N__19514;
    wire N__19511;
    wire N__19510;
    wire N__19507;
    wire N__19504;
    wire N__19501;
    wire N__19498;
    wire N__19493;
    wire N__19490;
    wire N__19489;
    wire N__19486;
    wire N__19485;
    wire N__19482;
    wire N__19479;
    wire N__19476;
    wire N__19469;
    wire N__19466;
    wire N__19463;
    wire N__19460;
    wire N__19457;
    wire N__19454;
    wire N__19451;
    wire N__19448;
    wire N__19445;
    wire N__19444;
    wire N__19443;
    wire N__19440;
    wire N__19437;
    wire N__19434;
    wire N__19427;
    wire N__19426;
    wire N__19423;
    wire N__19420;
    wire N__19415;
    wire N__19412;
    wire N__19409;
    wire N__19406;
    wire N__19403;
    wire N__19400;
    wire N__19399;
    wire N__19396;
    wire N__19393;
    wire N__19388;
    wire N__19387;
    wire N__19384;
    wire N__19381;
    wire N__19376;
    wire N__19373;
    wire N__19370;
    wire N__19367;
    wire N__19364;
    wire N__19361;
    wire N__19358;
    wire N__19355;
    wire N__19352;
    wire N__19349;
    wire N__19346;
    wire N__19343;
    wire N__19340;
    wire N__19337;
    wire N__19334;
    wire N__19331;
    wire N__19328;
    wire N__19325;
    wire N__19324;
    wire N__19321;
    wire N__19318;
    wire N__19315;
    wire N__19312;
    wire N__19307;
    wire N__19304;
    wire N__19301;
    wire N__19298;
    wire N__19295;
    wire N__19292;
    wire N__19289;
    wire N__19286;
    wire N__19283;
    wire N__19280;
    wire N__19277;
    wire N__19274;
    wire N__19271;
    wire N__19268;
    wire N__19265;
    wire N__19262;
    wire N__19259;
    wire N__19256;
    wire N__19253;
    wire N__19250;
    wire N__19247;
    wire N__19244;
    wire N__19241;
    wire N__19238;
    wire N__19235;
    wire N__19232;
    wire N__19229;
    wire N__19226;
    wire N__19223;
    wire N__19220;
    wire N__19217;
    wire N__19214;
    wire N__19211;
    wire N__19208;
    wire N__19205;
    wire N__19202;
    wire N__19199;
    wire N__19196;
    wire N__19193;
    wire N__19190;
    wire N__19187;
    wire N__19184;
    wire N__19181;
    wire N__19178;
    wire N__19175;
    wire N__19172;
    wire N__19169;
    wire N__19166;
    wire N__19163;
    wire N__19160;
    wire N__19157;
    wire N__19154;
    wire N__19151;
    wire N__19148;
    wire N__19145;
    wire N__19142;
    wire N__19139;
    wire N__19138;
    wire N__19137;
    wire N__19134;
    wire N__19129;
    wire N__19126;
    wire N__19121;
    wire N__19120;
    wire N__19117;
    wire N__19116;
    wire N__19113;
    wire N__19108;
    wire N__19105;
    wire N__19100;
    wire N__19099;
    wire N__19096;
    wire N__19095;
    wire N__19092;
    wire N__19089;
    wire N__19086;
    wire N__19083;
    wire N__19080;
    wire N__19073;
    wire N__19070;
    wire N__19067;
    wire N__19064;
    wire N__19063;
    wire N__19062;
    wire N__19059;
    wire N__19056;
    wire N__19053;
    wire N__19050;
    wire N__19043;
    wire N__19040;
    wire N__19037;
    wire N__19034;
    wire N__19031;
    wire N__19030;
    wire N__19027;
    wire N__19026;
    wire N__19019;
    wire N__19016;
    wire N__19015;
    wire N__19012;
    wire N__19009;
    wire N__19004;
    wire N__19003;
    wire N__19002;
    wire N__18999;
    wire N__18996;
    wire N__18993;
    wire N__18986;
    wire N__18983;
    wire N__18982;
    wire N__18979;
    wire N__18976;
    wire N__18971;
    wire N__18970;
    wire N__18967;
    wire N__18964;
    wire N__18959;
    wire N__18956;
    wire N__18953;
    wire N__18952;
    wire N__18951;
    wire N__18950;
    wire N__18949;
    wire N__18948;
    wire N__18947;
    wire N__18946;
    wire N__18945;
    wire N__18944;
    wire N__18943;
    wire N__18942;
    wire N__18941;
    wire N__18940;
    wire N__18939;
    wire N__18938;
    wire N__18937;
    wire N__18932;
    wire N__18915;
    wire N__18900;
    wire N__18897;
    wire N__18892;
    wire N__18891;
    wire N__18890;
    wire N__18889;
    wire N__18888;
    wire N__18887;
    wire N__18886;
    wire N__18885;
    wire N__18880;
    wire N__18875;
    wire N__18868;
    wire N__18863;
    wire N__18856;
    wire N__18851;
    wire N__18848;
    wire N__18847;
    wire N__18846;
    wire N__18843;
    wire N__18840;
    wire N__18837;
    wire N__18830;
    wire N__18827;
    wire N__18824;
    wire N__18821;
    wire N__18818;
    wire N__18815;
    wire N__18812;
    wire N__18809;
    wire N__18806;
    wire N__18803;
    wire N__18800;
    wire N__18797;
    wire N__18794;
    wire N__18791;
    wire N__18788;
    wire N__18785;
    wire N__18782;
    wire N__18779;
    wire N__18776;
    wire N__18773;
    wire N__18770;
    wire N__18767;
    wire N__18764;
    wire N__18761;
    wire N__18758;
    wire N__18755;
    wire N__18752;
    wire N__18749;
    wire N__18746;
    wire N__18743;
    wire N__18740;
    wire N__18737;
    wire N__18734;
    wire N__18731;
    wire N__18728;
    wire N__18725;
    wire N__18722;
    wire N__18719;
    wire N__18716;
    wire N__18713;
    wire N__18710;
    wire N__18707;
    wire N__18704;
    wire N__18701;
    wire N__18698;
    wire N__18695;
    wire N__18692;
    wire N__18689;
    wire N__18688;
    wire N__18687;
    wire N__18686;
    wire N__18685;
    wire N__18682;
    wire N__18681;
    wire N__18678;
    wire N__18677;
    wire N__18674;
    wire N__18673;
    wire N__18668;
    wire N__18655;
    wire N__18650;
    wire N__18647;
    wire N__18644;
    wire N__18641;
    wire N__18638;
    wire N__18635;
    wire N__18632;
    wire N__18629;
    wire N__18626;
    wire N__18623;
    wire N__18620;
    wire N__18617;
    wire N__18614;
    wire N__18611;
    wire N__18608;
    wire N__18605;
    wire N__18602;
    wire N__18599;
    wire N__18596;
    wire N__18593;
    wire N__18590;
    wire N__18587;
    wire N__18584;
    wire N__18581;
    wire N__18578;
    wire N__18575;
    wire N__18572;
    wire N__18569;
    wire N__18566;
    wire N__18563;
    wire N__18560;
    wire N__18557;
    wire N__18554;
    wire N__18551;
    wire N__18548;
    wire N__18545;
    wire N__18542;
    wire N__18539;
    wire N__18536;
    wire N__18533;
    wire N__18530;
    wire N__18527;
    wire N__18524;
    wire N__18521;
    wire N__18518;
    wire N__18515;
    wire N__18512;
    wire N__18509;
    wire N__18506;
    wire N__18503;
    wire N__18500;
    wire N__18497;
    wire N__18494;
    wire N__18491;
    wire N__18488;
    wire N__18485;
    wire N__18482;
    wire N__18479;
    wire N__18476;
    wire N__18473;
    wire N__18470;
    wire N__18467;
    wire N__18464;
    wire N__18461;
    wire N__18458;
    wire N__18455;
    wire N__18452;
    wire N__18449;
    wire N__18446;
    wire N__18443;
    wire N__18440;
    wire N__18437;
    wire N__18434;
    wire N__18431;
    wire N__18428;
    wire N__18425;
    wire N__18422;
    wire N__18419;
    wire N__18416;
    wire N__18413;
    wire N__18410;
    wire N__18407;
    wire N__18404;
    wire N__18401;
    wire N__18398;
    wire N__18395;
    wire N__18392;
    wire N__18389;
    wire N__18386;
    wire N__18383;
    wire N__18380;
    wire N__18377;
    wire N__18374;
    wire N__18371;
    wire N__18368;
    wire N__18365;
    wire N__18362;
    wire N__18359;
    wire N__18356;
    wire N__18353;
    wire N__18350;
    wire N__18347;
    wire N__18344;
    wire N__18341;
    wire N__18338;
    wire N__18335;
    wire N__18332;
    wire N__18329;
    wire N__18326;
    wire N__18323;
    wire N__18320;
    wire N__18319;
    wire N__18314;
    wire N__18311;
    wire N__18308;
    wire N__18305;
    wire N__18302;
    wire N__18299;
    wire N__18296;
    wire N__18293;
    wire N__18290;
    wire N__18287;
    wire N__18284;
    wire N__18281;
    wire N__18278;
    wire N__18275;
    wire N__18272;
    wire N__18269;
    wire N__18266;
    wire N__18263;
    wire N__18260;
    wire N__18257;
    wire N__18254;
    wire N__18251;
    wire N__18248;
    wire N__18245;
    wire N__18242;
    wire N__18239;
    wire N__18236;
    wire N__18233;
    wire N__18230;
    wire N__18227;
    wire N__18224;
    wire N__18221;
    wire N__18218;
    wire N__18215;
    wire N__18212;
    wire N__18209;
    wire N__18206;
    wire N__18203;
    wire N__18200;
    wire N__18197;
    wire N__18194;
    wire N__18191;
    wire N__18188;
    wire N__18185;
    wire N__18182;
    wire N__18179;
    wire N__18176;
    wire N__18173;
    wire N__18170;
    wire N__18167;
    wire N__18164;
    wire N__18161;
    wire N__18158;
    wire N__18155;
    wire N__18152;
    wire N__18149;
    wire N__18146;
    wire N__18145;
    wire N__18144;
    wire N__18137;
    wire N__18134;
    wire GNDG0;
    wire VCCG0;
    wire \current_shift_inst.PI_CTRL.N_97 ;
    wire bfn_1_9_0_;
    wire \pwm_generator_inst.O_12 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_0 ;
    wire \pwm_generator_inst.O_13 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_1 ;
    wire \pwm_generator_inst.O_14 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_2 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_3 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_4 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_5 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_6 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_7 ;
    wire bfn_1_10_0_;
    wire \pwm_generator_inst.un3_threshold_acc_cry_8 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_9 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_10 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_11 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_12 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_13 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_14 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_15 ;
    wire bfn_1_11_0_;
    wire \pwm_generator_inst.un3_threshold_acc_cry_16 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_17 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_18 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_19 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_1_16 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_1_15 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_0 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_15 ;
    wire \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4 ;
    wire bfn_1_12_0_;
    wire \pwm_generator_inst.un2_threshold_acc_1_16 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_1 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_17 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_2 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_18 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_3 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_19 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_4 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_20 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_5 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_21 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_6 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_22 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_7 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_7 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_23 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_8 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0 ;
    wire bfn_1_13_0_;
    wire \pwm_generator_inst.un2_threshold_acc_1_24 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_9 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_10 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_11 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_12 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_13 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_14 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_25 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_15 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO ;
    wire bfn_1_14_0_;
    wire N_110_i_i;
    wire un7_start_stop;
    wire pwm_duty_input_5;
    wire pwm_duty_input_9;
    wire pwm_duty_input_8;
    wire \current_shift_inst.PI_CTRL.m7_2 ;
    wire pwm_duty_input_7;
    wire \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_0_3 ;
    wire pwm_duty_input_1;
    wire pwm_duty_input_3;
    wire pwm_duty_input_0;
    wire pwm_duty_input_2;
    wire \current_shift_inst.PI_CTRL.m14_2 ;
    wire pwm_duty_input_10;
    wire \current_shift_inst.PI_CTRL.N_19_cascade_ ;
    wire pwm_duty_input_4;
    wire \pwm_generator_inst.O_0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_0 ;
    wire bfn_2_7_0_;
    wire \pwm_generator_inst.O_1 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_1 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_0 ;
    wire \pwm_generator_inst.O_2 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_2 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_1 ;
    wire \pwm_generator_inst.O_3 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_3 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_2 ;
    wire \pwm_generator_inst.O_4 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_4 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_3 ;
    wire \pwm_generator_inst.O_5 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_5 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_4 ;
    wire \pwm_generator_inst.O_6 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_6 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_5 ;
    wire \pwm_generator_inst.O_7 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_7 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_6 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_7 ;
    wire \pwm_generator_inst.O_8 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_8 ;
    wire bfn_2_8_0_;
    wire \pwm_generator_inst.O_9 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_9 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_8 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_9 ;
    wire \pwm_generator_inst.un3_threshold_acc ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_10 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_11 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_12 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_13 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_14 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_15 ;
    wire bfn_2_9_0_;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_16 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_17 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_18 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_15 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_17 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_ ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_18 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_18_cascade_ ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_16 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_13 ;
    wire \pwm_generator_inst.O_10 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_10 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_12 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.N_98_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_96 ;
    wire \current_shift_inst.PI_CTRL.N_178 ;
    wire \current_shift_inst.PI_CTRL.N_91 ;
    wire un2_counter_7_cascade_;
    wire \pwm_generator_inst.un19_threshold_acc_axb_0 ;
    wire bfn_3_9_0_;
    wire \pwm_generator_inst.un19_threshold_acc_axb_1 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_0 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_2 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_1 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_3 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_2 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_3 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_5 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_4 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_6 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_5 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_7 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_6 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_7 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_8 ;
    wire bfn_3_10_0_;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO ;
    wire \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_8 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9 ;
    wire \current_shift_inst.PI_CTRL.N_27 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_14 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_4 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_31 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_9_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_118 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ;
    wire bfn_4_7_0_;
    wire un5_counter_cry_1;
    wire counterZ0Z_3;
    wire un5_counter_cry_2;
    wire counterZ0Z_4;
    wire un5_counter_cry_3;
    wire counterZ0Z_5;
    wire un5_counter_cry_4;
    wire counterZ0Z_6;
    wire un5_counter_cry_5;
    wire un5_counter_cry_6;
    wire counterZ0Z_8;
    wire un5_counter_cry_7;
    wire un5_counter_cry_8;
    wire counterZ0Z_9;
    wire bfn_4_8_0_;
    wire un5_counter_cry_9;
    wire counterZ0Z_11;
    wire un5_counter_cry_10;
    wire counterZ0Z_12;
    wire un5_counter_cry_11;
    wire counter_RNO_0Z0Z_12;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5 ;
    wire pwm_duty_input_6;
    wire N_28_mux;
    wire i8_mux;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ;
    wire bfn_4_13_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto3 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto4 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ;
    wire bfn_4_14_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ;
    wire bfn_4_15_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ;
    wire bfn_4_16_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ;
    wire \current_shift_inst.PI_CTRL.un8_enablelto31 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_12 ;
    wire counter_RNO_0Z0Z_7;
    wire counterZ0Z_7;
    wire counterZ0Z_1;
    wire counterZ0Z_2;
    wire un2_counter_5_cascade_;
    wire counterZ0Z_0;
    wire un2_counter_9_cascade_;
    wire clk_10khz_RNIIENAZ0Z2_cascade_;
    wire \pwm_generator_inst.threshold_ACCZ0Z_2 ;
    wire un2_counter_8;
    wire counter_RNO_0Z0Z_10;
    wire un2_counter_9;
    wire un2_counter_7;
    wire counterZ0Z_10;
    wire \pwm_generator_inst.threshold_ACCZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_10_31_cascade_ ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_11_31 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_9_31 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_8_31 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_25 ;
    wire clk_10khz_i;
    wire clk_10khz_RNIIENAZ0Z2;
    wire \pwm_generator_inst.threshold_ACCZ0Z_7 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_1 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_4 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_3 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_2_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_2 ;
    wire \current_shift_inst.PI_CTRL.N_47_21 ;
    wire \current_shift_inst.PI_CTRL.N_43 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31_cascade_ ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31 ;
    wire \current_shift_inst.PI_CTRL.N_46_21 ;
    wire \current_shift_inst.PI_CTRL.N_46_21_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_44 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_7 ;
    wire bfn_7_17_0_;
    wire \current_shift_inst.control_input_1_cry_0 ;
    wire \current_shift_inst.control_input_1_cry_1 ;
    wire \current_shift_inst.control_input_1_cry_2 ;
    wire \current_shift_inst.control_input_1_cry_3 ;
    wire \current_shift_inst.control_input_1_cry_4 ;
    wire \current_shift_inst.control_input_1_cry_5 ;
    wire \current_shift_inst.control_input_1_cry_6 ;
    wire \current_shift_inst.control_input_1_cry_7 ;
    wire bfn_7_18_0_;
    wire \current_shift_inst.control_input_1_cry_8 ;
    wire \current_shift_inst.control_input_1_cry_9 ;
    wire \current_shift_inst.control_input_1_cry_10 ;
    wire \current_shift_inst.control_input_1_cry_11 ;
    wire \current_shift_inst.control_input_1_cry_12 ;
    wire \current_shift_inst.control_input_1_cry_13 ;
    wire \current_shift_inst.control_input_1_cry_14 ;
    wire \current_shift_inst.control_input_1_cry_15 ;
    wire bfn_7_19_0_;
    wire \current_shift_inst.control_input_1_cry_16 ;
    wire \current_shift_inst.control_input_1_cry_17 ;
    wire \current_shift_inst.control_input_1_cry_18 ;
    wire \current_shift_inst.control_input_1_cry_19 ;
    wire \current_shift_inst.control_input_1_cry_20 ;
    wire \current_shift_inst.control_input_1_cry_21 ;
    wire \current_shift_inst.control_input_1_cry_22 ;
    wire \current_shift_inst.control_input_1_cry_23 ;
    wire bfn_7_20_0_;
    wire \current_shift_inst.control_input_1_cry_24 ;
    wire il_min_comp2_c;
    wire il_max_comp2_c;
    wire \pwm_generator_inst.threshold_ACCZ0Z_0 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_6 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_3 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_5 ;
    wire bfn_8_11_0_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_1 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ1Z_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_8 ;
    wire bfn_8_12_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_9 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_16 ;
    wire bfn_8_13_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_17 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \current_shift_inst.PI_CTRL.un1_enablelt3_0 ;
    wire \current_shift_inst.PI_CTRL.N_47_16 ;
    wire \current_shift_inst.PI_CTRL.N_46_16 ;
    wire \current_shift_inst.PI_CTRL.N_76 ;
    wire \current_shift_inst.PI_CTRL.N_75 ;
    wire bfn_8_17_0_;
    wire \current_shift_inst.z_i_0_31 ;
    wire \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CO ;
    wire \current_shift_inst.un38_control_input_0_cry_0 ;
    wire \current_shift_inst.un38_control_input_0_cry_1 ;
    wire \current_shift_inst.un38_control_input_0_cry_3_c_invZ0 ;
    wire \current_shift_inst.un38_control_input_0_cry_2 ;
    wire \current_shift_inst.un38_control_input_0_cry_3 ;
    wire \current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0Z_0 ;
    wire \current_shift_inst.un38_control_input_0_cry_4 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIVQKU1_5 ;
    wire \current_shift_inst.control_input_1_axb_0 ;
    wire \current_shift_inst.un38_control_input_0_cry_5 ;
    wire \current_shift_inst.un38_control_input_0_cry_6 ;
    wire \current_shift_inst.control_input_1_axb_1 ;
    wire bfn_8_18_0_;
    wire \current_shift_inst.control_input_1_axb_2 ;
    wire \current_shift_inst.un38_control_input_0_cry_7 ;
    wire \current_shift_inst.control_input_1_axb_3 ;
    wire \current_shift_inst.un38_control_input_0_cry_8 ;
    wire \current_shift_inst.control_input_1_axb_4 ;
    wire \current_shift_inst.un38_control_input_0_cry_9 ;
    wire \current_shift_inst.control_input_1_axb_5 ;
    wire \current_shift_inst.un38_control_input_0_cry_10 ;
    wire \current_shift_inst.control_input_1_axb_6 ;
    wire \current_shift_inst.un38_control_input_0_cry_11 ;
    wire \current_shift_inst.control_input_1_axb_7 ;
    wire \current_shift_inst.un38_control_input_0_cry_12 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIR0UI_13 ;
    wire \current_shift_inst.control_input_1_axb_8 ;
    wire \current_shift_inst.un38_control_input_0_cry_13 ;
    wire \current_shift_inst.un38_control_input_0_cry_14 ;
    wire \current_shift_inst.control_input_1_axb_9 ;
    wire bfn_8_19_0_;
    wire \current_shift_inst.control_input_1_axb_10 ;
    wire \current_shift_inst.un38_control_input_0_cry_15 ;
    wire \current_shift_inst.control_input_1_axb_11 ;
    wire \current_shift_inst.un38_control_input_0_cry_16 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIH6661_17 ;
    wire \current_shift_inst.control_input_1_axb_12 ;
    wire \current_shift_inst.un38_control_input_0_cry_17 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIAL3J_18 ;
    wire \current_shift_inst.control_input_1_axb_13 ;
    wire \current_shift_inst.un38_control_input_0_cry_18 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI4H5J_19 ;
    wire \current_shift_inst.control_input_1_axb_14 ;
    wire \current_shift_inst.un38_control_input_0_cry_19 ;
    wire \current_shift_inst.control_input_1_axb_15 ;
    wire \current_shift_inst.un38_control_input_0_cry_20 ;
    wire \current_shift_inst.control_input_1_axb_16 ;
    wire \current_shift_inst.un38_control_input_0_cry_21 ;
    wire \current_shift_inst.un38_control_input_0_cry_22 ;
    wire \current_shift_inst.control_input_1_axb_17 ;
    wire bfn_8_20_0_;
    wire \current_shift_inst.control_input_1_axb_18 ;
    wire \current_shift_inst.un38_control_input_0_cry_23 ;
    wire \current_shift_inst.control_input_1_axb_19 ;
    wire \current_shift_inst.un38_control_input_0_cry_24 ;
    wire \current_shift_inst.control_input_1_axb_20 ;
    wire \current_shift_inst.un38_control_input_0_cry_25 ;
    wire \current_shift_inst.control_input_1_axb_21 ;
    wire \current_shift_inst.un38_control_input_0_cry_26 ;
    wire \current_shift_inst.control_input_1_axb_22 ;
    wire \current_shift_inst.un38_control_input_0_cry_27 ;
    wire \current_shift_inst.control_input_1_axb_23 ;
    wire \current_shift_inst.un38_control_input_0_cry_28 ;
    wire \current_shift_inst.control_input_1_axb_24 ;
    wire \current_shift_inst.un38_control_input_0_cry_29 ;
    wire \current_shift_inst.un38_control_input_0_cry_30 ;
    wire \current_shift_inst.control_input_1_cry_24_THRU_CO ;
    wire bfn_8_21_0_;
    wire \current_shift_inst.phase_valid_RNISLORZ0Z2 ;
    wire il_min_comp2_D1;
    wire il_max_comp1_c;
    wire \pwm_generator_inst.thresholdZ0Z_0 ;
    wire \pwm_generator_inst.counter_i_0 ;
    wire bfn_9_8_0_;
    wire \pwm_generator_inst.thresholdZ0Z_1 ;
    wire \pwm_generator_inst.counter_i_1 ;
    wire \pwm_generator_inst.un14_counter_cry_0 ;
    wire \pwm_generator_inst.thresholdZ0Z_2 ;
    wire \pwm_generator_inst.counter_i_2 ;
    wire \pwm_generator_inst.un14_counter_cry_1 ;
    wire \pwm_generator_inst.thresholdZ0Z_3 ;
    wire \pwm_generator_inst.counter_i_3 ;
    wire \pwm_generator_inst.un14_counter_cry_2 ;
    wire \pwm_generator_inst.thresholdZ0Z_4 ;
    wire \pwm_generator_inst.counter_i_4 ;
    wire \pwm_generator_inst.un14_counter_cry_3 ;
    wire \pwm_generator_inst.thresholdZ0Z_5 ;
    wire \pwm_generator_inst.counter_i_5 ;
    wire \pwm_generator_inst.un14_counter_cry_4 ;
    wire \pwm_generator_inst.thresholdZ0Z_6 ;
    wire \pwm_generator_inst.counter_i_6 ;
    wire \pwm_generator_inst.un14_counter_cry_5 ;
    wire \pwm_generator_inst.thresholdZ0Z_7 ;
    wire \pwm_generator_inst.counter_i_7 ;
    wire \pwm_generator_inst.un14_counter_cry_6 ;
    wire \pwm_generator_inst.un14_counter_cry_7 ;
    wire \pwm_generator_inst.thresholdZ0Z_8 ;
    wire \pwm_generator_inst.counter_i_8 ;
    wire bfn_9_9_0_;
    wire \pwm_generator_inst.thresholdZ0Z_9 ;
    wire \pwm_generator_inst.counter_i_9 ;
    wire \pwm_generator_inst.un14_counter_cry_8 ;
    wire \pwm_generator_inst.un14_counter_cry_9 ;
    wire pwm_output_c;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_0 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0 ;
    wire \current_shift_inst.control_inputZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_0 ;
    wire bfn_9_13_0_;
    wire \current_shift_inst.control_inputZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_0 ;
    wire \current_shift_inst.control_inputZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_1 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0 ;
    wire \current_shift_inst.control_inputZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_2 ;
    wire N_702_g;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_4 ;
    wire \current_shift_inst.control_inputZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_3 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_5 ;
    wire \current_shift_inst.control_inputZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_4 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_6 ;
    wire \current_shift_inst.control_inputZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_5 ;
    wire \current_shift_inst.control_inputZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_6 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_7 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_8 ;
    wire \current_shift_inst.control_inputZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ;
    wire bfn_9_14_0_;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_9 ;
    wire \current_shift_inst.control_inputZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_8 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_10 ;
    wire \current_shift_inst.control_inputZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_9 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_11 ;
    wire \current_shift_inst.control_inputZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_10 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_12 ;
    wire \current_shift_inst.control_inputZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_11 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_13 ;
    wire \current_shift_inst.control_inputZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_12 ;
    wire \current_shift_inst.control_inputZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_13 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_15 ;
    wire \current_shift_inst.control_inputZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_14 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_15 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_16 ;
    wire \current_shift_inst.control_inputZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ;
    wire bfn_9_15_0_;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_17 ;
    wire \current_shift_inst.control_inputZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_18 ;
    wire \current_shift_inst.control_inputZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_19 ;
    wire \current_shift_inst.control_inputZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_18 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_20 ;
    wire \current_shift_inst.control_inputZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_21 ;
    wire \current_shift_inst.control_inputZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_22 ;
    wire \current_shift_inst.control_inputZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_21 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_23 ;
    wire \current_shift_inst.control_inputZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_22 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_23 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_24 ;
    wire \current_shift_inst.control_inputZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ;
    wire bfn_9_16_0_;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_25 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_29 ;
    wire \current_shift_inst.control_inputZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_31 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ;
    wire \current_shift_inst.un38_control_input_0_cry_1_c_RNOZ0 ;
    wire \current_shift_inst.N_1717_i ;
    wire \current_shift_inst.un38_control_input_0_cry_2_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3_cascade_ ;
    wire \current_shift_inst.un38_control_input_0_cry_4_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIK3CV_7 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIP5T51_13 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIER9V_5 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJDBL1_10 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIE6961_18 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIHVAV_6 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI7DM51_10 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI53NU1_6 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI7H2J_17 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIIKQI_10 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIU4VI_14 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIBU361_16 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIBBPU1_7 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI1PG21_9 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNINKG81_27 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIR32K_22 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPB581_22 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJ3381_21 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIVQF91_30 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIAO7K_27 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI4D1J_16 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIKKJ81_29 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIHCE81_26 ;
    wire bfn_9_21_0_;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_2 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_3 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_4 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_5 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_6 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_7 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_8 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_9 ;
    wire bfn_9_22_0_;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_10 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_11 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_12 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_13 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_14 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_15 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_16 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_17 ;
    wire bfn_9_23_0_;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_18 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_19 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_20 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_21 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_22 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_23 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_24 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_25 ;
    wire bfn_9_24_0_;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_26 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_27 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_28 ;
    wire \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_29 ;
    wire \current_shift_inst.timer_phase.N_188_i_g ;
    wire \current_shift_inst.timer_phase.counterZ0Z_0 ;
    wire bfn_9_25_0_;
    wire \current_shift_inst.timer_phase.counterZ0Z_1 ;
    wire \current_shift_inst.timer_phase.counter_cry_0 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_2 ;
    wire \current_shift_inst.timer_phase.counter_cry_1 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_3 ;
    wire \current_shift_inst.timer_phase.counter_cry_2 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_4 ;
    wire \current_shift_inst.timer_phase.counter_cry_3 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_5 ;
    wire \current_shift_inst.timer_phase.counter_cry_4 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_6 ;
    wire \current_shift_inst.timer_phase.counter_cry_5 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_7 ;
    wire \current_shift_inst.timer_phase.counter_cry_6 ;
    wire \current_shift_inst.timer_phase.counter_cry_7 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_8 ;
    wire bfn_9_26_0_;
    wire \current_shift_inst.timer_phase.counterZ0Z_9 ;
    wire \current_shift_inst.timer_phase.counter_cry_8 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_10 ;
    wire \current_shift_inst.timer_phase.counter_cry_9 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_11 ;
    wire \current_shift_inst.timer_phase.counter_cry_10 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_12 ;
    wire \current_shift_inst.timer_phase.counter_cry_11 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_13 ;
    wire \current_shift_inst.timer_phase.counter_cry_12 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_14 ;
    wire \current_shift_inst.timer_phase.counter_cry_13 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_15 ;
    wire \current_shift_inst.timer_phase.counter_cry_14 ;
    wire \current_shift_inst.timer_phase.counter_cry_15 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_16 ;
    wire bfn_9_27_0_;
    wire \current_shift_inst.timer_phase.counterZ0Z_17 ;
    wire \current_shift_inst.timer_phase.counter_cry_16 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_18 ;
    wire \current_shift_inst.timer_phase.counter_cry_17 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_19 ;
    wire \current_shift_inst.timer_phase.counter_cry_18 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_20 ;
    wire \current_shift_inst.timer_phase.counter_cry_19 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_21 ;
    wire \current_shift_inst.timer_phase.counter_cry_20 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_22 ;
    wire \current_shift_inst.timer_phase.counter_cry_21 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_23 ;
    wire \current_shift_inst.timer_phase.counter_cry_22 ;
    wire \current_shift_inst.timer_phase.counter_cry_23 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_24 ;
    wire bfn_9_28_0_;
    wire \current_shift_inst.timer_phase.counterZ0Z_25 ;
    wire \current_shift_inst.timer_phase.counter_cry_24 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_26 ;
    wire \current_shift_inst.timer_phase.counter_cry_25 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_27 ;
    wire \current_shift_inst.timer_phase.counter_cry_26 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_28 ;
    wire \current_shift_inst.timer_phase.counter_cry_27 ;
    wire \current_shift_inst.timer_phase.counter_cry_28 ;
    wire \current_shift_inst.timer_phase.counterZ0Z_29 ;
    wire il_max_comp1_D1;
    wire \pwm_generator_inst.un1_counterlto2_0_cascade_ ;
    wire \pwm_generator_inst.un1_counterlt9_cascade_ ;
    wire \pwm_generator_inst.un1_counterlto9_2 ;
    wire \pwm_generator_inst.counterZ0Z_0 ;
    wire bfn_10_9_0_;
    wire \pwm_generator_inst.counterZ0Z_1 ;
    wire \pwm_generator_inst.counter_cry_0 ;
    wire \pwm_generator_inst.counterZ0Z_2 ;
    wire \pwm_generator_inst.counter_cry_1 ;
    wire \pwm_generator_inst.counterZ0Z_3 ;
    wire \pwm_generator_inst.counter_cry_2 ;
    wire \pwm_generator_inst.counterZ0Z_4 ;
    wire \pwm_generator_inst.counter_cry_3 ;
    wire \pwm_generator_inst.counterZ0Z_5 ;
    wire \pwm_generator_inst.counter_cry_4 ;
    wire \pwm_generator_inst.counterZ0Z_6 ;
    wire \pwm_generator_inst.counter_cry_5 ;
    wire \pwm_generator_inst.counterZ0Z_7 ;
    wire \pwm_generator_inst.counter_cry_6 ;
    wire \pwm_generator_inst.counter_cry_7 ;
    wire \pwm_generator_inst.counterZ0Z_8 ;
    wire bfn_10_10_0_;
    wire \pwm_generator_inst.un1_counter_0 ;
    wire \pwm_generator_inst.counter_cry_8 ;
    wire \pwm_generator_inst.counterZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.time_passed11 ;
    wire \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa ;
    wire G_407;
    wire bfn_10_14_0_;
    wire G_406;
    wire \current_shift_inst.z_cry_0 ;
    wire \current_shift_inst.z_cry_1 ;
    wire \current_shift_inst.z_cry_2 ;
    wire \current_shift_inst.z_cry_3 ;
    wire \current_shift_inst.z_cry_4 ;
    wire \current_shift_inst.z_cry_5 ;
    wire \current_shift_inst.z_cry_6 ;
    wire \current_shift_inst.z_cry_7 ;
    wire bfn_10_15_0_;
    wire \current_shift_inst.z_cry_8 ;
    wire \current_shift_inst.z_cry_9 ;
    wire \current_shift_inst.z_cry_10 ;
    wire \current_shift_inst.z_cry_11 ;
    wire \current_shift_inst.z_cry_12 ;
    wire \current_shift_inst.z_cry_13 ;
    wire \current_shift_inst.z_cry_14 ;
    wire \current_shift_inst.z_cry_15 ;
    wire bfn_10_16_0_;
    wire \current_shift_inst.z_cry_16 ;
    wire \current_shift_inst.z_cry_17 ;
    wire \current_shift_inst.z_cry_18 ;
    wire \current_shift_inst.z_cry_19 ;
    wire \current_shift_inst.z_cry_20 ;
    wire \current_shift_inst.z_cry_21 ;
    wire \current_shift_inst.z_cry_22 ;
    wire \current_shift_inst.z_cry_23 ;
    wire bfn_10_17_0_;
    wire \current_shift_inst.z_cry_24 ;
    wire \current_shift_inst.z_cry_25 ;
    wire \current_shift_inst.z_cry_26 ;
    wire \current_shift_inst.z_cry_27 ;
    wire \current_shift_inst.z_cry_28 ;
    wire \current_shift_inst.z_cry_29 ;
    wire \current_shift_inst.z_cry_30 ;
    wire \current_shift_inst.elapsed_time_ns_phase_1 ;
    wire bfn_10_18_0_;
    wire \current_shift_inst.elapsed_time_ns_phase_2 ;
    wire \current_shift_inst.z_5_2 ;
    wire \current_shift_inst.z_5_cry_1 ;
    wire \current_shift_inst.elapsed_time_ns_phase_3 ;
    wire \current_shift_inst.z_5_3 ;
    wire \current_shift_inst.z_5_cry_2 ;
    wire \current_shift_inst.elapsed_time_ns_phase_4 ;
    wire \current_shift_inst.z_5_4 ;
    wire \current_shift_inst.z_5_cry_3 ;
    wire \current_shift_inst.elapsed_time_ns_phase_5 ;
    wire \current_shift_inst.z_5_5 ;
    wire \current_shift_inst.z_5_cry_4 ;
    wire \current_shift_inst.elapsed_time_ns_phase_6 ;
    wire \current_shift_inst.z_5_6 ;
    wire \current_shift_inst.z_5_cry_5 ;
    wire \current_shift_inst.elapsed_time_ns_phase_7 ;
    wire \current_shift_inst.z_5_7 ;
    wire \current_shift_inst.z_5_cry_6 ;
    wire \current_shift_inst.z_5_8 ;
    wire \current_shift_inst.z_5_cry_7 ;
    wire \current_shift_inst.z_5_cry_8 ;
    wire \current_shift_inst.z_5_9 ;
    wire bfn_10_19_0_;
    wire \current_shift_inst.elapsed_time_ns_phase_10 ;
    wire \current_shift_inst.z_5_10 ;
    wire \current_shift_inst.z_5_cry_9 ;
    wire \current_shift_inst.z_5_11 ;
    wire \current_shift_inst.z_5_cry_10 ;
    wire \current_shift_inst.z_5_12 ;
    wire \current_shift_inst.z_5_cry_11 ;
    wire \current_shift_inst.z_5_13 ;
    wire \current_shift_inst.z_5_cry_12 ;
    wire \current_shift_inst.z_5_14 ;
    wire \current_shift_inst.z_5_cry_13 ;
    wire \current_shift_inst.z_5_15 ;
    wire \current_shift_inst.z_5_cry_14 ;
    wire \current_shift_inst.z_5_16 ;
    wire \current_shift_inst.z_5_cry_15 ;
    wire \current_shift_inst.z_5_cry_16 ;
    wire \current_shift_inst.elapsed_time_ns_phase_17 ;
    wire \current_shift_inst.z_5_17 ;
    wire bfn_10_20_0_;
    wire \current_shift_inst.elapsed_time_ns_phase_18 ;
    wire \current_shift_inst.z_5_18 ;
    wire \current_shift_inst.z_5_cry_17 ;
    wire \current_shift_inst.z_5_19 ;
    wire \current_shift_inst.z_5_cry_18 ;
    wire \current_shift_inst.z_5_20 ;
    wire \current_shift_inst.z_5_cry_19 ;
    wire \current_shift_inst.z_5_21 ;
    wire \current_shift_inst.z_5_cry_20 ;
    wire \current_shift_inst.elapsed_time_ns_phase_22 ;
    wire \current_shift_inst.z_5_22 ;
    wire \current_shift_inst.z_5_cry_21 ;
    wire \current_shift_inst.z_5_23 ;
    wire \current_shift_inst.z_5_cry_22 ;
    wire \current_shift_inst.z_5_24 ;
    wire \current_shift_inst.z_5_cry_23 ;
    wire \current_shift_inst.z_5_cry_24 ;
    wire \current_shift_inst.z_5_25 ;
    wire bfn_10_21_0_;
    wire \current_shift_inst.z_5_26 ;
    wire \current_shift_inst.z_5_cry_25 ;
    wire \current_shift_inst.elapsed_time_ns_phase_27 ;
    wire \current_shift_inst.z_5_27 ;
    wire \current_shift_inst.z_5_cry_26 ;
    wire \current_shift_inst.z_5_28 ;
    wire \current_shift_inst.z_5_cry_27 ;
    wire \current_shift_inst.z_5_29 ;
    wire \current_shift_inst.z_5_cry_28 ;
    wire CONSTANT_ONE_NET;
    wire \current_shift_inst.z_5_30 ;
    wire \current_shift_inst.z_5_cry_29 ;
    wire \current_shift_inst.z_5_cry_30 ;
    wire \current_shift_inst.z_5_cry_30_THRU_CO ;
    wire s4_phy_c;
    wire il_min_comp1_c;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ;
    wire bfn_11_8_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7 ;
    wire bfn_11_9_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17 ;
    wire bfn_11_10_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19 ;
    wire il_min_comp1_D1;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ;
    wire \current_shift_inst.elapsed_time_ns_1_fast_31 ;
    wire \current_shift_inst.un38_control_input_0 ;
    wire bfn_11_14_0_;
    wire \current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0 ;
    wire \current_shift_inst.un4_control_input_cry_1 ;
    wire \current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0 ;
    wire \current_shift_inst.un4_control_input_cry_2 ;
    wire \current_shift_inst.un4_control_input_cry_3_c_RNINL4GZ0 ;
    wire \current_shift_inst.un4_control_input_cry_3 ;
    wire \current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0 ;
    wire \current_shift_inst.un4_control_input_cry_4 ;
    wire \current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0 ;
    wire \current_shift_inst.un4_control_input_cry_5 ;
    wire \current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0 ;
    wire \current_shift_inst.un4_control_input_cry_6 ;
    wire \current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0 ;
    wire \current_shift_inst.un4_control_input_cry_7 ;
    wire \current_shift_inst.un4_control_input_cry_8 ;
    wire bfn_11_15_0_;
    wire \current_shift_inst.un4_control_input_cry_9 ;
    wire \current_shift_inst.un4_control_input_cry_10_c_RNIJLTGZ0 ;
    wire \current_shift_inst.un4_control_input_cry_10 ;
    wire \current_shift_inst.un4_control_input_cry_11 ;
    wire \current_shift_inst.un4_control_input_cry_12 ;
    wire \current_shift_inst.un4_control_input_cry_13 ;
    wire \current_shift_inst.un4_control_input_cry_14 ;
    wire \current_shift_inst.un4_control_input_cry_15 ;
    wire \current_shift_inst.un4_control_input_cry_16 ;
    wire bfn_11_16_0_;
    wire \current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0 ;
    wire \current_shift_inst.un4_control_input_cry_17 ;
    wire \current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0 ;
    wire \current_shift_inst.un4_control_input_cry_18 ;
    wire \current_shift_inst.un4_control_input_cry_19 ;
    wire \current_shift_inst.un4_control_input_cry_20 ;
    wire \current_shift_inst.un4_control_input_cry_21 ;
    wire \current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0 ;
    wire \current_shift_inst.un4_control_input_cry_22 ;
    wire \current_shift_inst.un4_control_input_cry_23 ;
    wire \current_shift_inst.un4_control_input_cry_24 ;
    wire bfn_11_17_0_;
    wire \current_shift_inst.un4_control_input_cry_25 ;
    wire \current_shift_inst.un4_control_input_cry_26 ;
    wire \current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0 ;
    wire \current_shift_inst.un4_control_input_cry_27 ;
    wire \current_shift_inst.un4_control_input_cry_28 ;
    wire \current_shift_inst.un4_control_input_cry_29 ;
    wire \current_shift_inst.un4_control_input_cry_30 ;
    wire \current_shift_inst.elapsed_time_ns_phase_9 ;
    wire \current_shift_inst.un4_control_input_cry_9_c_RNIALDJZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIO0U12_8 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNILORI_11 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIOSSI_12 ;
    wire \current_shift_inst.elapsed_time_ns_phase_13 ;
    wire \current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJTQ51_12 ;
    wire \current_shift_inst.elapsed_time_ns_phase_8 ;
    wire \current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIN7DV_8 ;
    wire \current_shift_inst.elapsed_time_ns_phase_28 ;
    wire \current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIDS8K_28 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5S981_24 ;
    wire \current_shift_inst.elapsed_time_ns_phase_11 ;
    wire \current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0 ;
    wire \current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0 ;
    wire \current_shift_inst.elapsed_time_ns_phase_12 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIDLO51_11 ;
    wire \current_shift_inst.elapsed_time_ns_phase_30 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31 ;
    wire \current_shift_inst.elapsed_time_ns_phase_31 ;
    wire \current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0 ;
    wire \current_shift_inst.un38_control_input_0_axb_31 ;
    wire \current_shift_inst.elapsed_time_ns_phase_19 ;
    wire \current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPC571_19 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI190J_15 ;
    wire \current_shift_inst.elapsed_time_ns_phase_16 ;
    wire \current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5M161_15 ;
    wire \current_shift_inst.elapsed_time_ns_phase_14 ;
    wire \current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0 ;
    wire \current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0 ;
    wire \current_shift_inst.elapsed_time_ns_phase_15 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIVDV51_14 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIDR081_20 ;
    wire \current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0 ;
    wire \current_shift_inst.elapsed_time_ns_phase_20 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNILRVJ_20 ;
    wire \current_shift_inst.elapsed_time_ns_phase_21 ;
    wire \current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIOV0K_21 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIU73K_23 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI7K6K_26 ;
    wire il_max_comp2_D1;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst1.start_timer_hc_0_sqmuxa_cascade_ ;
    wire \phase_controller_inst1.N_88 ;
    wire \phase_controller_inst1.hc_time_passed ;
    wire \current_shift_inst.un4_control_input_axb_5 ;
    wire \current_shift_inst.un4_control_input_axb_6 ;
    wire \current_shift_inst.un4_control_input_axb_7 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ;
    wire \current_shift_inst.un4_control_input_axb_3 ;
    wire \current_shift_inst.un4_control_input_axb_4 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_1 ;
    wire \current_shift_inst.un4_control_input_axb_1 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_2 ;
    wire \current_shift_inst.un4_control_input_axb_2 ;
    wire \current_shift_inst.un4_control_input_axb_24 ;
    wire \current_shift_inst.un4_control_input_axb_15 ;
    wire \current_shift_inst.un4_control_input_axb_11 ;
    wire \current_shift_inst.un4_control_input_axb_19 ;
    wire \current_shift_inst.un4_control_input_axb_10 ;
    wire \current_shift_inst.un4_control_input_axb_12 ;
    wire \current_shift_inst.un4_control_input_axb_14 ;
    wire \current_shift_inst.un4_control_input_axb_18 ;
    wire \current_shift_inst.un4_control_input_axb_29 ;
    wire \current_shift_inst.un4_control_input_axb_22 ;
    wire \current_shift_inst.un4_control_input_axb_26 ;
    wire \current_shift_inst.un4_control_input_axb_27 ;
    wire \current_shift_inst.un4_control_input_axb_30 ;
    wire \current_shift_inst.un4_control_input_axb_21 ;
    wire \current_shift_inst.un4_control_input_axb_25 ;
    wire \current_shift_inst.un4_control_input_axb_20 ;
    wire \current_shift_inst.z_31 ;
    wire \current_shift_inst.z_i_31 ;
    wire \current_shift_inst.un4_control_input_axb_28 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI1C4K_24 ;
    wire \current_shift_inst.elapsed_time_ns_phase_26 ;
    wire \current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIB4C81_25 ;
    wire \current_shift_inst.elapsed_time_ns_phase_25 ;
    wire \current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI4G5K_25 ;
    wire \current_shift_inst.elapsed_time_ns_phase_29 ;
    wire \current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI7OAK_29 ;
    wire \current_shift_inst.elapsed_time_ns_phase_24 ;
    wire \current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0 ;
    wire \current_shift_inst.elapsed_time_ns_phase_23 ;
    wire \current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIVJ781_23 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1Z0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1Z0Z_6_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6_cascade_ ;
    wire \phase_controller_slave.start_timer_hc_0_sqmuxa_cascade_ ;
    wire s3_phy_c;
    wire \phase_controller_slave.stateZ0Z_1 ;
    wire il_min_comp2_D2;
    wire il_max_comp2_D2;
    wire \phase_controller_slave.stateZ0Z_3 ;
    wire \current_shift_inst.timer_phase.N_192_i ;
    wire \current_shift_inst.timer_phase.running_i ;
    wire clk_12mhz;
    wire GB_BUFFER_clk_12mhz_THRU_CO;
    wire \delay_measurement_inst.delay_hc_timer.N_321_i ;
    wire \current_shift_inst.N_199_cascade_ ;
    wire \current_shift_inst.timer_s1.N_187_i ;
    wire \current_shift_inst.phase_validZ0 ;
    wire \current_shift_inst.start_timer_sZ0Z1 ;
    wire \current_shift_inst.stop_timer_sZ0Z1 ;
    wire \current_shift_inst.meas_stateZ0Z_0 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto5Z0Z_3_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un1_startlt8 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_13 ;
    wire il_max_comp1_D2;
    wire \phase_controller_inst1.N_86_cascade_ ;
    wire \phase_controller_inst1.stateZ0Z_3 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_3 ;
    wire bfn_13_13_0_;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_4 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_5 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_6 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_7 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_10 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_11 ;
    wire bfn_13_14_0_;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_12 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_14 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_15 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_18 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_19 ;
    wire bfn_13_15_0_;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_20 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_21 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_22 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_24 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_25 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_26 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_27 ;
    wire bfn_13_16_0_;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_28 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_29 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_30 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ;
    wire \current_shift_inst.timer_s1.N_187_i_g ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ;
    wire \current_shift_inst.S1_riseZ0 ;
    wire s1_phy_c;
    wire \current_shift_inst.S1_syncZ0Z0 ;
    wire \current_shift_inst.S3_sync_prevZ0 ;
    wire \current_shift_inst.S3_riseZ0 ;
    wire \current_shift_inst.S1_syncZ0Z1 ;
    wire \current_shift_inst.S1_sync_prevZ0 ;
    wire \current_shift_inst.S3_syncZ0Z0 ;
    wire \current_shift_inst.S3_syncZ0Z1 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13_cascade_ ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_1 ;
    wire bfn_13_19_0_;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_9 ;
    wire bfn_13_20_0_;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_16 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_17 ;
    wire bfn_13_21_0_;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_18 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_i_19 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_19 ;
    wire \phase_controller_slave.stateZ0Z_0 ;
    wire \phase_controller_slave.stateZ0Z_4 ;
    wire \phase_controller_slave.start_timer_tr_0_sqmuxa ;
    wire \phase_controller_slave.N_210_cascade_ ;
    wire \phase_controller_slave.stoper_tr.time_passed11_cascade_ ;
    wire \phase_controller_slave.tr_time_passed ;
    wire \phase_controller_slave.stoper_tr.time_passed_1_sqmuxa ;
    wire bfn_13_23_0_;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7 ;
    wire bfn_13_24_0_;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15 ;
    wire bfn_13_25_0_;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19 ;
    wire \current_shift_inst.start_timer_phaseZ0 ;
    wire \current_shift_inst.timer_phase.runningZ0 ;
    wire \current_shift_inst.stop_timer_phaseZ0 ;
    wire \current_shift_inst.timer_phase.N_188_i ;
    wire s2_phy_c;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_3_cascade_ ;
    wire \delay_measurement_inst.stop_timer_hcZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt14_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt30_0 ;
    wire \delay_measurement_inst.delay_hc_timer.runningZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_2_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_11 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_1 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_2_tz ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a1_1_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_0 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_1_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_1 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt30 ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto13_3Z0Z_1_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto13 ;
    wire measured_delay_hc_20;
    wire \phase_controller_inst1.stoper_hc.un1_startlto30_2_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un1_startlt15 ;
    wire \delay_measurement_inst.tr_stateZ0Z_0 ;
    wire \delay_measurement_inst.prev_tr_sigZ0 ;
    wire \delay_measurement_inst.tr_state_RNIMR6LZ0Z_0_cascade_ ;
    wire \phase_controller_inst1.stateZ0Z_2 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_8 ;
    wire \current_shift_inst.un4_control_input_axb_8 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_23 ;
    wire \current_shift_inst.un4_control_input_axb_23 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_9 ;
    wire \current_shift_inst.un4_control_input_axb_9 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_16 ;
    wire \current_shift_inst.un4_control_input_axb_16 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_17 ;
    wire \current_shift_inst.un4_control_input_axb_17 ;
    wire \current_shift_inst.timer_s1.elapsed_time_ns_s1_13 ;
    wire \current_shift_inst.un4_control_input_axb_13 ;
    wire measured_delay_hc_15;
    wire measured_delay_hc_14;
    wire measured_delay_hc_6;
    wire measured_delay_hc_2;
    wire measured_delay_hc_9;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8 ;
    wire \phase_controller_slave.stoper_hc.time_passed_1_sqmuxa ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3Z0Z_3_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_5Z0Z_3 ;
    wire \phase_controller_slave.stoper_hc.time_passed11_cascade_ ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0 ;
    wire start_stop_c;
    wire shift_flag_start;
    wire \phase_controller_slave.un1_startZ0 ;
    wire \phase_controller_slave.stoper_tr.time_passed11 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ;
    wire bfn_14_22_0_;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7 ;
    wire bfn_14_23_0_;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15 ;
    wire bfn_14_24_0_;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18 ;
    wire delay_tr_input_c;
    wire delay_tr_d1;
    wire delay_tr_d2;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_4 ;
    wire \delay_measurement_inst.elapsed_time_hc_1 ;
    wire \delay_measurement_inst.elapsed_time_hc_2 ;
    wire \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6 ;
    wire bfn_15_7_0_;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.elapsed_time_hc_5 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_hc_reg3lto6 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_hc_reg3lto9 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.elapsed_time_hc_10 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.elapsed_time_hc_11 ;
    wire bfn_15_8_0_;
    wire \delay_measurement_inst.elapsed_time_hc_12 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.elapsed_time_hc_13 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_hc_reg3lto14 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_hc_reg3lto15 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.elapsed_time_hc_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ;
    wire bfn_15_9_0_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ;
    wire bfn_15_10_0_;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ;
    wire \delay_measurement_inst.delay_hc_timer.N_321_i_g ;
    wire measured_delay_hc_10;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2 ;
    wire \current_shift_inst.timer_s1.runningZ0 ;
    wire \delay_measurement_inst.elapsed_time_hc_3 ;
    wire measured_delay_hc_3;
    wire \delay_measurement_inst.elapsed_time_hc_4 ;
    wire measured_delay_hc_4;
    wire \delay_measurement_inst.hc_stateZ0Z_0 ;
    wire \delay_measurement_inst.start_timer_hcZ0 ;
    wire \delay_measurement_inst.prev_hc_sigZ0 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_0 ;
    wire bfn_15_13_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_1 ;
    wire \current_shift_inst.timer_s1.counter_cry_0 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_2 ;
    wire \current_shift_inst.timer_s1.counter_cry_1 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_3 ;
    wire \current_shift_inst.timer_s1.counter_cry_2 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_4 ;
    wire \current_shift_inst.timer_s1.counter_cry_3 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_5 ;
    wire \current_shift_inst.timer_s1.counter_cry_4 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_5 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_7 ;
    wire \current_shift_inst.timer_s1.counter_cry_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_7 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_8 ;
    wire bfn_15_14_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_9 ;
    wire \current_shift_inst.timer_s1.counter_cry_8 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_10 ;
    wire \current_shift_inst.timer_s1.counter_cry_9 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_11 ;
    wire \current_shift_inst.timer_s1.counter_cry_10 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_12 ;
    wire \current_shift_inst.timer_s1.counter_cry_11 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_13 ;
    wire \current_shift_inst.timer_s1.counter_cry_12 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_13 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_15 ;
    wire \current_shift_inst.timer_s1.counter_cry_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_15 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_16 ;
    wire bfn_15_15_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_17 ;
    wire \current_shift_inst.timer_s1.counter_cry_16 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_18 ;
    wire \current_shift_inst.timer_s1.counter_cry_17 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_19 ;
    wire \current_shift_inst.timer_s1.counter_cry_18 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_20 ;
    wire \current_shift_inst.timer_s1.counter_cry_19 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_21 ;
    wire \current_shift_inst.timer_s1.counter_cry_20 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_21 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_23 ;
    wire \current_shift_inst.timer_s1.counter_cry_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_23 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_24 ;
    wire bfn_15_16_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_25 ;
    wire \current_shift_inst.timer_s1.counter_cry_24 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_26 ;
    wire \current_shift_inst.timer_s1.counter_cry_25 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_27 ;
    wire \current_shift_inst.timer_s1.counter_cry_26 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_28 ;
    wire \current_shift_inst.timer_s1.counter_cry_27 ;
    wire \current_shift_inst.timer_s1.running_i ;
    wire \current_shift_inst.timer_s1.counter_cry_28 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_29 ;
    wire \current_shift_inst.timer_s1.N_191_i ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_0 ;
    wire bfn_15_17_0_;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_1 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ1Z_6 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_8 ;
    wire bfn_15_18_0_;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_9 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_16 ;
    wire bfn_15_19_0_;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_17 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_18 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_i_19 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_slave.stoper_hc.time_passed11 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.N_20_li ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3 ;
    wire \delay_measurement_inst.stop_timer_trZ0 ;
    wire \delay_measurement_inst.start_timer_trZ0 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6 ;
    wire measured_delay_tr_7;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6 ;
    wire measured_delay_tr_8;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ;
    wire \phase_controller_slave.start_timer_trZ0 ;
    wire \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19 ;
    wire \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ;
    wire \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15 ;
    wire \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ;
    wire bfn_16_7_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ;
    wire bfn_16_8_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ;
    wire bfn_16_9_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ;
    wire bfn_16_10_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.running_i ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_hc_timer.N_322_i ;
    wire measured_delay_hc_12;
    wire measured_delay_hc_11;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9 ;
    wire \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_5 ;
    wire \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_6_cascade_ ;
    wire \delay_measurement_inst.tr_state_RNIMR6LZ0Z_0 ;
    wire \delay_measurement_inst.delay_tr_timer.N_375_cascade_ ;
    wire \delay_measurement_inst.N_265_i_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.runningZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_4 ;
    wire \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_6_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_364 ;
    wire \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_5 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_6_19_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_0_19 ;
    wire \delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_409 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_400_cascade_ ;
    wire \delay_measurement_inst.N_394_1_cascade_ ;
    wire \delay_measurement_inst.N_394_1 ;
    wire measured_delay_tr_12;
    wire measured_delay_tr_10;
    wire measured_delay_tr_6;
    wire measured_delay_tr_3;
    wire measured_delay_tr_5;
    wire \delay_measurement_inst.elapsed_time_tr_1 ;
    wire measured_delay_tr_1;
    wire measured_delay_tr_2;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_inst1.start_timer_hcZ0 ;
    wire \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ;
    wire \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ;
    wire \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ;
    wire \phase_controller_slave.start_timer_hcZ0 ;
    wire \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ;
    wire red_c_i;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_8 ;
    wire measured_delay_hc_16;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlt31 ;
    wire measured_delay_hc_1;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_1 ;
    wire bfn_16_19_0_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_9 ;
    wire bfn_16_20_0_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_17 ;
    wire bfn_16_21_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_19 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ;
    wire measured_delay_tr_19;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ;
    wire measured_delay_tr_11;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ;
    wire measured_delay_tr_13;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ;
    wire delay_hc_input_c;
    wire delay_hc_d1;
    wire delay_hc_d2;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_2 ;
    wire measured_delay_hc_25;
    wire measured_delay_hc_26;
    wire measured_delay_hc_23;
    wire \delay_measurement_inst.elapsed_time_hc_8 ;
    wire measured_delay_hc_8;
    wire \delay_measurement_inst.elapsed_time_hc_7 ;
    wire measured_delay_hc_7;
    wire measured_delay_hc_24;
    wire measured_delay_hc_0;
    wire \delay_measurement_inst.elapsed_time_hc_18 ;
    wire measured_delay_hc_18;
    wire \delay_measurement_inst.elapsed_time_hc_19 ;
    wire \delay_measurement_inst.delay_hc_reg3lto31_0_0 ;
    wire measured_delay_hc_19;
    wire measured_delay_hc_21;
    wire measured_delay_hc_22;
    wire \delay_measurement_inst.un1_elapsed_time_hc ;
    wire \delay_measurement_inst.elapsed_time_hc_17 ;
    wire \delay_measurement_inst.delay_hc_reg3 ;
    wire measured_delay_hc_17;
    wire bfn_17_11_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_7 ;
    wire bfn_17_12_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_15 ;
    wire bfn_17_13_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_23 ;
    wire bfn_17_14_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.running_i ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.N_324_i ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_7_19 ;
    wire \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_4 ;
    wire \delay_measurement_inst.elapsed_time_tr_2 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16 ;
    wire measured_delay_tr_17;
    wire \delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20 ;
    wire measured_delay_tr_18;
    wire \phase_controller_inst1.N_83 ;
    wire \phase_controller_inst1.stateZ0Z_4 ;
    wire \phase_controller_inst1.N_83_cascade_ ;
    wire \phase_controller_inst1.T01_0_sqmuxa ;
    wire \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa_cascade_ ;
    wire \phase_controller_inst1.stateZ0Z_1 ;
    wire \phase_controller_inst1.tr_time_passed ;
    wire il_min_comp1_D2;
    wire \phase_controller_inst1.stateZ0Z_0 ;
    wire \phase_controller_inst1.stoper_tr.time_passed11_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.time_passed11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ;
    wire \phase_controller_slave.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa ;
    wire measured_delay_tr_16;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ;
    wire measured_delay_hc_29;
    wire measured_delay_hc_28;
    wire measured_delay_hc_30;
    wire measured_delay_hc_27;
    wire \phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_4 ;
    wire measured_delay_hc_13;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_13 ;
    wire measured_delay_hc_31;
    wire measured_delay_hc_5;
    wire \phase_controller_inst1.stoper_hc.un1_startlt31_0 ;
    wire \phase_controller_slave.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa ;
    wire \delay_measurement_inst.N_410 ;
    wire \delay_measurement_inst.N_358 ;
    wire \delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15 ;
    wire measured_delay_tr_4;
    wire \delay_measurement_inst.N_265_i_0 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ;
    wire \delay_measurement_inst.elapsed_time_tr_3 ;
    wire bfn_18_13_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.elapsed_time_tr_4 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.elapsed_time_tr_5 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.elapsed_time_tr_6 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.elapsed_time_tr_7 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.elapsed_time_tr_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.elapsed_time_tr_9 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.elapsed_time_tr_10 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ;
    wire \delay_measurement_inst.elapsed_time_tr_11 ;
    wire bfn_18_14_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.elapsed_time_tr_12 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.elapsed_time_tr_13 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.elapsed_time_tr_15 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.elapsed_time_tr_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.elapsed_time_tr_17 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.elapsed_time_tr_18 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ;
    wire \delay_measurement_inst.elapsed_time_tr_19 ;
    wire bfn_18_15_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ;
    wire bfn_18_16_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.elapsed_time_tr_31 ;
    wire \delay_measurement_inst.delay_tr_timer.N_323_i ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ;
    wire bfn_18_17_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7 ;
    wire bfn_18_18_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17 ;
    wire bfn_18_19_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst1.start_timer_trZ0 ;
    wire \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ;
    wire \phase_controller_inst1.stoper_tr.N_21 ;
    wire \delay_measurement_inst.N_271_1 ;
    wire \delay_measurement_inst.elapsed_time_tr_14 ;
    wire \delay_measurement_inst.N_265_i ;
    wire measured_delay_tr_14;
    wire \phase_controller_slave.hc_time_passed ;
    wire \phase_controller_slave.stateZ0Z_2 ;
    wire \phase_controller_slave.N_211 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13 ;
    wire measured_delay_tr_15;
    wire measured_delay_tr_9;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0Z0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ;
    wire _gnd_net_;
    wire clk_100mhz_0;
    wire \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ;
    wire red_c_g;

    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .TEST_MODE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FILTER_RANGE=3'b001;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVR=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVQ=3'b011;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVF=7'b1000010;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__31943),
            .RESETB(N__40529),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(clk_100mhz_0));
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__28856),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__28849),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15}),
            .ADDSUBBOT(),
            .A({dangling_wire_16,N__18887,N__18890,N__18888,N__18891,N__18889,N__19120,N__19100,N__19064,N__20811,N__19139,N__18846,N__19002,N__18970,N__19015,N__18982}),
            .C({dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31,dangling_wire_32}),
            .B({dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,N__28855,N__28852,dangling_wire_40,dangling_wire_41,dangling_wire_42,N__28850,N__28854,N__28851,N__28853}),
            .OHOLDTOP(),
            .O({dangling_wire_43,dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,dangling_wire_48,\pwm_generator_inst.un2_threshold_acc_1_25 ,\pwm_generator_inst.un2_threshold_acc_1_24 ,\pwm_generator_inst.un2_threshold_acc_1_23 ,\pwm_generator_inst.un2_threshold_acc_1_22 ,\pwm_generator_inst.un2_threshold_acc_1_21 ,\pwm_generator_inst.un2_threshold_acc_1_20 ,\pwm_generator_inst.un2_threshold_acc_1_19 ,\pwm_generator_inst.un2_threshold_acc_1_18 ,\pwm_generator_inst.un2_threshold_acc_1_17 ,\pwm_generator_inst.un2_threshold_acc_1_16 ,\pwm_generator_inst.un2_threshold_acc_1_15 ,\pwm_generator_inst.O_14 ,\pwm_generator_inst.O_13 ,\pwm_generator_inst.O_12 ,\pwm_generator_inst.un3_threshold_acc ,\pwm_generator_inst.O_10 ,\pwm_generator_inst.O_9 ,\pwm_generator_inst.O_8 ,\pwm_generator_inst.O_7 ,\pwm_generator_inst.O_6 ,\pwm_generator_inst.O_5 ,\pwm_generator_inst.O_4 ,\pwm_generator_inst.O_3 ,\pwm_generator_inst.O_2 ,\pwm_generator_inst.O_1 ,\pwm_generator_inst.O_0 }));
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__28731),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__28817),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64}),
            .ADDSUBBOT(),
            .A({dangling_wire_65,N__18950,N__18943,N__18948,N__18942,N__18949,N__18941,N__18951,N__18938,N__18944,N__18937,N__18945,N__18939,N__18946,N__18940,N__18947}),
            .C({dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73,dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81}),
            .B({dangling_wire_82,dangling_wire_83,dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,N__28823,N__28820,dangling_wire_89,dangling_wire_90,dangling_wire_91,N__28818,N__28822,N__28819,N__28821}),
            .OHOLDTOP(),
            .O({dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,\pwm_generator_inst.un2_threshold_acc_2_1_16 ,\pwm_generator_inst.un2_threshold_acc_2_1_15 ,\pwm_generator_inst.un2_threshold_acc_2_14 ,\pwm_generator_inst.un2_threshold_acc_2_13 ,\pwm_generator_inst.un2_threshold_acc_2_12 ,\pwm_generator_inst.un2_threshold_acc_2_11 ,\pwm_generator_inst.un2_threshold_acc_2_10 ,\pwm_generator_inst.un2_threshold_acc_2_9 ,\pwm_generator_inst.un2_threshold_acc_2_8 ,\pwm_generator_inst.un2_threshold_acc_2_7 ,\pwm_generator_inst.un2_threshold_acc_2_6 ,\pwm_generator_inst.un2_threshold_acc_2_5 ,\pwm_generator_inst.un2_threshold_acc_2_4 ,\pwm_generator_inst.un2_threshold_acc_2_3 ,\pwm_generator_inst.un2_threshold_acc_2_2 ,\pwm_generator_inst.un2_threshold_acc_2_1 ,\pwm_generator_inst.un2_threshold_acc_2_0 }));
    PRE_IO_GBUF reset_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__48351),
            .GLOBALBUFFEROUTPUT(red_c_g));
    IO_PAD reset_ibuf_gb_io_iopad (
            .OE(N__48353),
            .DIN(N__48352),
            .DOUT(N__48351),
            .PACKAGEPIN(reset));
    defparam reset_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam reset_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO reset_ibuf_gb_io_preio (
            .PADOEN(N__48353),
            .PADOUT(N__48352),
            .PADIN(N__48351),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD start_stop_ibuf_iopad (
            .OE(N__48342),
            .DIN(N__48341),
            .DOUT(N__48340),
            .PACKAGEPIN(start_stop));
    defparam start_stop_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam start_stop_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO start_stop_ibuf_preio (
            .PADOEN(N__48342),
            .PADOUT(N__48341),
            .PADIN(N__48340),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(start_stop_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp2_ibuf_iopad (
            .OE(N__48333),
            .DIN(N__48332),
            .DOUT(N__48331),
            .PACKAGEPIN(il_max_comp2));
    defparam il_max_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp2_ibuf_preio (
            .PADOEN(N__48333),
            .PADOUT(N__48332),
            .PADIN(N__48331),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_output_obuf_iopad (
            .OE(N__48324),
            .DIN(N__48323),
            .DOUT(N__48322),
            .PACKAGEPIN(pwm_output));
    defparam pwm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam pwm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO pwm_output_obuf_preio (
            .PADOEN(N__48324),
            .PADOUT(N__48323),
            .PADIN(N__48322),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23270),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp1_ibuf_iopad (
            .OE(N__48315),
            .DIN(N__48314),
            .DOUT(N__48313),
            .PACKAGEPIN(il_max_comp1));
    defparam il_max_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp1_ibuf_preio (
            .PADOEN(N__48315),
            .PADOUT(N__48314),
            .PADIN(N__48313),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s2_phy_obuf_iopad (
            .OE(N__48306),
            .DIN(N__48305),
            .DOUT(N__48304),
            .PACKAGEPIN(s2_phy));
    defparam s2_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s2_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s2_phy_obuf_preio (
            .PADOEN(N__48306),
            .PADOUT(N__48305),
            .PADIN(N__48304),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__33443),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_hc_input_ibuf_iopad (
            .OE(N__48297),
            .DIN(N__48296),
            .DOUT(N__48295),
            .PACKAGEPIN(delay_hc_input));
    defparam delay_hc_input_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam delay_hc_input_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_hc_input_ibuf_preio (
            .PADOEN(N__48297),
            .PADOUT(N__48296),
            .PADIN(N__48295),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_hc_input_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_tr_input_ibuf_iopad (
            .OE(N__48288),
            .DIN(N__48287),
            .DOUT(N__48286),
            .PACKAGEPIN(delay_tr_input));
    defparam delay_tr_input_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam delay_tr_input_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_tr_input_ibuf_preio (
            .PADOEN(N__48288),
            .PADOUT(N__48287),
            .PADIN(N__48286),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_tr_input_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp2_ibuf_iopad (
            .OE(N__48279),
            .DIN(N__48278),
            .DOUT(N__48277),
            .PACKAGEPIN(il_min_comp2));
    defparam il_min_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp2_ibuf_preio (
            .PADOEN(N__48279),
            .PADOUT(N__48278),
            .PADIN(N__48277),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s1_phy_obuf_iopad (
            .OE(N__48270),
            .DIN(N__48269),
            .DOUT(N__48268),
            .PACKAGEPIN(s1_phy));
    defparam s1_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s1_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s1_phy_obuf_preio (
            .PADOEN(N__48270),
            .PADOUT(N__48269),
            .PADIN(N__48268),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__32888),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s4_phy_obuf_iopad (
            .OE(N__48261),
            .DIN(N__48260),
            .DOUT(N__48259),
            .PACKAGEPIN(s4_phy));
    defparam s4_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s4_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s4_phy_obuf_preio (
            .PADOEN(N__48261),
            .PADOUT(N__48260),
            .PADIN(N__48259),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__28436),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp1_ibuf_iopad (
            .OE(N__48252),
            .DIN(N__48251),
            .DOUT(N__48250),
            .PACKAGEPIN(il_min_comp1));
    defparam il_min_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp1_ibuf_preio (
            .PADOEN(N__48252),
            .PADOUT(N__48251),
            .PADIN(N__48250),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s3_phy_obuf_iopad (
            .OE(N__48243),
            .DIN(N__48242),
            .DOUT(N__48241),
            .PACKAGEPIN(s3_phy));
    defparam s3_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s3_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s3_phy_obuf_preio (
            .PADOEN(N__48243),
            .PADOUT(N__48242),
            .PADIN(N__48241),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__31913),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__11547 (
            .O(N__48224),
            .I(N__48221));
    LocalMux I__11546 (
            .O(N__48221),
            .I(N__48218));
    Odrv4 I__11545 (
            .O(N__48218),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9 ));
    InMux I__11544 (
            .O(N__48215),
            .I(N__48211));
    InMux I__11543 (
            .O(N__48214),
            .I(N__48208));
    LocalMux I__11542 (
            .O(N__48211),
            .I(N__48205));
    LocalMux I__11541 (
            .O(N__48208),
            .I(N__48202));
    Odrv4 I__11540 (
            .O(N__48205),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    Odrv4 I__11539 (
            .O(N__48202),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    CascadeMux I__11538 (
            .O(N__48197),
            .I(N__48192));
    CascadeMux I__11537 (
            .O(N__48196),
            .I(N__48189));
    CascadeMux I__11536 (
            .O(N__48195),
            .I(N__48186));
    InMux I__11535 (
            .O(N__48192),
            .I(N__48164));
    InMux I__11534 (
            .O(N__48189),
            .I(N__48164));
    InMux I__11533 (
            .O(N__48186),
            .I(N__48164));
    InMux I__11532 (
            .O(N__48185),
            .I(N__48164));
    InMux I__11531 (
            .O(N__48184),
            .I(N__48159));
    InMux I__11530 (
            .O(N__48183),
            .I(N__48159));
    CascadeMux I__11529 (
            .O(N__48182),
            .I(N__48150));
    CascadeMux I__11528 (
            .O(N__48181),
            .I(N__48146));
    CascadeMux I__11527 (
            .O(N__48180),
            .I(N__48142));
    CascadeMux I__11526 (
            .O(N__48179),
            .I(N__48139));
    InMux I__11525 (
            .O(N__48178),
            .I(N__48126));
    InMux I__11524 (
            .O(N__48177),
            .I(N__48126));
    InMux I__11523 (
            .O(N__48176),
            .I(N__48126));
    InMux I__11522 (
            .O(N__48175),
            .I(N__48126));
    InMux I__11521 (
            .O(N__48174),
            .I(N__48126));
    InMux I__11520 (
            .O(N__48173),
            .I(N__48126));
    LocalMux I__11519 (
            .O(N__48164),
            .I(N__48121));
    LocalMux I__11518 (
            .O(N__48159),
            .I(N__48121));
    InMux I__11517 (
            .O(N__48158),
            .I(N__48118));
    InMux I__11516 (
            .O(N__48157),
            .I(N__48115));
    InMux I__11515 (
            .O(N__48156),
            .I(N__48110));
    InMux I__11514 (
            .O(N__48155),
            .I(N__48110));
    InMux I__11513 (
            .O(N__48154),
            .I(N__48093));
    InMux I__11512 (
            .O(N__48153),
            .I(N__48093));
    InMux I__11511 (
            .O(N__48150),
            .I(N__48093));
    InMux I__11510 (
            .O(N__48149),
            .I(N__48093));
    InMux I__11509 (
            .O(N__48146),
            .I(N__48093));
    InMux I__11508 (
            .O(N__48145),
            .I(N__48093));
    InMux I__11507 (
            .O(N__48142),
            .I(N__48093));
    InMux I__11506 (
            .O(N__48139),
            .I(N__48093));
    LocalMux I__11505 (
            .O(N__48126),
            .I(N__48088));
    Span4Mux_v I__11504 (
            .O(N__48121),
            .I(N__48088));
    LocalMux I__11503 (
            .O(N__48118),
            .I(N__48085));
    LocalMux I__11502 (
            .O(N__48115),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    LocalMux I__11501 (
            .O(N__48110),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    LocalMux I__11500 (
            .O(N__48093),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv4 I__11499 (
            .O(N__48088),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv4 I__11498 (
            .O(N__48085),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    CascadeMux I__11497 (
            .O(N__48074),
            .I(N__48068));
    CascadeMux I__11496 (
            .O(N__48073),
            .I(N__48056));
    CascadeMux I__11495 (
            .O(N__48072),
            .I(N__48053));
    CascadeMux I__11494 (
            .O(N__48071),
            .I(N__48050));
    InMux I__11493 (
            .O(N__48068),
            .I(N__48042));
    InMux I__11492 (
            .O(N__48067),
            .I(N__48042));
    CascadeMux I__11491 (
            .O(N__48066),
            .I(N__48039));
    CascadeMux I__11490 (
            .O(N__48065),
            .I(N__48036));
    CascadeMux I__11489 (
            .O(N__48064),
            .I(N__48033));
    CascadeMux I__11488 (
            .O(N__48063),
            .I(N__48030));
    InMux I__11487 (
            .O(N__48062),
            .I(N__48015));
    InMux I__11486 (
            .O(N__48061),
            .I(N__48015));
    InMux I__11485 (
            .O(N__48060),
            .I(N__48015));
    InMux I__11484 (
            .O(N__48059),
            .I(N__48015));
    InMux I__11483 (
            .O(N__48056),
            .I(N__48002));
    InMux I__11482 (
            .O(N__48053),
            .I(N__48002));
    InMux I__11481 (
            .O(N__48050),
            .I(N__48002));
    InMux I__11480 (
            .O(N__48049),
            .I(N__48002));
    InMux I__11479 (
            .O(N__48048),
            .I(N__48002));
    InMux I__11478 (
            .O(N__48047),
            .I(N__48002));
    LocalMux I__11477 (
            .O(N__48042),
            .I(N__47999));
    InMux I__11476 (
            .O(N__48039),
            .I(N__47988));
    InMux I__11475 (
            .O(N__48036),
            .I(N__47988));
    InMux I__11474 (
            .O(N__48033),
            .I(N__47988));
    InMux I__11473 (
            .O(N__48030),
            .I(N__47988));
    InMux I__11472 (
            .O(N__48029),
            .I(N__47983));
    InMux I__11471 (
            .O(N__48028),
            .I(N__47983));
    InMux I__11470 (
            .O(N__48027),
            .I(N__47974));
    InMux I__11469 (
            .O(N__48026),
            .I(N__47974));
    InMux I__11468 (
            .O(N__48025),
            .I(N__47974));
    InMux I__11467 (
            .O(N__48024),
            .I(N__47974));
    LocalMux I__11466 (
            .O(N__48015),
            .I(N__47969));
    LocalMux I__11465 (
            .O(N__48002),
            .I(N__47969));
    Span4Mux_h I__11464 (
            .O(N__47999),
            .I(N__47966));
    InMux I__11463 (
            .O(N__47998),
            .I(N__47961));
    InMux I__11462 (
            .O(N__47997),
            .I(N__47961));
    LocalMux I__11461 (
            .O(N__47988),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    LocalMux I__11460 (
            .O(N__47983),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    LocalMux I__11459 (
            .O(N__47974),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__11458 (
            .O(N__47969),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__11457 (
            .O(N__47966),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    LocalMux I__11456 (
            .O(N__47961),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    CascadeMux I__11455 (
            .O(N__47948),
            .I(N__47943));
    CascadeMux I__11454 (
            .O(N__47947),
            .I(N__47937));
    CascadeMux I__11453 (
            .O(N__47946),
            .I(N__47934));
    InMux I__11452 (
            .O(N__47943),
            .I(N__47930));
    InMux I__11451 (
            .O(N__47942),
            .I(N__47923));
    InMux I__11450 (
            .O(N__47941),
            .I(N__47923));
    InMux I__11449 (
            .O(N__47940),
            .I(N__47923));
    InMux I__11448 (
            .O(N__47937),
            .I(N__47916));
    InMux I__11447 (
            .O(N__47934),
            .I(N__47916));
    InMux I__11446 (
            .O(N__47933),
            .I(N__47916));
    LocalMux I__11445 (
            .O(N__47930),
            .I(N__47903));
    LocalMux I__11444 (
            .O(N__47923),
            .I(N__47903));
    LocalMux I__11443 (
            .O(N__47916),
            .I(N__47903));
    InMux I__11442 (
            .O(N__47915),
            .I(N__47898));
    InMux I__11441 (
            .O(N__47914),
            .I(N__47898));
    CascadeMux I__11440 (
            .O(N__47913),
            .I(N__47895));
    InMux I__11439 (
            .O(N__47912),
            .I(N__47879));
    InMux I__11438 (
            .O(N__47911),
            .I(N__47879));
    InMux I__11437 (
            .O(N__47910),
            .I(N__47879));
    Span4Mux_v I__11436 (
            .O(N__47903),
            .I(N__47874));
    LocalMux I__11435 (
            .O(N__47898),
            .I(N__47874));
    InMux I__11434 (
            .O(N__47895),
            .I(N__47867));
    InMux I__11433 (
            .O(N__47894),
            .I(N__47867));
    InMux I__11432 (
            .O(N__47893),
            .I(N__47850));
    InMux I__11431 (
            .O(N__47892),
            .I(N__47850));
    InMux I__11430 (
            .O(N__47891),
            .I(N__47850));
    InMux I__11429 (
            .O(N__47890),
            .I(N__47850));
    InMux I__11428 (
            .O(N__47889),
            .I(N__47850));
    InMux I__11427 (
            .O(N__47888),
            .I(N__47850));
    InMux I__11426 (
            .O(N__47887),
            .I(N__47850));
    InMux I__11425 (
            .O(N__47886),
            .I(N__47850));
    LocalMux I__11424 (
            .O(N__47879),
            .I(N__47845));
    Span4Mux_h I__11423 (
            .O(N__47874),
            .I(N__47845));
    InMux I__11422 (
            .O(N__47873),
            .I(N__47840));
    InMux I__11421 (
            .O(N__47872),
            .I(N__47840));
    LocalMux I__11420 (
            .O(N__47867),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    LocalMux I__11419 (
            .O(N__47850),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__11418 (
            .O(N__47845),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    LocalMux I__11417 (
            .O(N__47840),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    InMux I__11416 (
            .O(N__47831),
            .I(N__47828));
    LocalMux I__11415 (
            .O(N__47828),
            .I(N__47825));
    Span4Mux_v I__11414 (
            .O(N__47825),
            .I(N__47821));
    InMux I__11413 (
            .O(N__47824),
            .I(N__47818));
    Sp12to4 I__11412 (
            .O(N__47821),
            .I(N__47813));
    LocalMux I__11411 (
            .O(N__47818),
            .I(N__47813));
    Odrv12 I__11410 (
            .O(N__47813),
            .I(\phase_controller_inst1.stoper_tr.N_21 ));
    InMux I__11409 (
            .O(N__47810),
            .I(N__47807));
    LocalMux I__11408 (
            .O(N__47807),
            .I(N__47803));
    CascadeMux I__11407 (
            .O(N__47806),
            .I(N__47800));
    Span4Mux_h I__11406 (
            .O(N__47803),
            .I(N__47797));
    InMux I__11405 (
            .O(N__47800),
            .I(N__47794));
    Span4Mux_v I__11404 (
            .O(N__47797),
            .I(N__47791));
    LocalMux I__11403 (
            .O(N__47794),
            .I(N__47788));
    Odrv4 I__11402 (
            .O(N__47791),
            .I(\delay_measurement_inst.N_271_1 ));
    Odrv4 I__11401 (
            .O(N__47788),
            .I(\delay_measurement_inst.N_271_1 ));
    InMux I__11400 (
            .O(N__47783),
            .I(N__47776));
    InMux I__11399 (
            .O(N__47782),
            .I(N__47773));
    InMux I__11398 (
            .O(N__47781),
            .I(N__47770));
    InMux I__11397 (
            .O(N__47780),
            .I(N__47767));
    InMux I__11396 (
            .O(N__47779),
            .I(N__47764));
    LocalMux I__11395 (
            .O(N__47776),
            .I(N__47761));
    LocalMux I__11394 (
            .O(N__47773),
            .I(N__47756));
    LocalMux I__11393 (
            .O(N__47770),
            .I(N__47756));
    LocalMux I__11392 (
            .O(N__47767),
            .I(N__47753));
    LocalMux I__11391 (
            .O(N__47764),
            .I(N__47750));
    Span4Mux_v I__11390 (
            .O(N__47761),
            .I(N__47745));
    Span4Mux_v I__11389 (
            .O(N__47756),
            .I(N__47745));
    Span4Mux_h I__11388 (
            .O(N__47753),
            .I(N__47742));
    Odrv12 I__11387 (
            .O(N__47750),
            .I(\delay_measurement_inst.elapsed_time_tr_14 ));
    Odrv4 I__11386 (
            .O(N__47745),
            .I(\delay_measurement_inst.elapsed_time_tr_14 ));
    Odrv4 I__11385 (
            .O(N__47742),
            .I(\delay_measurement_inst.elapsed_time_tr_14 ));
    InMux I__11384 (
            .O(N__47735),
            .I(N__47732));
    LocalMux I__11383 (
            .O(N__47732),
            .I(N__47729));
    Span4Mux_v I__11382 (
            .O(N__47729),
            .I(N__47726));
    Span4Mux_v I__11381 (
            .O(N__47726),
            .I(N__47720));
    InMux I__11380 (
            .O(N__47725),
            .I(N__47713));
    InMux I__11379 (
            .O(N__47724),
            .I(N__47713));
    InMux I__11378 (
            .O(N__47723),
            .I(N__47713));
    Odrv4 I__11377 (
            .O(N__47720),
            .I(\delay_measurement_inst.N_265_i ));
    LocalMux I__11376 (
            .O(N__47713),
            .I(\delay_measurement_inst.N_265_i ));
    InMux I__11375 (
            .O(N__47708),
            .I(N__47701));
    InMux I__11374 (
            .O(N__47707),
            .I(N__47701));
    InMux I__11373 (
            .O(N__47706),
            .I(N__47698));
    LocalMux I__11372 (
            .O(N__47701),
            .I(N__47695));
    LocalMux I__11371 (
            .O(N__47698),
            .I(N__47691));
    Span4Mux_h I__11370 (
            .O(N__47695),
            .I(N__47688));
    CascadeMux I__11369 (
            .O(N__47694),
            .I(N__47685));
    Span4Mux_h I__11368 (
            .O(N__47691),
            .I(N__47681));
    Span4Mux_h I__11367 (
            .O(N__47688),
            .I(N__47678));
    InMux I__11366 (
            .O(N__47685),
            .I(N__47673));
    InMux I__11365 (
            .O(N__47684),
            .I(N__47673));
    Odrv4 I__11364 (
            .O(N__47681),
            .I(measured_delay_tr_14));
    Odrv4 I__11363 (
            .O(N__47678),
            .I(measured_delay_tr_14));
    LocalMux I__11362 (
            .O(N__47673),
            .I(measured_delay_tr_14));
    InMux I__11361 (
            .O(N__47666),
            .I(N__47660));
    InMux I__11360 (
            .O(N__47665),
            .I(N__47657));
    InMux I__11359 (
            .O(N__47664),
            .I(N__47652));
    InMux I__11358 (
            .O(N__47663),
            .I(N__47652));
    LocalMux I__11357 (
            .O(N__47660),
            .I(N__47649));
    LocalMux I__11356 (
            .O(N__47657),
            .I(\phase_controller_slave.hc_time_passed ));
    LocalMux I__11355 (
            .O(N__47652),
            .I(\phase_controller_slave.hc_time_passed ));
    Odrv12 I__11354 (
            .O(N__47649),
            .I(\phase_controller_slave.hc_time_passed ));
    InMux I__11353 (
            .O(N__47642),
            .I(N__47638));
    CascadeMux I__11352 (
            .O(N__47641),
            .I(N__47634));
    LocalMux I__11351 (
            .O(N__47638),
            .I(N__47631));
    InMux I__11350 (
            .O(N__47637),
            .I(N__47628));
    InMux I__11349 (
            .O(N__47634),
            .I(N__47625));
    Span4Mux_h I__11348 (
            .O(N__47631),
            .I(N__47622));
    LocalMux I__11347 (
            .O(N__47628),
            .I(\phase_controller_slave.stateZ0Z_2 ));
    LocalMux I__11346 (
            .O(N__47625),
            .I(\phase_controller_slave.stateZ0Z_2 ));
    Odrv4 I__11345 (
            .O(N__47622),
            .I(\phase_controller_slave.stateZ0Z_2 ));
    InMux I__11344 (
            .O(N__47615),
            .I(N__47612));
    LocalMux I__11343 (
            .O(N__47612),
            .I(N__47609));
    Odrv12 I__11342 (
            .O(N__47609),
            .I(\phase_controller_slave.N_211 ));
    InMux I__11341 (
            .O(N__47606),
            .I(N__47599));
    InMux I__11340 (
            .O(N__47605),
            .I(N__47599));
    InMux I__11339 (
            .O(N__47604),
            .I(N__47590));
    LocalMux I__11338 (
            .O(N__47599),
            .I(N__47587));
    InMux I__11337 (
            .O(N__47598),
            .I(N__47578));
    InMux I__11336 (
            .O(N__47597),
            .I(N__47578));
    InMux I__11335 (
            .O(N__47596),
            .I(N__47578));
    InMux I__11334 (
            .O(N__47595),
            .I(N__47578));
    InMux I__11333 (
            .O(N__47594),
            .I(N__47573));
    InMux I__11332 (
            .O(N__47593),
            .I(N__47573));
    LocalMux I__11331 (
            .O(N__47590),
            .I(N__47570));
    Span4Mux_v I__11330 (
            .O(N__47587),
            .I(N__47567));
    LocalMux I__11329 (
            .O(N__47578),
            .I(N__47564));
    LocalMux I__11328 (
            .O(N__47573),
            .I(N__47561));
    Span4Mux_v I__11327 (
            .O(N__47570),
            .I(N__47558));
    Span4Mux_h I__11326 (
            .O(N__47567),
            .I(N__47555));
    Span4Mux_v I__11325 (
            .O(N__47564),
            .I(N__47552));
    Span4Mux_v I__11324 (
            .O(N__47561),
            .I(N__47547));
    Span4Mux_h I__11323 (
            .O(N__47558),
            .I(N__47547));
    Odrv4 I__11322 (
            .O(N__47555),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13 ));
    Odrv4 I__11321 (
            .O(N__47552),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13 ));
    Odrv4 I__11320 (
            .O(N__47547),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13 ));
    InMux I__11319 (
            .O(N__47540),
            .I(N__47531));
    InMux I__11318 (
            .O(N__47539),
            .I(N__47527));
    InMux I__11317 (
            .O(N__47538),
            .I(N__47524));
    InMux I__11316 (
            .O(N__47537),
            .I(N__47521));
    InMux I__11315 (
            .O(N__47536),
            .I(N__47513));
    InMux I__11314 (
            .O(N__47535),
            .I(N__47513));
    InMux I__11313 (
            .O(N__47534),
            .I(N__47513));
    LocalMux I__11312 (
            .O(N__47531),
            .I(N__47510));
    InMux I__11311 (
            .O(N__47530),
            .I(N__47507));
    LocalMux I__11310 (
            .O(N__47527),
            .I(N__47502));
    LocalMux I__11309 (
            .O(N__47524),
            .I(N__47502));
    LocalMux I__11308 (
            .O(N__47521),
            .I(N__47499));
    InMux I__11307 (
            .O(N__47520),
            .I(N__47496));
    LocalMux I__11306 (
            .O(N__47513),
            .I(N__47493));
    Span4Mux_h I__11305 (
            .O(N__47510),
            .I(N__47488));
    LocalMux I__11304 (
            .O(N__47507),
            .I(N__47488));
    Span4Mux_v I__11303 (
            .O(N__47502),
            .I(N__47484));
    Span4Mux_h I__11302 (
            .O(N__47499),
            .I(N__47481));
    LocalMux I__11301 (
            .O(N__47496),
            .I(N__47478));
    Span4Mux_v I__11300 (
            .O(N__47493),
            .I(N__47475));
    Span4Mux_v I__11299 (
            .O(N__47488),
            .I(N__47472));
    InMux I__11298 (
            .O(N__47487),
            .I(N__47469));
    Span4Mux_v I__11297 (
            .O(N__47484),
            .I(N__47466));
    Span4Mux_v I__11296 (
            .O(N__47481),
            .I(N__47463));
    Span4Mux_h I__11295 (
            .O(N__47478),
            .I(N__47456));
    Span4Mux_v I__11294 (
            .O(N__47475),
            .I(N__47456));
    Span4Mux_v I__11293 (
            .O(N__47472),
            .I(N__47456));
    LocalMux I__11292 (
            .O(N__47469),
            .I(measured_delay_tr_15));
    Odrv4 I__11291 (
            .O(N__47466),
            .I(measured_delay_tr_15));
    Odrv4 I__11290 (
            .O(N__47463),
            .I(measured_delay_tr_15));
    Odrv4 I__11289 (
            .O(N__47456),
            .I(measured_delay_tr_15));
    CascadeMux I__11288 (
            .O(N__47447),
            .I(N__47444));
    InMux I__11287 (
            .O(N__47444),
            .I(N__47439));
    InMux I__11286 (
            .O(N__47443),
            .I(N__47436));
    CascadeMux I__11285 (
            .O(N__47442),
            .I(N__47432));
    LocalMux I__11284 (
            .O(N__47439),
            .I(N__47429));
    LocalMux I__11283 (
            .O(N__47436),
            .I(N__47426));
    InMux I__11282 (
            .O(N__47435),
            .I(N__47421));
    InMux I__11281 (
            .O(N__47432),
            .I(N__47421));
    Span4Mux_v I__11280 (
            .O(N__47429),
            .I(N__47418));
    Span4Mux_h I__11279 (
            .O(N__47426),
            .I(N__47413));
    LocalMux I__11278 (
            .O(N__47421),
            .I(N__47413));
    Span4Mux_h I__11277 (
            .O(N__47418),
            .I(N__47410));
    Span4Mux_v I__11276 (
            .O(N__47413),
            .I(N__47407));
    Odrv4 I__11275 (
            .O(N__47410),
            .I(measured_delay_tr_9));
    Odrv4 I__11274 (
            .O(N__47407),
            .I(measured_delay_tr_9));
    InMux I__11273 (
            .O(N__47402),
            .I(N__47397));
    InMux I__11272 (
            .O(N__47401),
            .I(N__47392));
    InMux I__11271 (
            .O(N__47400),
            .I(N__47392));
    LocalMux I__11270 (
            .O(N__47397),
            .I(N__47387));
    LocalMux I__11269 (
            .O(N__47392),
            .I(N__47384));
    InMux I__11268 (
            .O(N__47391),
            .I(N__47379));
    InMux I__11267 (
            .O(N__47390),
            .I(N__47379));
    Span4Mux_v I__11266 (
            .O(N__47387),
            .I(N__47376));
    Span4Mux_v I__11265 (
            .O(N__47384),
            .I(N__47371));
    LocalMux I__11264 (
            .O(N__47379),
            .I(N__47371));
    Span4Mux_h I__11263 (
            .O(N__47376),
            .I(N__47366));
    Span4Mux_h I__11262 (
            .O(N__47371),
            .I(N__47366));
    Odrv4 I__11261 (
            .O(N__47366),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0Z0Z_6 ));
    CascadeMux I__11260 (
            .O(N__47363),
            .I(N__47360));
    InMux I__11259 (
            .O(N__47360),
            .I(N__47357));
    LocalMux I__11258 (
            .O(N__47357),
            .I(N__47354));
    Odrv12 I__11257 (
            .O(N__47354),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ));
    ClkMux I__11256 (
            .O(N__47351),
            .I(N__46862));
    ClkMux I__11255 (
            .O(N__47350),
            .I(N__46862));
    ClkMux I__11254 (
            .O(N__47349),
            .I(N__46862));
    ClkMux I__11253 (
            .O(N__47348),
            .I(N__46862));
    ClkMux I__11252 (
            .O(N__47347),
            .I(N__46862));
    ClkMux I__11251 (
            .O(N__47346),
            .I(N__46862));
    ClkMux I__11250 (
            .O(N__47345),
            .I(N__46862));
    ClkMux I__11249 (
            .O(N__47344),
            .I(N__46862));
    ClkMux I__11248 (
            .O(N__47343),
            .I(N__46862));
    ClkMux I__11247 (
            .O(N__47342),
            .I(N__46862));
    ClkMux I__11246 (
            .O(N__47341),
            .I(N__46862));
    ClkMux I__11245 (
            .O(N__47340),
            .I(N__46862));
    ClkMux I__11244 (
            .O(N__47339),
            .I(N__46862));
    ClkMux I__11243 (
            .O(N__47338),
            .I(N__46862));
    ClkMux I__11242 (
            .O(N__47337),
            .I(N__46862));
    ClkMux I__11241 (
            .O(N__47336),
            .I(N__46862));
    ClkMux I__11240 (
            .O(N__47335),
            .I(N__46862));
    ClkMux I__11239 (
            .O(N__47334),
            .I(N__46862));
    ClkMux I__11238 (
            .O(N__47333),
            .I(N__46862));
    ClkMux I__11237 (
            .O(N__47332),
            .I(N__46862));
    ClkMux I__11236 (
            .O(N__47331),
            .I(N__46862));
    ClkMux I__11235 (
            .O(N__47330),
            .I(N__46862));
    ClkMux I__11234 (
            .O(N__47329),
            .I(N__46862));
    ClkMux I__11233 (
            .O(N__47328),
            .I(N__46862));
    ClkMux I__11232 (
            .O(N__47327),
            .I(N__46862));
    ClkMux I__11231 (
            .O(N__47326),
            .I(N__46862));
    ClkMux I__11230 (
            .O(N__47325),
            .I(N__46862));
    ClkMux I__11229 (
            .O(N__47324),
            .I(N__46862));
    ClkMux I__11228 (
            .O(N__47323),
            .I(N__46862));
    ClkMux I__11227 (
            .O(N__47322),
            .I(N__46862));
    ClkMux I__11226 (
            .O(N__47321),
            .I(N__46862));
    ClkMux I__11225 (
            .O(N__47320),
            .I(N__46862));
    ClkMux I__11224 (
            .O(N__47319),
            .I(N__46862));
    ClkMux I__11223 (
            .O(N__47318),
            .I(N__46862));
    ClkMux I__11222 (
            .O(N__47317),
            .I(N__46862));
    ClkMux I__11221 (
            .O(N__47316),
            .I(N__46862));
    ClkMux I__11220 (
            .O(N__47315),
            .I(N__46862));
    ClkMux I__11219 (
            .O(N__47314),
            .I(N__46862));
    ClkMux I__11218 (
            .O(N__47313),
            .I(N__46862));
    ClkMux I__11217 (
            .O(N__47312),
            .I(N__46862));
    ClkMux I__11216 (
            .O(N__47311),
            .I(N__46862));
    ClkMux I__11215 (
            .O(N__47310),
            .I(N__46862));
    ClkMux I__11214 (
            .O(N__47309),
            .I(N__46862));
    ClkMux I__11213 (
            .O(N__47308),
            .I(N__46862));
    ClkMux I__11212 (
            .O(N__47307),
            .I(N__46862));
    ClkMux I__11211 (
            .O(N__47306),
            .I(N__46862));
    ClkMux I__11210 (
            .O(N__47305),
            .I(N__46862));
    ClkMux I__11209 (
            .O(N__47304),
            .I(N__46862));
    ClkMux I__11208 (
            .O(N__47303),
            .I(N__46862));
    ClkMux I__11207 (
            .O(N__47302),
            .I(N__46862));
    ClkMux I__11206 (
            .O(N__47301),
            .I(N__46862));
    ClkMux I__11205 (
            .O(N__47300),
            .I(N__46862));
    ClkMux I__11204 (
            .O(N__47299),
            .I(N__46862));
    ClkMux I__11203 (
            .O(N__47298),
            .I(N__46862));
    ClkMux I__11202 (
            .O(N__47297),
            .I(N__46862));
    ClkMux I__11201 (
            .O(N__47296),
            .I(N__46862));
    ClkMux I__11200 (
            .O(N__47295),
            .I(N__46862));
    ClkMux I__11199 (
            .O(N__47294),
            .I(N__46862));
    ClkMux I__11198 (
            .O(N__47293),
            .I(N__46862));
    ClkMux I__11197 (
            .O(N__47292),
            .I(N__46862));
    ClkMux I__11196 (
            .O(N__47291),
            .I(N__46862));
    ClkMux I__11195 (
            .O(N__47290),
            .I(N__46862));
    ClkMux I__11194 (
            .O(N__47289),
            .I(N__46862));
    ClkMux I__11193 (
            .O(N__47288),
            .I(N__46862));
    ClkMux I__11192 (
            .O(N__47287),
            .I(N__46862));
    ClkMux I__11191 (
            .O(N__47286),
            .I(N__46862));
    ClkMux I__11190 (
            .O(N__47285),
            .I(N__46862));
    ClkMux I__11189 (
            .O(N__47284),
            .I(N__46862));
    ClkMux I__11188 (
            .O(N__47283),
            .I(N__46862));
    ClkMux I__11187 (
            .O(N__47282),
            .I(N__46862));
    ClkMux I__11186 (
            .O(N__47281),
            .I(N__46862));
    ClkMux I__11185 (
            .O(N__47280),
            .I(N__46862));
    ClkMux I__11184 (
            .O(N__47279),
            .I(N__46862));
    ClkMux I__11183 (
            .O(N__47278),
            .I(N__46862));
    ClkMux I__11182 (
            .O(N__47277),
            .I(N__46862));
    ClkMux I__11181 (
            .O(N__47276),
            .I(N__46862));
    ClkMux I__11180 (
            .O(N__47275),
            .I(N__46862));
    ClkMux I__11179 (
            .O(N__47274),
            .I(N__46862));
    ClkMux I__11178 (
            .O(N__47273),
            .I(N__46862));
    ClkMux I__11177 (
            .O(N__47272),
            .I(N__46862));
    ClkMux I__11176 (
            .O(N__47271),
            .I(N__46862));
    ClkMux I__11175 (
            .O(N__47270),
            .I(N__46862));
    ClkMux I__11174 (
            .O(N__47269),
            .I(N__46862));
    ClkMux I__11173 (
            .O(N__47268),
            .I(N__46862));
    ClkMux I__11172 (
            .O(N__47267),
            .I(N__46862));
    ClkMux I__11171 (
            .O(N__47266),
            .I(N__46862));
    ClkMux I__11170 (
            .O(N__47265),
            .I(N__46862));
    ClkMux I__11169 (
            .O(N__47264),
            .I(N__46862));
    ClkMux I__11168 (
            .O(N__47263),
            .I(N__46862));
    ClkMux I__11167 (
            .O(N__47262),
            .I(N__46862));
    ClkMux I__11166 (
            .O(N__47261),
            .I(N__46862));
    ClkMux I__11165 (
            .O(N__47260),
            .I(N__46862));
    ClkMux I__11164 (
            .O(N__47259),
            .I(N__46862));
    ClkMux I__11163 (
            .O(N__47258),
            .I(N__46862));
    ClkMux I__11162 (
            .O(N__47257),
            .I(N__46862));
    ClkMux I__11161 (
            .O(N__47256),
            .I(N__46862));
    ClkMux I__11160 (
            .O(N__47255),
            .I(N__46862));
    ClkMux I__11159 (
            .O(N__47254),
            .I(N__46862));
    ClkMux I__11158 (
            .O(N__47253),
            .I(N__46862));
    ClkMux I__11157 (
            .O(N__47252),
            .I(N__46862));
    ClkMux I__11156 (
            .O(N__47251),
            .I(N__46862));
    ClkMux I__11155 (
            .O(N__47250),
            .I(N__46862));
    ClkMux I__11154 (
            .O(N__47249),
            .I(N__46862));
    ClkMux I__11153 (
            .O(N__47248),
            .I(N__46862));
    ClkMux I__11152 (
            .O(N__47247),
            .I(N__46862));
    ClkMux I__11151 (
            .O(N__47246),
            .I(N__46862));
    ClkMux I__11150 (
            .O(N__47245),
            .I(N__46862));
    ClkMux I__11149 (
            .O(N__47244),
            .I(N__46862));
    ClkMux I__11148 (
            .O(N__47243),
            .I(N__46862));
    ClkMux I__11147 (
            .O(N__47242),
            .I(N__46862));
    ClkMux I__11146 (
            .O(N__47241),
            .I(N__46862));
    ClkMux I__11145 (
            .O(N__47240),
            .I(N__46862));
    ClkMux I__11144 (
            .O(N__47239),
            .I(N__46862));
    ClkMux I__11143 (
            .O(N__47238),
            .I(N__46862));
    ClkMux I__11142 (
            .O(N__47237),
            .I(N__46862));
    ClkMux I__11141 (
            .O(N__47236),
            .I(N__46862));
    ClkMux I__11140 (
            .O(N__47235),
            .I(N__46862));
    ClkMux I__11139 (
            .O(N__47234),
            .I(N__46862));
    ClkMux I__11138 (
            .O(N__47233),
            .I(N__46862));
    ClkMux I__11137 (
            .O(N__47232),
            .I(N__46862));
    ClkMux I__11136 (
            .O(N__47231),
            .I(N__46862));
    ClkMux I__11135 (
            .O(N__47230),
            .I(N__46862));
    ClkMux I__11134 (
            .O(N__47229),
            .I(N__46862));
    ClkMux I__11133 (
            .O(N__47228),
            .I(N__46862));
    ClkMux I__11132 (
            .O(N__47227),
            .I(N__46862));
    ClkMux I__11131 (
            .O(N__47226),
            .I(N__46862));
    ClkMux I__11130 (
            .O(N__47225),
            .I(N__46862));
    ClkMux I__11129 (
            .O(N__47224),
            .I(N__46862));
    ClkMux I__11128 (
            .O(N__47223),
            .I(N__46862));
    ClkMux I__11127 (
            .O(N__47222),
            .I(N__46862));
    ClkMux I__11126 (
            .O(N__47221),
            .I(N__46862));
    ClkMux I__11125 (
            .O(N__47220),
            .I(N__46862));
    ClkMux I__11124 (
            .O(N__47219),
            .I(N__46862));
    ClkMux I__11123 (
            .O(N__47218),
            .I(N__46862));
    ClkMux I__11122 (
            .O(N__47217),
            .I(N__46862));
    ClkMux I__11121 (
            .O(N__47216),
            .I(N__46862));
    ClkMux I__11120 (
            .O(N__47215),
            .I(N__46862));
    ClkMux I__11119 (
            .O(N__47214),
            .I(N__46862));
    ClkMux I__11118 (
            .O(N__47213),
            .I(N__46862));
    ClkMux I__11117 (
            .O(N__47212),
            .I(N__46862));
    ClkMux I__11116 (
            .O(N__47211),
            .I(N__46862));
    ClkMux I__11115 (
            .O(N__47210),
            .I(N__46862));
    ClkMux I__11114 (
            .O(N__47209),
            .I(N__46862));
    ClkMux I__11113 (
            .O(N__47208),
            .I(N__46862));
    ClkMux I__11112 (
            .O(N__47207),
            .I(N__46862));
    ClkMux I__11111 (
            .O(N__47206),
            .I(N__46862));
    ClkMux I__11110 (
            .O(N__47205),
            .I(N__46862));
    ClkMux I__11109 (
            .O(N__47204),
            .I(N__46862));
    ClkMux I__11108 (
            .O(N__47203),
            .I(N__46862));
    ClkMux I__11107 (
            .O(N__47202),
            .I(N__46862));
    ClkMux I__11106 (
            .O(N__47201),
            .I(N__46862));
    ClkMux I__11105 (
            .O(N__47200),
            .I(N__46862));
    ClkMux I__11104 (
            .O(N__47199),
            .I(N__46862));
    ClkMux I__11103 (
            .O(N__47198),
            .I(N__46862));
    ClkMux I__11102 (
            .O(N__47197),
            .I(N__46862));
    ClkMux I__11101 (
            .O(N__47196),
            .I(N__46862));
    ClkMux I__11100 (
            .O(N__47195),
            .I(N__46862));
    ClkMux I__11099 (
            .O(N__47194),
            .I(N__46862));
    ClkMux I__11098 (
            .O(N__47193),
            .I(N__46862));
    ClkMux I__11097 (
            .O(N__47192),
            .I(N__46862));
    ClkMux I__11096 (
            .O(N__47191),
            .I(N__46862));
    ClkMux I__11095 (
            .O(N__47190),
            .I(N__46862));
    ClkMux I__11094 (
            .O(N__47189),
            .I(N__46862));
    GlobalMux I__11093 (
            .O(N__46862),
            .I(clk_100mhz_0));
    CEMux I__11092 (
            .O(N__46859),
            .I(N__46853));
    CEMux I__11091 (
            .O(N__46858),
            .I(N__46849));
    CEMux I__11090 (
            .O(N__46857),
            .I(N__46846));
    CEMux I__11089 (
            .O(N__46856),
            .I(N__46843));
    LocalMux I__11088 (
            .O(N__46853),
            .I(N__46840));
    CEMux I__11087 (
            .O(N__46852),
            .I(N__46837));
    LocalMux I__11086 (
            .O(N__46849),
            .I(N__46834));
    LocalMux I__11085 (
            .O(N__46846),
            .I(N__46831));
    LocalMux I__11084 (
            .O(N__46843),
            .I(N__46828));
    Span4Mux_v I__11083 (
            .O(N__46840),
            .I(N__46823));
    LocalMux I__11082 (
            .O(N__46837),
            .I(N__46820));
    Span4Mux_v I__11081 (
            .O(N__46834),
            .I(N__46817));
    Span4Mux_h I__11080 (
            .O(N__46831),
            .I(N__46812));
    Span4Mux_h I__11079 (
            .O(N__46828),
            .I(N__46812));
    CEMux I__11078 (
            .O(N__46827),
            .I(N__46809));
    CEMux I__11077 (
            .O(N__46826),
            .I(N__46806));
    Span4Mux_h I__11076 (
            .O(N__46823),
            .I(N__46801));
    Span4Mux_v I__11075 (
            .O(N__46820),
            .I(N__46801));
    Span4Mux_h I__11074 (
            .O(N__46817),
            .I(N__46796));
    Span4Mux_h I__11073 (
            .O(N__46812),
            .I(N__46796));
    LocalMux I__11072 (
            .O(N__46809),
            .I(N__46793));
    LocalMux I__11071 (
            .O(N__46806),
            .I(N__46790));
    Odrv4 I__11070 (
            .O(N__46801),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv4 I__11069 (
            .O(N__46796),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv4 I__11068 (
            .O(N__46793),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv12 I__11067 (
            .O(N__46790),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ));
    CascadeMux I__11066 (
            .O(N__46781),
            .I(N__46774));
    InMux I__11065 (
            .O(N__46780),
            .I(N__46770));
    InMux I__11064 (
            .O(N__46779),
            .I(N__46767));
    InMux I__11063 (
            .O(N__46778),
            .I(N__46764));
    InMux I__11062 (
            .O(N__46777),
            .I(N__46761));
    InMux I__11061 (
            .O(N__46774),
            .I(N__46758));
    InMux I__11060 (
            .O(N__46773),
            .I(N__46755));
    LocalMux I__11059 (
            .O(N__46770),
            .I(N__46752));
    LocalMux I__11058 (
            .O(N__46767),
            .I(N__46749));
    LocalMux I__11057 (
            .O(N__46764),
            .I(N__46746));
    LocalMux I__11056 (
            .O(N__46761),
            .I(N__46698));
    LocalMux I__11055 (
            .O(N__46758),
            .I(N__46624));
    LocalMux I__11054 (
            .O(N__46755),
            .I(N__46621));
    Glb2LocalMux I__11053 (
            .O(N__46752),
            .I(N__46298));
    Glb2LocalMux I__11052 (
            .O(N__46749),
            .I(N__46298));
    Glb2LocalMux I__11051 (
            .O(N__46746),
            .I(N__46298));
    SRMux I__11050 (
            .O(N__46745),
            .I(N__46298));
    SRMux I__11049 (
            .O(N__46744),
            .I(N__46298));
    SRMux I__11048 (
            .O(N__46743),
            .I(N__46298));
    SRMux I__11047 (
            .O(N__46742),
            .I(N__46298));
    SRMux I__11046 (
            .O(N__46741),
            .I(N__46298));
    SRMux I__11045 (
            .O(N__46740),
            .I(N__46298));
    SRMux I__11044 (
            .O(N__46739),
            .I(N__46298));
    SRMux I__11043 (
            .O(N__46738),
            .I(N__46298));
    SRMux I__11042 (
            .O(N__46737),
            .I(N__46298));
    SRMux I__11041 (
            .O(N__46736),
            .I(N__46298));
    SRMux I__11040 (
            .O(N__46735),
            .I(N__46298));
    SRMux I__11039 (
            .O(N__46734),
            .I(N__46298));
    SRMux I__11038 (
            .O(N__46733),
            .I(N__46298));
    SRMux I__11037 (
            .O(N__46732),
            .I(N__46298));
    SRMux I__11036 (
            .O(N__46731),
            .I(N__46298));
    SRMux I__11035 (
            .O(N__46730),
            .I(N__46298));
    SRMux I__11034 (
            .O(N__46729),
            .I(N__46298));
    SRMux I__11033 (
            .O(N__46728),
            .I(N__46298));
    SRMux I__11032 (
            .O(N__46727),
            .I(N__46298));
    SRMux I__11031 (
            .O(N__46726),
            .I(N__46298));
    SRMux I__11030 (
            .O(N__46725),
            .I(N__46298));
    SRMux I__11029 (
            .O(N__46724),
            .I(N__46298));
    SRMux I__11028 (
            .O(N__46723),
            .I(N__46298));
    SRMux I__11027 (
            .O(N__46722),
            .I(N__46298));
    SRMux I__11026 (
            .O(N__46721),
            .I(N__46298));
    SRMux I__11025 (
            .O(N__46720),
            .I(N__46298));
    SRMux I__11024 (
            .O(N__46719),
            .I(N__46298));
    SRMux I__11023 (
            .O(N__46718),
            .I(N__46298));
    SRMux I__11022 (
            .O(N__46717),
            .I(N__46298));
    SRMux I__11021 (
            .O(N__46716),
            .I(N__46298));
    SRMux I__11020 (
            .O(N__46715),
            .I(N__46298));
    SRMux I__11019 (
            .O(N__46714),
            .I(N__46298));
    SRMux I__11018 (
            .O(N__46713),
            .I(N__46298));
    SRMux I__11017 (
            .O(N__46712),
            .I(N__46298));
    SRMux I__11016 (
            .O(N__46711),
            .I(N__46298));
    SRMux I__11015 (
            .O(N__46710),
            .I(N__46298));
    SRMux I__11014 (
            .O(N__46709),
            .I(N__46298));
    SRMux I__11013 (
            .O(N__46708),
            .I(N__46298));
    SRMux I__11012 (
            .O(N__46707),
            .I(N__46298));
    SRMux I__11011 (
            .O(N__46706),
            .I(N__46298));
    SRMux I__11010 (
            .O(N__46705),
            .I(N__46298));
    SRMux I__11009 (
            .O(N__46704),
            .I(N__46298));
    SRMux I__11008 (
            .O(N__46703),
            .I(N__46298));
    SRMux I__11007 (
            .O(N__46702),
            .I(N__46298));
    SRMux I__11006 (
            .O(N__46701),
            .I(N__46298));
    Glb2LocalMux I__11005 (
            .O(N__46698),
            .I(N__46298));
    SRMux I__11004 (
            .O(N__46697),
            .I(N__46298));
    SRMux I__11003 (
            .O(N__46696),
            .I(N__46298));
    SRMux I__11002 (
            .O(N__46695),
            .I(N__46298));
    SRMux I__11001 (
            .O(N__46694),
            .I(N__46298));
    SRMux I__11000 (
            .O(N__46693),
            .I(N__46298));
    SRMux I__10999 (
            .O(N__46692),
            .I(N__46298));
    SRMux I__10998 (
            .O(N__46691),
            .I(N__46298));
    SRMux I__10997 (
            .O(N__46690),
            .I(N__46298));
    SRMux I__10996 (
            .O(N__46689),
            .I(N__46298));
    SRMux I__10995 (
            .O(N__46688),
            .I(N__46298));
    SRMux I__10994 (
            .O(N__46687),
            .I(N__46298));
    SRMux I__10993 (
            .O(N__46686),
            .I(N__46298));
    SRMux I__10992 (
            .O(N__46685),
            .I(N__46298));
    SRMux I__10991 (
            .O(N__46684),
            .I(N__46298));
    SRMux I__10990 (
            .O(N__46683),
            .I(N__46298));
    SRMux I__10989 (
            .O(N__46682),
            .I(N__46298));
    SRMux I__10988 (
            .O(N__46681),
            .I(N__46298));
    SRMux I__10987 (
            .O(N__46680),
            .I(N__46298));
    SRMux I__10986 (
            .O(N__46679),
            .I(N__46298));
    SRMux I__10985 (
            .O(N__46678),
            .I(N__46298));
    SRMux I__10984 (
            .O(N__46677),
            .I(N__46298));
    SRMux I__10983 (
            .O(N__46676),
            .I(N__46298));
    SRMux I__10982 (
            .O(N__46675),
            .I(N__46298));
    SRMux I__10981 (
            .O(N__46674),
            .I(N__46298));
    SRMux I__10980 (
            .O(N__46673),
            .I(N__46298));
    SRMux I__10979 (
            .O(N__46672),
            .I(N__46298));
    SRMux I__10978 (
            .O(N__46671),
            .I(N__46298));
    SRMux I__10977 (
            .O(N__46670),
            .I(N__46298));
    SRMux I__10976 (
            .O(N__46669),
            .I(N__46298));
    SRMux I__10975 (
            .O(N__46668),
            .I(N__46298));
    SRMux I__10974 (
            .O(N__46667),
            .I(N__46298));
    SRMux I__10973 (
            .O(N__46666),
            .I(N__46298));
    SRMux I__10972 (
            .O(N__46665),
            .I(N__46298));
    SRMux I__10971 (
            .O(N__46664),
            .I(N__46298));
    SRMux I__10970 (
            .O(N__46663),
            .I(N__46298));
    SRMux I__10969 (
            .O(N__46662),
            .I(N__46298));
    SRMux I__10968 (
            .O(N__46661),
            .I(N__46298));
    SRMux I__10967 (
            .O(N__46660),
            .I(N__46298));
    SRMux I__10966 (
            .O(N__46659),
            .I(N__46298));
    SRMux I__10965 (
            .O(N__46658),
            .I(N__46298));
    SRMux I__10964 (
            .O(N__46657),
            .I(N__46298));
    SRMux I__10963 (
            .O(N__46656),
            .I(N__46298));
    SRMux I__10962 (
            .O(N__46655),
            .I(N__46298));
    SRMux I__10961 (
            .O(N__46654),
            .I(N__46298));
    SRMux I__10960 (
            .O(N__46653),
            .I(N__46298));
    SRMux I__10959 (
            .O(N__46652),
            .I(N__46298));
    SRMux I__10958 (
            .O(N__46651),
            .I(N__46298));
    SRMux I__10957 (
            .O(N__46650),
            .I(N__46298));
    SRMux I__10956 (
            .O(N__46649),
            .I(N__46298));
    SRMux I__10955 (
            .O(N__46648),
            .I(N__46298));
    SRMux I__10954 (
            .O(N__46647),
            .I(N__46298));
    SRMux I__10953 (
            .O(N__46646),
            .I(N__46298));
    SRMux I__10952 (
            .O(N__46645),
            .I(N__46298));
    SRMux I__10951 (
            .O(N__46644),
            .I(N__46298));
    SRMux I__10950 (
            .O(N__46643),
            .I(N__46298));
    SRMux I__10949 (
            .O(N__46642),
            .I(N__46298));
    SRMux I__10948 (
            .O(N__46641),
            .I(N__46298));
    SRMux I__10947 (
            .O(N__46640),
            .I(N__46298));
    SRMux I__10946 (
            .O(N__46639),
            .I(N__46298));
    SRMux I__10945 (
            .O(N__46638),
            .I(N__46298));
    SRMux I__10944 (
            .O(N__46637),
            .I(N__46298));
    SRMux I__10943 (
            .O(N__46636),
            .I(N__46298));
    SRMux I__10942 (
            .O(N__46635),
            .I(N__46298));
    SRMux I__10941 (
            .O(N__46634),
            .I(N__46298));
    SRMux I__10940 (
            .O(N__46633),
            .I(N__46298));
    SRMux I__10939 (
            .O(N__46632),
            .I(N__46298));
    SRMux I__10938 (
            .O(N__46631),
            .I(N__46298));
    SRMux I__10937 (
            .O(N__46630),
            .I(N__46298));
    SRMux I__10936 (
            .O(N__46629),
            .I(N__46298));
    SRMux I__10935 (
            .O(N__46628),
            .I(N__46298));
    SRMux I__10934 (
            .O(N__46627),
            .I(N__46298));
    Glb2LocalMux I__10933 (
            .O(N__46624),
            .I(N__46298));
    Glb2LocalMux I__10932 (
            .O(N__46621),
            .I(N__46298));
    SRMux I__10931 (
            .O(N__46620),
            .I(N__46298));
    SRMux I__10930 (
            .O(N__46619),
            .I(N__46298));
    SRMux I__10929 (
            .O(N__46618),
            .I(N__46298));
    SRMux I__10928 (
            .O(N__46617),
            .I(N__46298));
    SRMux I__10927 (
            .O(N__46616),
            .I(N__46298));
    SRMux I__10926 (
            .O(N__46615),
            .I(N__46298));
    SRMux I__10925 (
            .O(N__46614),
            .I(N__46298));
    SRMux I__10924 (
            .O(N__46613),
            .I(N__46298));
    SRMux I__10923 (
            .O(N__46612),
            .I(N__46298));
    SRMux I__10922 (
            .O(N__46611),
            .I(N__46298));
    SRMux I__10921 (
            .O(N__46610),
            .I(N__46298));
    SRMux I__10920 (
            .O(N__46609),
            .I(N__46298));
    SRMux I__10919 (
            .O(N__46608),
            .I(N__46298));
    SRMux I__10918 (
            .O(N__46607),
            .I(N__46298));
    SRMux I__10917 (
            .O(N__46606),
            .I(N__46298));
    SRMux I__10916 (
            .O(N__46605),
            .I(N__46298));
    SRMux I__10915 (
            .O(N__46604),
            .I(N__46298));
    SRMux I__10914 (
            .O(N__46603),
            .I(N__46298));
    SRMux I__10913 (
            .O(N__46602),
            .I(N__46298));
    SRMux I__10912 (
            .O(N__46601),
            .I(N__46298));
    SRMux I__10911 (
            .O(N__46600),
            .I(N__46298));
    SRMux I__10910 (
            .O(N__46599),
            .I(N__46298));
    SRMux I__10909 (
            .O(N__46598),
            .I(N__46298));
    SRMux I__10908 (
            .O(N__46597),
            .I(N__46298));
    SRMux I__10907 (
            .O(N__46596),
            .I(N__46298));
    SRMux I__10906 (
            .O(N__46595),
            .I(N__46298));
    GlobalMux I__10905 (
            .O(N__46298),
            .I(N__46295));
    gio2CtrlBuf I__10904 (
            .O(N__46295),
            .I(red_c_g));
    InMux I__10903 (
            .O(N__46292),
            .I(N__46288));
    InMux I__10902 (
            .O(N__46291),
            .I(N__46285));
    LocalMux I__10901 (
            .O(N__46288),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    LocalMux I__10900 (
            .O(N__46285),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__10899 (
            .O(N__46280),
            .I(N__46277));
    LocalMux I__10898 (
            .O(N__46277),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12 ));
    InMux I__10897 (
            .O(N__46274),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ));
    InMux I__10896 (
            .O(N__46271),
            .I(N__46267));
    InMux I__10895 (
            .O(N__46270),
            .I(N__46264));
    LocalMux I__10894 (
            .O(N__46267),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    LocalMux I__10893 (
            .O(N__46264),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__10892 (
            .O(N__46259),
            .I(N__46256));
    LocalMux I__10891 (
            .O(N__46256),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13 ));
    InMux I__10890 (
            .O(N__46253),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ));
    InMux I__10889 (
            .O(N__46250),
            .I(N__46246));
    InMux I__10888 (
            .O(N__46249),
            .I(N__46243));
    LocalMux I__10887 (
            .O(N__46246),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    LocalMux I__10886 (
            .O(N__46243),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__10885 (
            .O(N__46238),
            .I(N__46235));
    LocalMux I__10884 (
            .O(N__46235),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14 ));
    InMux I__10883 (
            .O(N__46232),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ));
    InMux I__10882 (
            .O(N__46229),
            .I(N__46226));
    LocalMux I__10881 (
            .O(N__46226),
            .I(N__46222));
    InMux I__10880 (
            .O(N__46225),
            .I(N__46219));
    Odrv4 I__10879 (
            .O(N__46222),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    LocalMux I__10878 (
            .O(N__46219),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__10877 (
            .O(N__46214),
            .I(N__46211));
    LocalMux I__10876 (
            .O(N__46211),
            .I(N__46208));
    Odrv4 I__10875 (
            .O(N__46208),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15 ));
    InMux I__10874 (
            .O(N__46205),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ));
    InMux I__10873 (
            .O(N__46202),
            .I(N__46198));
    InMux I__10872 (
            .O(N__46201),
            .I(N__46195));
    LocalMux I__10871 (
            .O(N__46198),
            .I(N__46192));
    LocalMux I__10870 (
            .O(N__46195),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv4 I__10869 (
            .O(N__46192),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    InMux I__10868 (
            .O(N__46187),
            .I(N__46184));
    LocalMux I__10867 (
            .O(N__46184),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16 ));
    InMux I__10866 (
            .O(N__46181),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ));
    InMux I__10865 (
            .O(N__46178),
            .I(N__46174));
    InMux I__10864 (
            .O(N__46177),
            .I(N__46171));
    LocalMux I__10863 (
            .O(N__46174),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    LocalMux I__10862 (
            .O(N__46171),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__10861 (
            .O(N__46166),
            .I(N__46163));
    LocalMux I__10860 (
            .O(N__46163),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17 ));
    InMux I__10859 (
            .O(N__46160),
            .I(bfn_18_19_0_));
    InMux I__10858 (
            .O(N__46157),
            .I(N__46153));
    InMux I__10857 (
            .O(N__46156),
            .I(N__46150));
    LocalMux I__10856 (
            .O(N__46153),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    LocalMux I__10855 (
            .O(N__46150),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__10854 (
            .O(N__46145),
            .I(N__46142));
    LocalMux I__10853 (
            .O(N__46142),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18 ));
    InMux I__10852 (
            .O(N__46139),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ));
    InMux I__10851 (
            .O(N__46136),
            .I(N__46132));
    InMux I__10850 (
            .O(N__46135),
            .I(N__46129));
    LocalMux I__10849 (
            .O(N__46132),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    LocalMux I__10848 (
            .O(N__46129),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__10847 (
            .O(N__46124),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17 ));
    InMux I__10846 (
            .O(N__46121),
            .I(N__46118));
    LocalMux I__10845 (
            .O(N__46118),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19 ));
    CascadeMux I__10844 (
            .O(N__46115),
            .I(N__46112));
    InMux I__10843 (
            .O(N__46112),
            .I(N__46108));
    InMux I__10842 (
            .O(N__46111),
            .I(N__46105));
    LocalMux I__10841 (
            .O(N__46108),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    LocalMux I__10840 (
            .O(N__46105),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__10839 (
            .O(N__46100),
            .I(N__46097));
    LocalMux I__10838 (
            .O(N__46097),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4 ));
    InMux I__10837 (
            .O(N__46094),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ));
    InMux I__10836 (
            .O(N__46091),
            .I(N__46087));
    InMux I__10835 (
            .O(N__46090),
            .I(N__46084));
    LocalMux I__10834 (
            .O(N__46087),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    LocalMux I__10833 (
            .O(N__46084),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__10832 (
            .O(N__46079),
            .I(N__46076));
    LocalMux I__10831 (
            .O(N__46076),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5 ));
    InMux I__10830 (
            .O(N__46073),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ));
    InMux I__10829 (
            .O(N__46070),
            .I(N__46066));
    InMux I__10828 (
            .O(N__46069),
            .I(N__46063));
    LocalMux I__10827 (
            .O(N__46066),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    LocalMux I__10826 (
            .O(N__46063),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__10825 (
            .O(N__46058),
            .I(N__46055));
    LocalMux I__10824 (
            .O(N__46055),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6 ));
    InMux I__10823 (
            .O(N__46052),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ));
    InMux I__10822 (
            .O(N__46049),
            .I(N__46045));
    InMux I__10821 (
            .O(N__46048),
            .I(N__46042));
    LocalMux I__10820 (
            .O(N__46045),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    LocalMux I__10819 (
            .O(N__46042),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__10818 (
            .O(N__46037),
            .I(N__46034));
    LocalMux I__10817 (
            .O(N__46034),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7 ));
    InMux I__10816 (
            .O(N__46031),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ));
    InMux I__10815 (
            .O(N__46028),
            .I(N__46024));
    InMux I__10814 (
            .O(N__46027),
            .I(N__46021));
    LocalMux I__10813 (
            .O(N__46024),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    LocalMux I__10812 (
            .O(N__46021),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__10811 (
            .O(N__46016),
            .I(N__46013));
    LocalMux I__10810 (
            .O(N__46013),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8 ));
    InMux I__10809 (
            .O(N__46010),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ));
    InMux I__10808 (
            .O(N__46007),
            .I(bfn_18_18_0_));
    InMux I__10807 (
            .O(N__46004),
            .I(N__46000));
    InMux I__10806 (
            .O(N__46003),
            .I(N__45997));
    LocalMux I__10805 (
            .O(N__46000),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    LocalMux I__10804 (
            .O(N__45997),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__10803 (
            .O(N__45992),
            .I(N__45989));
    LocalMux I__10802 (
            .O(N__45989),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10 ));
    InMux I__10801 (
            .O(N__45986),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ));
    InMux I__10800 (
            .O(N__45983),
            .I(N__45979));
    InMux I__10799 (
            .O(N__45982),
            .I(N__45976));
    LocalMux I__10798 (
            .O(N__45979),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    LocalMux I__10797 (
            .O(N__45976),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__10796 (
            .O(N__45971),
            .I(N__45968));
    LocalMux I__10795 (
            .O(N__45968),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11 ));
    InMux I__10794 (
            .O(N__45965),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ));
    InMux I__10793 (
            .O(N__45962),
            .I(N__45959));
    LocalMux I__10792 (
            .O(N__45959),
            .I(N__45955));
    CascadeMux I__10791 (
            .O(N__45958),
            .I(N__45951));
    Span4Mux_h I__10790 (
            .O(N__45955),
            .I(N__45948));
    InMux I__10789 (
            .O(N__45954),
            .I(N__45945));
    InMux I__10788 (
            .O(N__45951),
            .I(N__45942));
    Odrv4 I__10787 (
            .O(N__45948),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    LocalMux I__10786 (
            .O(N__45945),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    LocalMux I__10785 (
            .O(N__45942),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    CascadeMux I__10784 (
            .O(N__45935),
            .I(N__45932));
    InMux I__10783 (
            .O(N__45932),
            .I(N__45929));
    LocalMux I__10782 (
            .O(N__45929),
            .I(N__45926));
    Span4Mux_h I__10781 (
            .O(N__45926),
            .I(N__45923));
    Odrv4 I__10780 (
            .O(N__45923),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    InMux I__10779 (
            .O(N__45920),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__10778 (
            .O(N__45917),
            .I(N__45914));
    LocalMux I__10777 (
            .O(N__45914),
            .I(N__45910));
    InMux I__10776 (
            .O(N__45913),
            .I(N__45907));
    Span4Mux_h I__10775 (
            .O(N__45910),
            .I(N__45904));
    LocalMux I__10774 (
            .O(N__45907),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    Odrv4 I__10773 (
            .O(N__45904),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    CascadeMux I__10772 (
            .O(N__45899),
            .I(N__45895));
    CascadeMux I__10771 (
            .O(N__45898),
            .I(N__45892));
    InMux I__10770 (
            .O(N__45895),
            .I(N__45886));
    InMux I__10769 (
            .O(N__45892),
            .I(N__45886));
    InMux I__10768 (
            .O(N__45891),
            .I(N__45883));
    LocalMux I__10767 (
            .O(N__45886),
            .I(N__45880));
    LocalMux I__10766 (
            .O(N__45883),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    Odrv4 I__10765 (
            .O(N__45880),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    InMux I__10764 (
            .O(N__45875),
            .I(N__45872));
    LocalMux I__10763 (
            .O(N__45872),
            .I(N__45869));
    Span4Mux_v I__10762 (
            .O(N__45869),
            .I(N__45866));
    Odrv4 I__10761 (
            .O(N__45866),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    InMux I__10760 (
            .O(N__45863),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__10759 (
            .O(N__45860),
            .I(N__45856));
    InMux I__10758 (
            .O(N__45859),
            .I(N__45853));
    LocalMux I__10757 (
            .O(N__45856),
            .I(N__45850));
    LocalMux I__10756 (
            .O(N__45853),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    Odrv4 I__10755 (
            .O(N__45850),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    CascadeMux I__10754 (
            .O(N__45845),
            .I(N__45841));
    CascadeMux I__10753 (
            .O(N__45844),
            .I(N__45838));
    InMux I__10752 (
            .O(N__45841),
            .I(N__45832));
    InMux I__10751 (
            .O(N__45838),
            .I(N__45832));
    InMux I__10750 (
            .O(N__45837),
            .I(N__45829));
    LocalMux I__10749 (
            .O(N__45832),
            .I(N__45826));
    LocalMux I__10748 (
            .O(N__45829),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    Odrv4 I__10747 (
            .O(N__45826),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    InMux I__10746 (
            .O(N__45821),
            .I(N__45818));
    LocalMux I__10745 (
            .O(N__45818),
            .I(N__45815));
    Span4Mux_v I__10744 (
            .O(N__45815),
            .I(N__45812));
    Odrv4 I__10743 (
            .O(N__45812),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30 ));
    InMux I__10742 (
            .O(N__45809),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__10741 (
            .O(N__45806),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ));
    CascadeMux I__10740 (
            .O(N__45803),
            .I(N__45798));
    InMux I__10739 (
            .O(N__45802),
            .I(N__45791));
    CascadeMux I__10738 (
            .O(N__45801),
            .I(N__45787));
    InMux I__10737 (
            .O(N__45798),
            .I(N__45782));
    InMux I__10736 (
            .O(N__45797),
            .I(N__45773));
    InMux I__10735 (
            .O(N__45796),
            .I(N__45773));
    InMux I__10734 (
            .O(N__45795),
            .I(N__45773));
    InMux I__10733 (
            .O(N__45794),
            .I(N__45773));
    LocalMux I__10732 (
            .O(N__45791),
            .I(N__45770));
    InMux I__10731 (
            .O(N__45790),
            .I(N__45765));
    InMux I__10730 (
            .O(N__45787),
            .I(N__45765));
    CascadeMux I__10729 (
            .O(N__45786),
            .I(N__45762));
    InMux I__10728 (
            .O(N__45785),
            .I(N__45757));
    LocalMux I__10727 (
            .O(N__45782),
            .I(N__45748));
    LocalMux I__10726 (
            .O(N__45773),
            .I(N__45748));
    Span4Mux_h I__10725 (
            .O(N__45770),
            .I(N__45748));
    LocalMux I__10724 (
            .O(N__45765),
            .I(N__45748));
    InMux I__10723 (
            .O(N__45762),
            .I(N__45741));
    InMux I__10722 (
            .O(N__45761),
            .I(N__45741));
    InMux I__10721 (
            .O(N__45760),
            .I(N__45741));
    LocalMux I__10720 (
            .O(N__45757),
            .I(N__45736));
    Span4Mux_v I__10719 (
            .O(N__45748),
            .I(N__45736));
    LocalMux I__10718 (
            .O(N__45741),
            .I(\delay_measurement_inst.elapsed_time_tr_31 ));
    Odrv4 I__10717 (
            .O(N__45736),
            .I(\delay_measurement_inst.elapsed_time_tr_31 ));
    CEMux I__10716 (
            .O(N__45731),
            .I(N__45728));
    LocalMux I__10715 (
            .O(N__45728),
            .I(N__45722));
    CEMux I__10714 (
            .O(N__45727),
            .I(N__45719));
    CEMux I__10713 (
            .O(N__45726),
            .I(N__45715));
    CEMux I__10712 (
            .O(N__45725),
            .I(N__45712));
    Span4Mux_v I__10711 (
            .O(N__45722),
            .I(N__45707));
    LocalMux I__10710 (
            .O(N__45719),
            .I(N__45707));
    CEMux I__10709 (
            .O(N__45718),
            .I(N__45704));
    LocalMux I__10708 (
            .O(N__45715),
            .I(N__45698));
    LocalMux I__10707 (
            .O(N__45712),
            .I(N__45698));
    Span4Mux_v I__10706 (
            .O(N__45707),
            .I(N__45693));
    LocalMux I__10705 (
            .O(N__45704),
            .I(N__45693));
    CEMux I__10704 (
            .O(N__45703),
            .I(N__45690));
    Span4Mux_v I__10703 (
            .O(N__45698),
            .I(N__45687));
    Span4Mux_h I__10702 (
            .O(N__45693),
            .I(N__45684));
    LocalMux I__10701 (
            .O(N__45690),
            .I(N__45681));
    Odrv4 I__10700 (
            .O(N__45687),
            .I(\delay_measurement_inst.delay_tr_timer.N_323_i ));
    Odrv4 I__10699 (
            .O(N__45684),
            .I(\delay_measurement_inst.delay_tr_timer.N_323_i ));
    Odrv12 I__10698 (
            .O(N__45681),
            .I(\delay_measurement_inst.delay_tr_timer.N_323_i ));
    InMux I__10697 (
            .O(N__45674),
            .I(N__45671));
    LocalMux I__10696 (
            .O(N__45671),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0 ));
    CascadeMux I__10695 (
            .O(N__45668),
            .I(N__45665));
    InMux I__10694 (
            .O(N__45665),
            .I(N__45661));
    InMux I__10693 (
            .O(N__45664),
            .I(N__45657));
    LocalMux I__10692 (
            .O(N__45661),
            .I(N__45654));
    InMux I__10691 (
            .O(N__45660),
            .I(N__45651));
    LocalMux I__10690 (
            .O(N__45657),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv4 I__10689 (
            .O(N__45654),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__10688 (
            .O(N__45651),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    InMux I__10687 (
            .O(N__45644),
            .I(N__45640));
    InMux I__10686 (
            .O(N__45643),
            .I(N__45637));
    LocalMux I__10685 (
            .O(N__45640),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    LocalMux I__10684 (
            .O(N__45637),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__10683 (
            .O(N__45632),
            .I(N__45629));
    LocalMux I__10682 (
            .O(N__45629),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2 ));
    InMux I__10681 (
            .O(N__45626),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ));
    InMux I__10680 (
            .O(N__45623),
            .I(N__45620));
    LocalMux I__10679 (
            .O(N__45620),
            .I(N__45617));
    Odrv4 I__10678 (
            .O(N__45617),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0 ));
    CascadeMux I__10677 (
            .O(N__45614),
            .I(N__45611));
    InMux I__10676 (
            .O(N__45611),
            .I(N__45607));
    InMux I__10675 (
            .O(N__45610),
            .I(N__45604));
    LocalMux I__10674 (
            .O(N__45607),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    LocalMux I__10673 (
            .O(N__45604),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__10672 (
            .O(N__45599),
            .I(N__45596));
    LocalMux I__10671 (
            .O(N__45596),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3 ));
    InMux I__10670 (
            .O(N__45593),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ));
    CascadeMux I__10669 (
            .O(N__45590),
            .I(N__45587));
    InMux I__10668 (
            .O(N__45587),
            .I(N__45584));
    LocalMux I__10667 (
            .O(N__45584),
            .I(N__45580));
    InMux I__10666 (
            .O(N__45583),
            .I(N__45576));
    Span4Mux_h I__10665 (
            .O(N__45580),
            .I(N__45573));
    InMux I__10664 (
            .O(N__45579),
            .I(N__45570));
    LocalMux I__10663 (
            .O(N__45576),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    Odrv4 I__10662 (
            .O(N__45573),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    LocalMux I__10661 (
            .O(N__45570),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    InMux I__10660 (
            .O(N__45563),
            .I(N__45560));
    LocalMux I__10659 (
            .O(N__45560),
            .I(N__45557));
    Span4Mux_v I__10658 (
            .O(N__45557),
            .I(N__45554));
    Odrv4 I__10657 (
            .O(N__45554),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    InMux I__10656 (
            .O(N__45551),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ));
    CascadeMux I__10655 (
            .O(N__45548),
            .I(N__45544));
    InMux I__10654 (
            .O(N__45547),
            .I(N__45541));
    InMux I__10653 (
            .O(N__45544),
            .I(N__45538));
    LocalMux I__10652 (
            .O(N__45541),
            .I(N__45534));
    LocalMux I__10651 (
            .O(N__45538),
            .I(N__45531));
    InMux I__10650 (
            .O(N__45537),
            .I(N__45528));
    Span4Mux_v I__10649 (
            .O(N__45534),
            .I(N__45525));
    Span4Mux_v I__10648 (
            .O(N__45531),
            .I(N__45522));
    LocalMux I__10647 (
            .O(N__45528),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    Odrv4 I__10646 (
            .O(N__45525),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    Odrv4 I__10645 (
            .O(N__45522),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    InMux I__10644 (
            .O(N__45515),
            .I(N__45512));
    LocalMux I__10643 (
            .O(N__45512),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    InMux I__10642 (
            .O(N__45509),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__10641 (
            .O(N__45506),
            .I(N__45499));
    InMux I__10640 (
            .O(N__45505),
            .I(N__45499));
    InMux I__10639 (
            .O(N__45504),
            .I(N__45496));
    LocalMux I__10638 (
            .O(N__45499),
            .I(N__45493));
    LocalMux I__10637 (
            .O(N__45496),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    Odrv4 I__10636 (
            .O(N__45493),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    InMux I__10635 (
            .O(N__45488),
            .I(N__45485));
    LocalMux I__10634 (
            .O(N__45485),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    InMux I__10633 (
            .O(N__45482),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__10632 (
            .O(N__45479),
            .I(N__45475));
    CascadeMux I__10631 (
            .O(N__45478),
            .I(N__45472));
    InMux I__10630 (
            .O(N__45475),
            .I(N__45466));
    InMux I__10629 (
            .O(N__45472),
            .I(N__45466));
    InMux I__10628 (
            .O(N__45471),
            .I(N__45463));
    LocalMux I__10627 (
            .O(N__45466),
            .I(N__45460));
    LocalMux I__10626 (
            .O(N__45463),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    Odrv4 I__10625 (
            .O(N__45460),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    InMux I__10624 (
            .O(N__45455),
            .I(N__45452));
    LocalMux I__10623 (
            .O(N__45452),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    InMux I__10622 (
            .O(N__45449),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ));
    CascadeMux I__10621 (
            .O(N__45446),
            .I(N__45442));
    CascadeMux I__10620 (
            .O(N__45445),
            .I(N__45439));
    InMux I__10619 (
            .O(N__45442),
            .I(N__45433));
    InMux I__10618 (
            .O(N__45439),
            .I(N__45433));
    InMux I__10617 (
            .O(N__45438),
            .I(N__45430));
    LocalMux I__10616 (
            .O(N__45433),
            .I(N__45427));
    LocalMux I__10615 (
            .O(N__45430),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    Odrv4 I__10614 (
            .O(N__45427),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    CascadeMux I__10613 (
            .O(N__45422),
            .I(N__45419));
    InMux I__10612 (
            .O(N__45419),
            .I(N__45416));
    LocalMux I__10611 (
            .O(N__45416),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    InMux I__10610 (
            .O(N__45413),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ));
    InMux I__10609 (
            .O(N__45410),
            .I(N__45403));
    InMux I__10608 (
            .O(N__45409),
            .I(N__45403));
    InMux I__10607 (
            .O(N__45408),
            .I(N__45400));
    LocalMux I__10606 (
            .O(N__45403),
            .I(N__45397));
    LocalMux I__10605 (
            .O(N__45400),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    Odrv4 I__10604 (
            .O(N__45397),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    InMux I__10603 (
            .O(N__45392),
            .I(N__45389));
    LocalMux I__10602 (
            .O(N__45389),
            .I(N__45386));
    Span4Mux_h I__10601 (
            .O(N__45386),
            .I(N__45383));
    Odrv4 I__10600 (
            .O(N__45383),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    InMux I__10599 (
            .O(N__45380),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ));
    InMux I__10598 (
            .O(N__45377),
            .I(N__45371));
    InMux I__10597 (
            .O(N__45376),
            .I(N__45371));
    LocalMux I__10596 (
            .O(N__45371),
            .I(N__45367));
    InMux I__10595 (
            .O(N__45370),
            .I(N__45364));
    Span4Mux_v I__10594 (
            .O(N__45367),
            .I(N__45361));
    LocalMux I__10593 (
            .O(N__45364),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    Odrv4 I__10592 (
            .O(N__45361),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    InMux I__10591 (
            .O(N__45356),
            .I(N__45353));
    LocalMux I__10590 (
            .O(N__45353),
            .I(N__45350));
    Span4Mux_h I__10589 (
            .O(N__45350),
            .I(N__45347));
    Odrv4 I__10588 (
            .O(N__45347),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    InMux I__10587 (
            .O(N__45344),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ));
    InMux I__10586 (
            .O(N__45341),
            .I(N__45337));
    CascadeMux I__10585 (
            .O(N__45340),
            .I(N__45333));
    LocalMux I__10584 (
            .O(N__45337),
            .I(N__45330));
    InMux I__10583 (
            .O(N__45336),
            .I(N__45327));
    InMux I__10582 (
            .O(N__45333),
            .I(N__45324));
    Odrv4 I__10581 (
            .O(N__45330),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    LocalMux I__10580 (
            .O(N__45327),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    LocalMux I__10579 (
            .O(N__45324),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    InMux I__10578 (
            .O(N__45317),
            .I(N__45314));
    LocalMux I__10577 (
            .O(N__45314),
            .I(N__45311));
    Span4Mux_h I__10576 (
            .O(N__45311),
            .I(N__45308));
    Odrv4 I__10575 (
            .O(N__45308),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    InMux I__10574 (
            .O(N__45305),
            .I(bfn_18_16_0_));
    InMux I__10573 (
            .O(N__45302),
            .I(N__45299));
    LocalMux I__10572 (
            .O(N__45299),
            .I(N__45294));
    InMux I__10571 (
            .O(N__45298),
            .I(N__45291));
    InMux I__10570 (
            .O(N__45297),
            .I(N__45288));
    Odrv4 I__10569 (
            .O(N__45294),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    LocalMux I__10568 (
            .O(N__45291),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    LocalMux I__10567 (
            .O(N__45288),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    InMux I__10566 (
            .O(N__45281),
            .I(N__45278));
    LocalMux I__10565 (
            .O(N__45278),
            .I(N__45274));
    InMux I__10564 (
            .O(N__45277),
            .I(N__45271));
    Span4Mux_v I__10563 (
            .O(N__45274),
            .I(N__45266));
    LocalMux I__10562 (
            .O(N__45271),
            .I(N__45266));
    Odrv4 I__10561 (
            .O(N__45266),
            .I(\delay_measurement_inst.elapsed_time_tr_12 ));
    InMux I__10560 (
            .O(N__45263),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__10559 (
            .O(N__45260),
            .I(N__45256));
    CascadeMux I__10558 (
            .O(N__45259),
            .I(N__45253));
    InMux I__10557 (
            .O(N__45256),
            .I(N__45247));
    InMux I__10556 (
            .O(N__45253),
            .I(N__45247));
    InMux I__10555 (
            .O(N__45252),
            .I(N__45244));
    LocalMux I__10554 (
            .O(N__45247),
            .I(N__45241));
    LocalMux I__10553 (
            .O(N__45244),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    Odrv4 I__10552 (
            .O(N__45241),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    InMux I__10551 (
            .O(N__45236),
            .I(N__45232));
    CascadeMux I__10550 (
            .O(N__45235),
            .I(N__45229));
    LocalMux I__10549 (
            .O(N__45232),
            .I(N__45226));
    InMux I__10548 (
            .O(N__45229),
            .I(N__45223));
    Span4Mux_h I__10547 (
            .O(N__45226),
            .I(N__45220));
    LocalMux I__10546 (
            .O(N__45223),
            .I(N__45217));
    Odrv4 I__10545 (
            .O(N__45220),
            .I(\delay_measurement_inst.elapsed_time_tr_13 ));
    Odrv4 I__10544 (
            .O(N__45217),
            .I(\delay_measurement_inst.elapsed_time_tr_13 ));
    InMux I__10543 (
            .O(N__45212),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ));
    CascadeMux I__10542 (
            .O(N__45209),
            .I(N__45205));
    CascadeMux I__10541 (
            .O(N__45208),
            .I(N__45202));
    InMux I__10540 (
            .O(N__45205),
            .I(N__45196));
    InMux I__10539 (
            .O(N__45202),
            .I(N__45196));
    InMux I__10538 (
            .O(N__45201),
            .I(N__45193));
    LocalMux I__10537 (
            .O(N__45196),
            .I(N__45190));
    LocalMux I__10536 (
            .O(N__45193),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    Odrv4 I__10535 (
            .O(N__45190),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    InMux I__10534 (
            .O(N__45185),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ));
    InMux I__10533 (
            .O(N__45182),
            .I(N__45176));
    InMux I__10532 (
            .O(N__45181),
            .I(N__45176));
    LocalMux I__10531 (
            .O(N__45176),
            .I(N__45172));
    InMux I__10530 (
            .O(N__45175),
            .I(N__45169));
    Span4Mux_h I__10529 (
            .O(N__45172),
            .I(N__45166));
    LocalMux I__10528 (
            .O(N__45169),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    Odrv4 I__10527 (
            .O(N__45166),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    InMux I__10526 (
            .O(N__45161),
            .I(N__45156));
    CascadeMux I__10525 (
            .O(N__45160),
            .I(N__45150));
    InMux I__10524 (
            .O(N__45159),
            .I(N__45147));
    LocalMux I__10523 (
            .O(N__45156),
            .I(N__45144));
    InMux I__10522 (
            .O(N__45155),
            .I(N__45139));
    InMux I__10521 (
            .O(N__45154),
            .I(N__45139));
    InMux I__10520 (
            .O(N__45153),
            .I(N__45134));
    InMux I__10519 (
            .O(N__45150),
            .I(N__45134));
    LocalMux I__10518 (
            .O(N__45147),
            .I(N__45131));
    Span4Mux_v I__10517 (
            .O(N__45144),
            .I(N__45128));
    LocalMux I__10516 (
            .O(N__45139),
            .I(N__45125));
    LocalMux I__10515 (
            .O(N__45134),
            .I(N__45122));
    Span4Mux_v I__10514 (
            .O(N__45131),
            .I(N__45117));
    Span4Mux_h I__10513 (
            .O(N__45128),
            .I(N__45117));
    Span4Mux_h I__10512 (
            .O(N__45125),
            .I(N__45114));
    Span4Mux_h I__10511 (
            .O(N__45122),
            .I(N__45111));
    Odrv4 I__10510 (
            .O(N__45117),
            .I(\delay_measurement_inst.elapsed_time_tr_15 ));
    Odrv4 I__10509 (
            .O(N__45114),
            .I(\delay_measurement_inst.elapsed_time_tr_15 ));
    Odrv4 I__10508 (
            .O(N__45111),
            .I(\delay_measurement_inst.elapsed_time_tr_15 ));
    InMux I__10507 (
            .O(N__45104),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ));
    InMux I__10506 (
            .O(N__45101),
            .I(N__45095));
    InMux I__10505 (
            .O(N__45100),
            .I(N__45095));
    LocalMux I__10504 (
            .O(N__45095),
            .I(N__45091));
    InMux I__10503 (
            .O(N__45094),
            .I(N__45088));
    Span4Mux_h I__10502 (
            .O(N__45091),
            .I(N__45085));
    LocalMux I__10501 (
            .O(N__45088),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    Odrv4 I__10500 (
            .O(N__45085),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    InMux I__10499 (
            .O(N__45080),
            .I(N__45077));
    LocalMux I__10498 (
            .O(N__45077),
            .I(N__45072));
    InMux I__10497 (
            .O(N__45076),
            .I(N__45067));
    InMux I__10496 (
            .O(N__45075),
            .I(N__45067));
    Odrv4 I__10495 (
            .O(N__45072),
            .I(\delay_measurement_inst.elapsed_time_tr_16 ));
    LocalMux I__10494 (
            .O(N__45067),
            .I(\delay_measurement_inst.elapsed_time_tr_16 ));
    InMux I__10493 (
            .O(N__45062),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__10492 (
            .O(N__45059),
            .I(N__45056));
    InMux I__10491 (
            .O(N__45056),
            .I(N__45052));
    InMux I__10490 (
            .O(N__45055),
            .I(N__45048));
    LocalMux I__10489 (
            .O(N__45052),
            .I(N__45045));
    InMux I__10488 (
            .O(N__45051),
            .I(N__45042));
    LocalMux I__10487 (
            .O(N__45048),
            .I(N__45039));
    Span4Mux_h I__10486 (
            .O(N__45045),
            .I(N__45036));
    LocalMux I__10485 (
            .O(N__45042),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    Odrv4 I__10484 (
            .O(N__45039),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    Odrv4 I__10483 (
            .O(N__45036),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    InMux I__10482 (
            .O(N__45029),
            .I(N__45026));
    LocalMux I__10481 (
            .O(N__45026),
            .I(N__45021));
    InMux I__10480 (
            .O(N__45025),
            .I(N__45018));
    InMux I__10479 (
            .O(N__45024),
            .I(N__45015));
    Odrv4 I__10478 (
            .O(N__45021),
            .I(\delay_measurement_inst.elapsed_time_tr_17 ));
    LocalMux I__10477 (
            .O(N__45018),
            .I(\delay_measurement_inst.elapsed_time_tr_17 ));
    LocalMux I__10476 (
            .O(N__45015),
            .I(\delay_measurement_inst.elapsed_time_tr_17 ));
    InMux I__10475 (
            .O(N__45008),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ));
    CascadeMux I__10474 (
            .O(N__45005),
            .I(N__45001));
    CascadeMux I__10473 (
            .O(N__45004),
            .I(N__44998));
    InMux I__10472 (
            .O(N__45001),
            .I(N__44993));
    InMux I__10471 (
            .O(N__44998),
            .I(N__44993));
    LocalMux I__10470 (
            .O(N__44993),
            .I(N__44989));
    InMux I__10469 (
            .O(N__44992),
            .I(N__44986));
    Span4Mux_v I__10468 (
            .O(N__44989),
            .I(N__44983));
    LocalMux I__10467 (
            .O(N__44986),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    Odrv4 I__10466 (
            .O(N__44983),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    InMux I__10465 (
            .O(N__44978),
            .I(N__44975));
    LocalMux I__10464 (
            .O(N__44975),
            .I(N__44970));
    InMux I__10463 (
            .O(N__44974),
            .I(N__44965));
    InMux I__10462 (
            .O(N__44973),
            .I(N__44965));
    Odrv4 I__10461 (
            .O(N__44970),
            .I(\delay_measurement_inst.elapsed_time_tr_18 ));
    LocalMux I__10460 (
            .O(N__44965),
            .I(\delay_measurement_inst.elapsed_time_tr_18 ));
    InMux I__10459 (
            .O(N__44960),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ));
    InMux I__10458 (
            .O(N__44957),
            .I(N__44954));
    LocalMux I__10457 (
            .O(N__44954),
            .I(N__44950));
    CascadeMux I__10456 (
            .O(N__44953),
            .I(N__44946));
    Span4Mux_h I__10455 (
            .O(N__44950),
            .I(N__44943));
    InMux I__10454 (
            .O(N__44949),
            .I(N__44940));
    InMux I__10453 (
            .O(N__44946),
            .I(N__44937));
    Odrv4 I__10452 (
            .O(N__44943),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    LocalMux I__10451 (
            .O(N__44940),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    LocalMux I__10450 (
            .O(N__44937),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    InMux I__10449 (
            .O(N__44930),
            .I(N__44927));
    LocalMux I__10448 (
            .O(N__44927),
            .I(N__44922));
    CascadeMux I__10447 (
            .O(N__44926),
            .I(N__44919));
    CascadeMux I__10446 (
            .O(N__44925),
            .I(N__44916));
    Span4Mux_h I__10445 (
            .O(N__44922),
            .I(N__44913));
    InMux I__10444 (
            .O(N__44919),
            .I(N__44910));
    InMux I__10443 (
            .O(N__44916),
            .I(N__44907));
    Odrv4 I__10442 (
            .O(N__44913),
            .I(\delay_measurement_inst.elapsed_time_tr_19 ));
    LocalMux I__10441 (
            .O(N__44910),
            .I(\delay_measurement_inst.elapsed_time_tr_19 ));
    LocalMux I__10440 (
            .O(N__44907),
            .I(\delay_measurement_inst.elapsed_time_tr_19 ));
    InMux I__10439 (
            .O(N__44900),
            .I(bfn_18_15_0_));
    InMux I__10438 (
            .O(N__44897),
            .I(N__44894));
    LocalMux I__10437 (
            .O(N__44894),
            .I(N__44890));
    InMux I__10436 (
            .O(N__44893),
            .I(N__44886));
    Span4Mux_v I__10435 (
            .O(N__44890),
            .I(N__44883));
    InMux I__10434 (
            .O(N__44889),
            .I(N__44880));
    LocalMux I__10433 (
            .O(N__44886),
            .I(N__44877));
    Odrv4 I__10432 (
            .O(N__44883),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__10431 (
            .O(N__44880),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    Odrv4 I__10430 (
            .O(N__44877),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    InMux I__10429 (
            .O(N__44870),
            .I(N__44867));
    LocalMux I__10428 (
            .O(N__44867),
            .I(N__44862));
    InMux I__10427 (
            .O(N__44866),
            .I(N__44859));
    InMux I__10426 (
            .O(N__44865),
            .I(N__44856));
    Span4Mux_v I__10425 (
            .O(N__44862),
            .I(N__44851));
    LocalMux I__10424 (
            .O(N__44859),
            .I(N__44851));
    LocalMux I__10423 (
            .O(N__44856),
            .I(\delay_measurement_inst.elapsed_time_tr_4 ));
    Odrv4 I__10422 (
            .O(N__44851),
            .I(\delay_measurement_inst.elapsed_time_tr_4 ));
    InMux I__10421 (
            .O(N__44846),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ));
    CascadeMux I__10420 (
            .O(N__44843),
            .I(N__44839));
    CascadeMux I__10419 (
            .O(N__44842),
            .I(N__44836));
    InMux I__10418 (
            .O(N__44839),
            .I(N__44830));
    InMux I__10417 (
            .O(N__44836),
            .I(N__44830));
    InMux I__10416 (
            .O(N__44835),
            .I(N__44827));
    LocalMux I__10415 (
            .O(N__44830),
            .I(N__44824));
    LocalMux I__10414 (
            .O(N__44827),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    Odrv4 I__10413 (
            .O(N__44824),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    CascadeMux I__10412 (
            .O(N__44819),
            .I(N__44816));
    InMux I__10411 (
            .O(N__44816),
            .I(N__44813));
    LocalMux I__10410 (
            .O(N__44813),
            .I(N__44808));
    InMux I__10409 (
            .O(N__44812),
            .I(N__44803));
    InMux I__10408 (
            .O(N__44811),
            .I(N__44803));
    Span4Mux_h I__10407 (
            .O(N__44808),
            .I(N__44800));
    LocalMux I__10406 (
            .O(N__44803),
            .I(N__44797));
    Odrv4 I__10405 (
            .O(N__44800),
            .I(\delay_measurement_inst.elapsed_time_tr_5 ));
    Odrv12 I__10404 (
            .O(N__44797),
            .I(\delay_measurement_inst.elapsed_time_tr_5 ));
    InMux I__10403 (
            .O(N__44792),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__10402 (
            .O(N__44789),
            .I(N__44785));
    CascadeMux I__10401 (
            .O(N__44788),
            .I(N__44782));
    InMux I__10400 (
            .O(N__44785),
            .I(N__44776));
    InMux I__10399 (
            .O(N__44782),
            .I(N__44776));
    InMux I__10398 (
            .O(N__44781),
            .I(N__44773));
    LocalMux I__10397 (
            .O(N__44776),
            .I(N__44770));
    LocalMux I__10396 (
            .O(N__44773),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    Odrv4 I__10395 (
            .O(N__44770),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    InMux I__10394 (
            .O(N__44765),
            .I(N__44762));
    LocalMux I__10393 (
            .O(N__44762),
            .I(N__44757));
    InMux I__10392 (
            .O(N__44761),
            .I(N__44752));
    InMux I__10391 (
            .O(N__44760),
            .I(N__44752));
    Span4Mux_h I__10390 (
            .O(N__44757),
            .I(N__44749));
    LocalMux I__10389 (
            .O(N__44752),
            .I(N__44746));
    Odrv4 I__10388 (
            .O(N__44749),
            .I(\delay_measurement_inst.elapsed_time_tr_6 ));
    Odrv4 I__10387 (
            .O(N__44746),
            .I(\delay_measurement_inst.elapsed_time_tr_6 ));
    InMux I__10386 (
            .O(N__44741),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ));
    InMux I__10385 (
            .O(N__44738),
            .I(N__44732));
    InMux I__10384 (
            .O(N__44737),
            .I(N__44732));
    LocalMux I__10383 (
            .O(N__44732),
            .I(N__44728));
    InMux I__10382 (
            .O(N__44731),
            .I(N__44725));
    Span4Mux_h I__10381 (
            .O(N__44728),
            .I(N__44722));
    LocalMux I__10380 (
            .O(N__44725),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    Odrv4 I__10379 (
            .O(N__44722),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    InMux I__10378 (
            .O(N__44717),
            .I(N__44712));
    InMux I__10377 (
            .O(N__44716),
            .I(N__44709));
    InMux I__10376 (
            .O(N__44715),
            .I(N__44706));
    LocalMux I__10375 (
            .O(N__44712),
            .I(N__44701));
    LocalMux I__10374 (
            .O(N__44709),
            .I(N__44701));
    LocalMux I__10373 (
            .O(N__44706),
            .I(N__44698));
    Span4Mux_h I__10372 (
            .O(N__44701),
            .I(N__44695));
    Span4Mux_h I__10371 (
            .O(N__44698),
            .I(N__44692));
    Odrv4 I__10370 (
            .O(N__44695),
            .I(\delay_measurement_inst.elapsed_time_tr_7 ));
    Odrv4 I__10369 (
            .O(N__44692),
            .I(\delay_measurement_inst.elapsed_time_tr_7 ));
    InMux I__10368 (
            .O(N__44687),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ));
    InMux I__10367 (
            .O(N__44684),
            .I(N__44678));
    InMux I__10366 (
            .O(N__44683),
            .I(N__44678));
    LocalMux I__10365 (
            .O(N__44678),
            .I(N__44674));
    InMux I__10364 (
            .O(N__44677),
            .I(N__44671));
    Span4Mux_h I__10363 (
            .O(N__44674),
            .I(N__44668));
    LocalMux I__10362 (
            .O(N__44671),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    Odrv4 I__10361 (
            .O(N__44668),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    InMux I__10360 (
            .O(N__44663),
            .I(N__44659));
    InMux I__10359 (
            .O(N__44662),
            .I(N__44656));
    LocalMux I__10358 (
            .O(N__44659),
            .I(N__44652));
    LocalMux I__10357 (
            .O(N__44656),
            .I(N__44649));
    InMux I__10356 (
            .O(N__44655),
            .I(N__44646));
    Span4Mux_v I__10355 (
            .O(N__44652),
            .I(N__44639));
    Span4Mux_v I__10354 (
            .O(N__44649),
            .I(N__44639));
    LocalMux I__10353 (
            .O(N__44646),
            .I(N__44639));
    Odrv4 I__10352 (
            .O(N__44639),
            .I(\delay_measurement_inst.elapsed_time_tr_8 ));
    InMux I__10351 (
            .O(N__44636),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__10350 (
            .O(N__44633),
            .I(N__44630));
    InMux I__10349 (
            .O(N__44630),
            .I(N__44626));
    InMux I__10348 (
            .O(N__44629),
            .I(N__44622));
    LocalMux I__10347 (
            .O(N__44626),
            .I(N__44619));
    InMux I__10346 (
            .O(N__44625),
            .I(N__44616));
    LocalMux I__10345 (
            .O(N__44622),
            .I(N__44613));
    Span4Mux_h I__10344 (
            .O(N__44619),
            .I(N__44610));
    LocalMux I__10343 (
            .O(N__44616),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    Odrv4 I__10342 (
            .O(N__44613),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    Odrv4 I__10341 (
            .O(N__44610),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    InMux I__10340 (
            .O(N__44603),
            .I(N__44598));
    InMux I__10339 (
            .O(N__44602),
            .I(N__44595));
    CascadeMux I__10338 (
            .O(N__44601),
            .I(N__44591));
    LocalMux I__10337 (
            .O(N__44598),
            .I(N__44586));
    LocalMux I__10336 (
            .O(N__44595),
            .I(N__44586));
    InMux I__10335 (
            .O(N__44594),
            .I(N__44581));
    InMux I__10334 (
            .O(N__44591),
            .I(N__44581));
    Span12Mux_v I__10333 (
            .O(N__44586),
            .I(N__44576));
    LocalMux I__10332 (
            .O(N__44581),
            .I(N__44576));
    Odrv12 I__10331 (
            .O(N__44576),
            .I(\delay_measurement_inst.elapsed_time_tr_9 ));
    InMux I__10330 (
            .O(N__44573),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ));
    CascadeMux I__10329 (
            .O(N__44570),
            .I(N__44566));
    CascadeMux I__10328 (
            .O(N__44569),
            .I(N__44563));
    InMux I__10327 (
            .O(N__44566),
            .I(N__44558));
    InMux I__10326 (
            .O(N__44563),
            .I(N__44558));
    LocalMux I__10325 (
            .O(N__44558),
            .I(N__44554));
    InMux I__10324 (
            .O(N__44557),
            .I(N__44551));
    Span4Mux_v I__10323 (
            .O(N__44554),
            .I(N__44548));
    LocalMux I__10322 (
            .O(N__44551),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    Odrv4 I__10321 (
            .O(N__44548),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    InMux I__10320 (
            .O(N__44543),
            .I(N__44539));
    InMux I__10319 (
            .O(N__44542),
            .I(N__44536));
    LocalMux I__10318 (
            .O(N__44539),
            .I(N__44533));
    LocalMux I__10317 (
            .O(N__44536),
            .I(N__44530));
    Span4Mux_h I__10316 (
            .O(N__44533),
            .I(N__44527));
    Span4Mux_h I__10315 (
            .O(N__44530),
            .I(N__44524));
    Odrv4 I__10314 (
            .O(N__44527),
            .I(\delay_measurement_inst.elapsed_time_tr_10 ));
    Odrv4 I__10313 (
            .O(N__44524),
            .I(\delay_measurement_inst.elapsed_time_tr_10 ));
    InMux I__10312 (
            .O(N__44519),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ));
    InMux I__10311 (
            .O(N__44516),
            .I(N__44512));
    CascadeMux I__10310 (
            .O(N__44515),
            .I(N__44508));
    LocalMux I__10309 (
            .O(N__44512),
            .I(N__44505));
    InMux I__10308 (
            .O(N__44511),
            .I(N__44502));
    InMux I__10307 (
            .O(N__44508),
            .I(N__44499));
    Odrv4 I__10306 (
            .O(N__44505),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    LocalMux I__10305 (
            .O(N__44502),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    LocalMux I__10304 (
            .O(N__44499),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    InMux I__10303 (
            .O(N__44492),
            .I(N__44489));
    LocalMux I__10302 (
            .O(N__44489),
            .I(N__44485));
    InMux I__10301 (
            .O(N__44488),
            .I(N__44482));
    Span4Mux_v I__10300 (
            .O(N__44485),
            .I(N__44477));
    LocalMux I__10299 (
            .O(N__44482),
            .I(N__44477));
    Odrv4 I__10298 (
            .O(N__44477),
            .I(\delay_measurement_inst.elapsed_time_tr_11 ));
    InMux I__10297 (
            .O(N__44474),
            .I(bfn_18_14_0_));
    CascadeMux I__10296 (
            .O(N__44471),
            .I(N__44468));
    InMux I__10295 (
            .O(N__44468),
            .I(N__44465));
    LocalMux I__10294 (
            .O(N__44465),
            .I(N__44462));
    Span4Mux_v I__10293 (
            .O(N__44462),
            .I(N__44459));
    Span4Mux_h I__10292 (
            .O(N__44459),
            .I(N__44456));
    Odrv4 I__10291 (
            .O(N__44456),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_16 ));
    CEMux I__10290 (
            .O(N__44453),
            .I(N__44450));
    LocalMux I__10289 (
            .O(N__44450),
            .I(N__44446));
    CEMux I__10288 (
            .O(N__44449),
            .I(N__44441));
    Span4Mux_v I__10287 (
            .O(N__44446),
            .I(N__44438));
    CEMux I__10286 (
            .O(N__44445),
            .I(N__44435));
    CEMux I__10285 (
            .O(N__44444),
            .I(N__44432));
    LocalMux I__10284 (
            .O(N__44441),
            .I(N__44429));
    Span4Mux_h I__10283 (
            .O(N__44438),
            .I(N__44424));
    LocalMux I__10282 (
            .O(N__44435),
            .I(N__44424));
    LocalMux I__10281 (
            .O(N__44432),
            .I(N__44421));
    Span4Mux_v I__10280 (
            .O(N__44429),
            .I(N__44418));
    Span4Mux_v I__10279 (
            .O(N__44424),
            .I(N__44414));
    Span4Mux_h I__10278 (
            .O(N__44421),
            .I(N__44411));
    Span4Mux_h I__10277 (
            .O(N__44418),
            .I(N__44408));
    CEMux I__10276 (
            .O(N__44417),
            .I(N__44405));
    Span4Mux_v I__10275 (
            .O(N__44414),
            .I(N__44402));
    Span4Mux_v I__10274 (
            .O(N__44411),
            .I(N__44399));
    Span4Mux_v I__10273 (
            .O(N__44408),
            .I(N__44394));
    LocalMux I__10272 (
            .O(N__44405),
            .I(N__44394));
    Odrv4 I__10271 (
            .O(N__44402),
            .I(\phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv4 I__10270 (
            .O(N__44399),
            .I(\phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv4 I__10269 (
            .O(N__44394),
            .I(\phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa ));
    InMux I__10268 (
            .O(N__44387),
            .I(N__44379));
    InMux I__10267 (
            .O(N__44386),
            .I(N__44379));
    InMux I__10266 (
            .O(N__44385),
            .I(N__44376));
    InMux I__10265 (
            .O(N__44384),
            .I(N__44373));
    LocalMux I__10264 (
            .O(N__44379),
            .I(N__44370));
    LocalMux I__10263 (
            .O(N__44376),
            .I(N__44365));
    LocalMux I__10262 (
            .O(N__44373),
            .I(N__44365));
    Span4Mux_v I__10261 (
            .O(N__44370),
            .I(N__44362));
    Odrv12 I__10260 (
            .O(N__44365),
            .I(measured_delay_tr_16));
    Odrv4 I__10259 (
            .O(N__44362),
            .I(measured_delay_tr_16));
    CascadeMux I__10258 (
            .O(N__44357),
            .I(N__44354));
    InMux I__10257 (
            .O(N__44354),
            .I(N__44351));
    LocalMux I__10256 (
            .O(N__44351),
            .I(N__44348));
    Span4Mux_h I__10255 (
            .O(N__44348),
            .I(N__44345));
    Odrv4 I__10254 (
            .O(N__44345),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ));
    InMux I__10253 (
            .O(N__44342),
            .I(N__44338));
    InMux I__10252 (
            .O(N__44341),
            .I(N__44335));
    LocalMux I__10251 (
            .O(N__44338),
            .I(measured_delay_hc_29));
    LocalMux I__10250 (
            .O(N__44335),
            .I(measured_delay_hc_29));
    InMux I__10249 (
            .O(N__44330),
            .I(N__44326));
    InMux I__10248 (
            .O(N__44329),
            .I(N__44323));
    LocalMux I__10247 (
            .O(N__44326),
            .I(measured_delay_hc_28));
    LocalMux I__10246 (
            .O(N__44323),
            .I(measured_delay_hc_28));
    CascadeMux I__10245 (
            .O(N__44318),
            .I(N__44314));
    InMux I__10244 (
            .O(N__44317),
            .I(N__44311));
    InMux I__10243 (
            .O(N__44314),
            .I(N__44308));
    LocalMux I__10242 (
            .O(N__44311),
            .I(measured_delay_hc_30));
    LocalMux I__10241 (
            .O(N__44308),
            .I(measured_delay_hc_30));
    InMux I__10240 (
            .O(N__44303),
            .I(N__44299));
    InMux I__10239 (
            .O(N__44302),
            .I(N__44296));
    LocalMux I__10238 (
            .O(N__44299),
            .I(measured_delay_hc_27));
    LocalMux I__10237 (
            .O(N__44296),
            .I(measured_delay_hc_27));
    InMux I__10236 (
            .O(N__44291),
            .I(N__44288));
    LocalMux I__10235 (
            .O(N__44288),
            .I(N__44285));
    Odrv4 I__10234 (
            .O(N__44285),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_4 ));
    InMux I__10233 (
            .O(N__44282),
            .I(N__44278));
    InMux I__10232 (
            .O(N__44281),
            .I(N__44275));
    LocalMux I__10231 (
            .O(N__44278),
            .I(N__44270));
    LocalMux I__10230 (
            .O(N__44275),
            .I(N__44267));
    InMux I__10229 (
            .O(N__44274),
            .I(N__44264));
    CascadeMux I__10228 (
            .O(N__44273),
            .I(N__44261));
    Span4Mux_h I__10227 (
            .O(N__44270),
            .I(N__44257));
    Span4Mux_v I__10226 (
            .O(N__44267),
            .I(N__44254));
    LocalMux I__10225 (
            .O(N__44264),
            .I(N__44251));
    InMux I__10224 (
            .O(N__44261),
            .I(N__44248));
    CascadeMux I__10223 (
            .O(N__44260),
            .I(N__44245));
    Span4Mux_h I__10222 (
            .O(N__44257),
            .I(N__44236));
    Span4Mux_h I__10221 (
            .O(N__44254),
            .I(N__44236));
    Span4Mux_v I__10220 (
            .O(N__44251),
            .I(N__44236));
    LocalMux I__10219 (
            .O(N__44248),
            .I(N__44236));
    InMux I__10218 (
            .O(N__44245),
            .I(N__44233));
    Span4Mux_v I__10217 (
            .O(N__44236),
            .I(N__44230));
    LocalMux I__10216 (
            .O(N__44233),
            .I(measured_delay_hc_13));
    Odrv4 I__10215 (
            .O(N__44230),
            .I(measured_delay_hc_13));
    CascadeMux I__10214 (
            .O(N__44225),
            .I(N__44222));
    InMux I__10213 (
            .O(N__44222),
            .I(N__44219));
    LocalMux I__10212 (
            .O(N__44219),
            .I(N__44216));
    Span4Mux_v I__10211 (
            .O(N__44216),
            .I(N__44213));
    Span4Mux_v I__10210 (
            .O(N__44213),
            .I(N__44210));
    Odrv4 I__10209 (
            .O(N__44210),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_13 ));
    CascadeMux I__10208 (
            .O(N__44207),
            .I(N__44201));
    InMux I__10207 (
            .O(N__44206),
            .I(N__44189));
    InMux I__10206 (
            .O(N__44205),
            .I(N__44189));
    InMux I__10205 (
            .O(N__44204),
            .I(N__44189));
    InMux I__10204 (
            .O(N__44201),
            .I(N__44189));
    CascadeMux I__10203 (
            .O(N__44200),
            .I(N__44174));
    CascadeMux I__10202 (
            .O(N__44199),
            .I(N__44170));
    CascadeMux I__10201 (
            .O(N__44198),
            .I(N__44161));
    LocalMux I__10200 (
            .O(N__44189),
            .I(N__44158));
    CascadeMux I__10199 (
            .O(N__44188),
            .I(N__44151));
    CascadeMux I__10198 (
            .O(N__44187),
            .I(N__44148));
    CascadeMux I__10197 (
            .O(N__44186),
            .I(N__44145));
    CascadeMux I__10196 (
            .O(N__44185),
            .I(N__44141));
    InMux I__10195 (
            .O(N__44184),
            .I(N__44126));
    InMux I__10194 (
            .O(N__44183),
            .I(N__44126));
    InMux I__10193 (
            .O(N__44182),
            .I(N__44126));
    InMux I__10192 (
            .O(N__44181),
            .I(N__44126));
    InMux I__10191 (
            .O(N__44180),
            .I(N__44126));
    InMux I__10190 (
            .O(N__44179),
            .I(N__44126));
    InMux I__10189 (
            .O(N__44178),
            .I(N__44109));
    InMux I__10188 (
            .O(N__44177),
            .I(N__44109));
    InMux I__10187 (
            .O(N__44174),
            .I(N__44109));
    InMux I__10186 (
            .O(N__44173),
            .I(N__44109));
    InMux I__10185 (
            .O(N__44170),
            .I(N__44109));
    InMux I__10184 (
            .O(N__44169),
            .I(N__44109));
    InMux I__10183 (
            .O(N__44168),
            .I(N__44109));
    InMux I__10182 (
            .O(N__44167),
            .I(N__44109));
    InMux I__10181 (
            .O(N__44166),
            .I(N__44100));
    InMux I__10180 (
            .O(N__44165),
            .I(N__44100));
    InMux I__10179 (
            .O(N__44164),
            .I(N__44100));
    InMux I__10178 (
            .O(N__44161),
            .I(N__44100));
    Span4Mux_v I__10177 (
            .O(N__44158),
            .I(N__44097));
    InMux I__10176 (
            .O(N__44157),
            .I(N__44094));
    InMux I__10175 (
            .O(N__44156),
            .I(N__44091));
    CascadeMux I__10174 (
            .O(N__44155),
            .I(N__44088));
    InMux I__10173 (
            .O(N__44154),
            .I(N__44081));
    InMux I__10172 (
            .O(N__44151),
            .I(N__44066));
    InMux I__10171 (
            .O(N__44148),
            .I(N__44066));
    InMux I__10170 (
            .O(N__44145),
            .I(N__44066));
    InMux I__10169 (
            .O(N__44144),
            .I(N__44066));
    InMux I__10168 (
            .O(N__44141),
            .I(N__44066));
    InMux I__10167 (
            .O(N__44140),
            .I(N__44066));
    InMux I__10166 (
            .O(N__44139),
            .I(N__44066));
    LocalMux I__10165 (
            .O(N__44126),
            .I(N__44063));
    LocalMux I__10164 (
            .O(N__44109),
            .I(N__44055));
    LocalMux I__10163 (
            .O(N__44100),
            .I(N__44055));
    Span4Mux_h I__10162 (
            .O(N__44097),
            .I(N__44052));
    LocalMux I__10161 (
            .O(N__44094),
            .I(N__44049));
    LocalMux I__10160 (
            .O(N__44091),
            .I(N__44046));
    InMux I__10159 (
            .O(N__44088),
            .I(N__44039));
    InMux I__10158 (
            .O(N__44087),
            .I(N__44039));
    InMux I__10157 (
            .O(N__44086),
            .I(N__44039));
    InMux I__10156 (
            .O(N__44085),
            .I(N__44034));
    InMux I__10155 (
            .O(N__44084),
            .I(N__44034));
    LocalMux I__10154 (
            .O(N__44081),
            .I(N__44031));
    LocalMux I__10153 (
            .O(N__44066),
            .I(N__44028));
    Span4Mux_h I__10152 (
            .O(N__44063),
            .I(N__44025));
    InMux I__10151 (
            .O(N__44062),
            .I(N__44018));
    InMux I__10150 (
            .O(N__44061),
            .I(N__44018));
    InMux I__10149 (
            .O(N__44060),
            .I(N__44018));
    Span4Mux_v I__10148 (
            .O(N__44055),
            .I(N__44014));
    Span4Mux_h I__10147 (
            .O(N__44052),
            .I(N__44009));
    Span4Mux_h I__10146 (
            .O(N__44049),
            .I(N__44009));
    Span4Mux_h I__10145 (
            .O(N__44046),
            .I(N__44006));
    LocalMux I__10144 (
            .O(N__44039),
            .I(N__44001));
    LocalMux I__10143 (
            .O(N__44034),
            .I(N__44001));
    Span4Mux_h I__10142 (
            .O(N__44031),
            .I(N__43998));
    Span4Mux_v I__10141 (
            .O(N__44028),
            .I(N__43995));
    Span4Mux_v I__10140 (
            .O(N__44025),
            .I(N__43990));
    LocalMux I__10139 (
            .O(N__44018),
            .I(N__43990));
    InMux I__10138 (
            .O(N__44017),
            .I(N__43987));
    Span4Mux_v I__10137 (
            .O(N__44014),
            .I(N__43984));
    Span4Mux_v I__10136 (
            .O(N__44009),
            .I(N__43979));
    Span4Mux_v I__10135 (
            .O(N__44006),
            .I(N__43979));
    Span12Mux_h I__10134 (
            .O(N__44001),
            .I(N__43976));
    Span4Mux_h I__10133 (
            .O(N__43998),
            .I(N__43969));
    Span4Mux_h I__10132 (
            .O(N__43995),
            .I(N__43969));
    Span4Mux_v I__10131 (
            .O(N__43990),
            .I(N__43969));
    LocalMux I__10130 (
            .O(N__43987),
            .I(measured_delay_hc_31));
    Odrv4 I__10129 (
            .O(N__43984),
            .I(measured_delay_hc_31));
    Odrv4 I__10128 (
            .O(N__43979),
            .I(measured_delay_hc_31));
    Odrv12 I__10127 (
            .O(N__43976),
            .I(measured_delay_hc_31));
    Odrv4 I__10126 (
            .O(N__43969),
            .I(measured_delay_hc_31));
    CascadeMux I__10125 (
            .O(N__43958),
            .I(N__43951));
    InMux I__10124 (
            .O(N__43957),
            .I(N__43948));
    InMux I__10123 (
            .O(N__43956),
            .I(N__43945));
    InMux I__10122 (
            .O(N__43955),
            .I(N__43942));
    InMux I__10121 (
            .O(N__43954),
            .I(N__43939));
    InMux I__10120 (
            .O(N__43951),
            .I(N__43936));
    LocalMux I__10119 (
            .O(N__43948),
            .I(N__43933));
    LocalMux I__10118 (
            .O(N__43945),
            .I(N__43930));
    LocalMux I__10117 (
            .O(N__43942),
            .I(N__43927));
    LocalMux I__10116 (
            .O(N__43939),
            .I(N__43924));
    LocalMux I__10115 (
            .O(N__43936),
            .I(measured_delay_hc_5));
    Odrv12 I__10114 (
            .O(N__43933),
            .I(measured_delay_hc_5));
    Odrv12 I__10113 (
            .O(N__43930),
            .I(measured_delay_hc_5));
    Odrv4 I__10112 (
            .O(N__43927),
            .I(measured_delay_hc_5));
    Odrv4 I__10111 (
            .O(N__43924),
            .I(measured_delay_hc_5));
    InMux I__10110 (
            .O(N__43913),
            .I(N__43901));
    InMux I__10109 (
            .O(N__43912),
            .I(N__43901));
    InMux I__10108 (
            .O(N__43911),
            .I(N__43901));
    InMux I__10107 (
            .O(N__43910),
            .I(N__43901));
    LocalMux I__10106 (
            .O(N__43901),
            .I(N__43889));
    InMux I__10105 (
            .O(N__43900),
            .I(N__43880));
    InMux I__10104 (
            .O(N__43899),
            .I(N__43880));
    InMux I__10103 (
            .O(N__43898),
            .I(N__43880));
    InMux I__10102 (
            .O(N__43897),
            .I(N__43875));
    InMux I__10101 (
            .O(N__43896),
            .I(N__43864));
    InMux I__10100 (
            .O(N__43895),
            .I(N__43864));
    InMux I__10099 (
            .O(N__43894),
            .I(N__43864));
    InMux I__10098 (
            .O(N__43893),
            .I(N__43864));
    InMux I__10097 (
            .O(N__43892),
            .I(N__43864));
    Span4Mux_h I__10096 (
            .O(N__43889),
            .I(N__43841));
    InMux I__10095 (
            .O(N__43888),
            .I(N__43836));
    InMux I__10094 (
            .O(N__43887),
            .I(N__43836));
    LocalMux I__10093 (
            .O(N__43880),
            .I(N__43833));
    InMux I__10092 (
            .O(N__43879),
            .I(N__43828));
    InMux I__10091 (
            .O(N__43878),
            .I(N__43828));
    LocalMux I__10090 (
            .O(N__43875),
            .I(N__43824));
    LocalMux I__10089 (
            .O(N__43864),
            .I(N__43821));
    InMux I__10088 (
            .O(N__43863),
            .I(N__43804));
    InMux I__10087 (
            .O(N__43862),
            .I(N__43804));
    InMux I__10086 (
            .O(N__43861),
            .I(N__43804));
    InMux I__10085 (
            .O(N__43860),
            .I(N__43804));
    InMux I__10084 (
            .O(N__43859),
            .I(N__43804));
    InMux I__10083 (
            .O(N__43858),
            .I(N__43804));
    InMux I__10082 (
            .O(N__43857),
            .I(N__43804));
    InMux I__10081 (
            .O(N__43856),
            .I(N__43804));
    InMux I__10080 (
            .O(N__43855),
            .I(N__43795));
    InMux I__10079 (
            .O(N__43854),
            .I(N__43795));
    InMux I__10078 (
            .O(N__43853),
            .I(N__43795));
    InMux I__10077 (
            .O(N__43852),
            .I(N__43795));
    InMux I__10076 (
            .O(N__43851),
            .I(N__43792));
    InMux I__10075 (
            .O(N__43850),
            .I(N__43777));
    InMux I__10074 (
            .O(N__43849),
            .I(N__43777));
    InMux I__10073 (
            .O(N__43848),
            .I(N__43777));
    InMux I__10072 (
            .O(N__43847),
            .I(N__43777));
    InMux I__10071 (
            .O(N__43846),
            .I(N__43777));
    InMux I__10070 (
            .O(N__43845),
            .I(N__43777));
    InMux I__10069 (
            .O(N__43844),
            .I(N__43777));
    Span4Mux_h I__10068 (
            .O(N__43841),
            .I(N__43772));
    LocalMux I__10067 (
            .O(N__43836),
            .I(N__43772));
    Sp12to4 I__10066 (
            .O(N__43833),
            .I(N__43767));
    LocalMux I__10065 (
            .O(N__43828),
            .I(N__43767));
    InMux I__10064 (
            .O(N__43827),
            .I(N__43764));
    Span4Mux_h I__10063 (
            .O(N__43824),
            .I(N__43761));
    Span12Mux_s11_h I__10062 (
            .O(N__43821),
            .I(N__43754));
    LocalMux I__10061 (
            .O(N__43804),
            .I(N__43754));
    LocalMux I__10060 (
            .O(N__43795),
            .I(N__43754));
    LocalMux I__10059 (
            .O(N__43792),
            .I(N__43749));
    LocalMux I__10058 (
            .O(N__43777),
            .I(N__43749));
    Span4Mux_h I__10057 (
            .O(N__43772),
            .I(N__43746));
    Span12Mux_v I__10056 (
            .O(N__43767),
            .I(N__43741));
    LocalMux I__10055 (
            .O(N__43764),
            .I(N__43741));
    Odrv4 I__10054 (
            .O(N__43761),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt31_0 ));
    Odrv12 I__10053 (
            .O(N__43754),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt31_0 ));
    Odrv12 I__10052 (
            .O(N__43749),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt31_0 ));
    Odrv4 I__10051 (
            .O(N__43746),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt31_0 ));
    Odrv12 I__10050 (
            .O(N__43741),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt31_0 ));
    CascadeMux I__10049 (
            .O(N__43730),
            .I(N__43727));
    InMux I__10048 (
            .O(N__43727),
            .I(N__43724));
    LocalMux I__10047 (
            .O(N__43724),
            .I(N__43721));
    Span4Mux_v I__10046 (
            .O(N__43721),
            .I(N__43718));
    Span4Mux_h I__10045 (
            .O(N__43718),
            .I(N__43715));
    Odrv4 I__10044 (
            .O(N__43715),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_5 ));
    CEMux I__10043 (
            .O(N__43712),
            .I(N__43708));
    CEMux I__10042 (
            .O(N__43711),
            .I(N__43704));
    LocalMux I__10041 (
            .O(N__43708),
            .I(N__43701));
    CEMux I__10040 (
            .O(N__43707),
            .I(N__43697));
    LocalMux I__10039 (
            .O(N__43704),
            .I(N__43694));
    Span4Mux_v I__10038 (
            .O(N__43701),
            .I(N__43691));
    CEMux I__10037 (
            .O(N__43700),
            .I(N__43688));
    LocalMux I__10036 (
            .O(N__43697),
            .I(N__43684));
    Span4Mux_v I__10035 (
            .O(N__43694),
            .I(N__43681));
    Span4Mux_h I__10034 (
            .O(N__43691),
            .I(N__43676));
    LocalMux I__10033 (
            .O(N__43688),
            .I(N__43676));
    CEMux I__10032 (
            .O(N__43687),
            .I(N__43673));
    Span4Mux_h I__10031 (
            .O(N__43684),
            .I(N__43670));
    Span4Mux_h I__10030 (
            .O(N__43681),
            .I(N__43667));
    Span4Mux_v I__10029 (
            .O(N__43676),
            .I(N__43662));
    LocalMux I__10028 (
            .O(N__43673),
            .I(N__43662));
    Span4Mux_h I__10027 (
            .O(N__43670),
            .I(N__43659));
    Span4Mux_v I__10026 (
            .O(N__43667),
            .I(N__43654));
    Span4Mux_h I__10025 (
            .O(N__43662),
            .I(N__43654));
    Odrv4 I__10024 (
            .O(N__43659),
            .I(\phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa ));
    Odrv4 I__10023 (
            .O(N__43654),
            .I(\phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa ));
    CascadeMux I__10022 (
            .O(N__43649),
            .I(N__43642));
    CascadeMux I__10021 (
            .O(N__43648),
            .I(N__43639));
    InMux I__10020 (
            .O(N__43647),
            .I(N__43635));
    InMux I__10019 (
            .O(N__43646),
            .I(N__43632));
    InMux I__10018 (
            .O(N__43645),
            .I(N__43623));
    InMux I__10017 (
            .O(N__43642),
            .I(N__43623));
    InMux I__10016 (
            .O(N__43639),
            .I(N__43623));
    InMux I__10015 (
            .O(N__43638),
            .I(N__43623));
    LocalMux I__10014 (
            .O(N__43635),
            .I(N__43620));
    LocalMux I__10013 (
            .O(N__43632),
            .I(N__43612));
    LocalMux I__10012 (
            .O(N__43623),
            .I(N__43612));
    Span4Mux_h I__10011 (
            .O(N__43620),
            .I(N__43612));
    InMux I__10010 (
            .O(N__43619),
            .I(N__43609));
    Odrv4 I__10009 (
            .O(N__43612),
            .I(\delay_measurement_inst.N_410 ));
    LocalMux I__10008 (
            .O(N__43609),
            .I(\delay_measurement_inst.N_410 ));
    CascadeMux I__10007 (
            .O(N__43604),
            .I(N__43598));
    CascadeMux I__10006 (
            .O(N__43603),
            .I(N__43595));
    CascadeMux I__10005 (
            .O(N__43602),
            .I(N__43588));
    CascadeMux I__10004 (
            .O(N__43601),
            .I(N__43585));
    InMux I__10003 (
            .O(N__43598),
            .I(N__43582));
    InMux I__10002 (
            .O(N__43595),
            .I(N__43577));
    InMux I__10001 (
            .O(N__43594),
            .I(N__43577));
    InMux I__10000 (
            .O(N__43593),
            .I(N__43566));
    InMux I__9999 (
            .O(N__43592),
            .I(N__43566));
    InMux I__9998 (
            .O(N__43591),
            .I(N__43566));
    InMux I__9997 (
            .O(N__43588),
            .I(N__43566));
    InMux I__9996 (
            .O(N__43585),
            .I(N__43566));
    LocalMux I__9995 (
            .O(N__43582),
            .I(N__43563));
    LocalMux I__9994 (
            .O(N__43577),
            .I(N__43560));
    LocalMux I__9993 (
            .O(N__43566),
            .I(N__43553));
    Span4Mux_h I__9992 (
            .O(N__43563),
            .I(N__43553));
    Span4Mux_h I__9991 (
            .O(N__43560),
            .I(N__43553));
    Odrv4 I__9990 (
            .O(N__43553),
            .I(\delay_measurement_inst.N_358 ));
    InMux I__9989 (
            .O(N__43550),
            .I(N__43547));
    LocalMux I__9988 (
            .O(N__43547),
            .I(N__43538));
    InMux I__9987 (
            .O(N__43546),
            .I(N__43527));
    InMux I__9986 (
            .O(N__43545),
            .I(N__43527));
    InMux I__9985 (
            .O(N__43544),
            .I(N__43527));
    InMux I__9984 (
            .O(N__43543),
            .I(N__43527));
    InMux I__9983 (
            .O(N__43542),
            .I(N__43527));
    InMux I__9982 (
            .O(N__43541),
            .I(N__43524));
    Span4Mux_v I__9981 (
            .O(N__43538),
            .I(N__43520));
    LocalMux I__9980 (
            .O(N__43527),
            .I(N__43517));
    LocalMux I__9979 (
            .O(N__43524),
            .I(N__43514));
    InMux I__9978 (
            .O(N__43523),
            .I(N__43511));
    Odrv4 I__9977 (
            .O(N__43520),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15 ));
    Odrv12 I__9976 (
            .O(N__43517),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15 ));
    Odrv4 I__9975 (
            .O(N__43514),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15 ));
    LocalMux I__9974 (
            .O(N__43511),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15 ));
    InMux I__9973 (
            .O(N__43502),
            .I(N__43498));
    CascadeMux I__9972 (
            .O(N__43501),
            .I(N__43494));
    LocalMux I__9971 (
            .O(N__43498),
            .I(N__43491));
    InMux I__9970 (
            .O(N__43497),
            .I(N__43488));
    InMux I__9969 (
            .O(N__43494),
            .I(N__43485));
    Span4Mux_v I__9968 (
            .O(N__43491),
            .I(N__43480));
    LocalMux I__9967 (
            .O(N__43488),
            .I(N__43480));
    LocalMux I__9966 (
            .O(N__43485),
            .I(N__43477));
    Span4Mux_v I__9965 (
            .O(N__43480),
            .I(N__43474));
    Span12Mux_h I__9964 (
            .O(N__43477),
            .I(N__43471));
    Span4Mux_v I__9963 (
            .O(N__43474),
            .I(N__43468));
    Odrv12 I__9962 (
            .O(N__43471),
            .I(measured_delay_tr_4));
    Odrv4 I__9961 (
            .O(N__43468),
            .I(measured_delay_tr_4));
    CEMux I__9960 (
            .O(N__43463),
            .I(N__43458));
    CEMux I__9959 (
            .O(N__43462),
            .I(N__43455));
    CEMux I__9958 (
            .O(N__43461),
            .I(N__43452));
    LocalMux I__9957 (
            .O(N__43458),
            .I(N__43448));
    LocalMux I__9956 (
            .O(N__43455),
            .I(N__43445));
    LocalMux I__9955 (
            .O(N__43452),
            .I(N__43442));
    CEMux I__9954 (
            .O(N__43451),
            .I(N__43439));
    Span4Mux_v I__9953 (
            .O(N__43448),
            .I(N__43434));
    Span4Mux_h I__9952 (
            .O(N__43445),
            .I(N__43434));
    Span4Mux_v I__9951 (
            .O(N__43442),
            .I(N__43429));
    LocalMux I__9950 (
            .O(N__43439),
            .I(N__43429));
    Odrv4 I__9949 (
            .O(N__43434),
            .I(\delay_measurement_inst.N_265_i_0 ));
    Odrv4 I__9948 (
            .O(N__43429),
            .I(\delay_measurement_inst.N_265_i_0 ));
    InMux I__9947 (
            .O(N__43424),
            .I(N__43420));
    InMux I__9946 (
            .O(N__43423),
            .I(N__43416));
    LocalMux I__9945 (
            .O(N__43420),
            .I(N__43413));
    InMux I__9944 (
            .O(N__43419),
            .I(N__43410));
    LocalMux I__9943 (
            .O(N__43416),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    Odrv4 I__9942 (
            .O(N__43413),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__9941 (
            .O(N__43410),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    CascadeMux I__9940 (
            .O(N__43403),
            .I(N__43398));
    CascadeMux I__9939 (
            .O(N__43402),
            .I(N__43395));
    InMux I__9938 (
            .O(N__43401),
            .I(N__43392));
    InMux I__9937 (
            .O(N__43398),
            .I(N__43389));
    InMux I__9936 (
            .O(N__43395),
            .I(N__43386));
    LocalMux I__9935 (
            .O(N__43392),
            .I(N__43383));
    LocalMux I__9934 (
            .O(N__43389),
            .I(N__43380));
    LocalMux I__9933 (
            .O(N__43386),
            .I(N__43377));
    Span4Mux_v I__9932 (
            .O(N__43383),
            .I(N__43370));
    Span4Mux_h I__9931 (
            .O(N__43380),
            .I(N__43370));
    Span4Mux_v I__9930 (
            .O(N__43377),
            .I(N__43370));
    Odrv4 I__9929 (
            .O(N__43370),
            .I(\delay_measurement_inst.elapsed_time_tr_3 ));
    InMux I__9928 (
            .O(N__43367),
            .I(N__43363));
    InMux I__9927 (
            .O(N__43366),
            .I(N__43359));
    LocalMux I__9926 (
            .O(N__43363),
            .I(N__43356));
    InMux I__9925 (
            .O(N__43362),
            .I(N__43353));
    LocalMux I__9924 (
            .O(N__43359),
            .I(\phase_controller_inst1.stoper_tr.time_passed11 ));
    Odrv4 I__9923 (
            .O(N__43356),
            .I(\phase_controller_inst1.stoper_tr.time_passed11 ));
    LocalMux I__9922 (
            .O(N__43353),
            .I(\phase_controller_inst1.stoper_tr.time_passed11 ));
    InMux I__9921 (
            .O(N__43346),
            .I(N__43338));
    InMux I__9920 (
            .O(N__43345),
            .I(N__43338));
    CascadeMux I__9919 (
            .O(N__43344),
            .I(N__43335));
    InMux I__9918 (
            .O(N__43343),
            .I(N__43330));
    LocalMux I__9917 (
            .O(N__43338),
            .I(N__43327));
    InMux I__9916 (
            .O(N__43335),
            .I(N__43320));
    InMux I__9915 (
            .O(N__43334),
            .I(N__43320));
    InMux I__9914 (
            .O(N__43333),
            .I(N__43320));
    LocalMux I__9913 (
            .O(N__43330),
            .I(N__43317));
    Span4Mux_h I__9912 (
            .O(N__43327),
            .I(N__43314));
    LocalMux I__9911 (
            .O(N__43320),
            .I(N__43311));
    Odrv4 I__9910 (
            .O(N__43317),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__9909 (
            .O(N__43314),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv12 I__9908 (
            .O(N__43311),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    CascadeMux I__9907 (
            .O(N__43304),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ));
    CascadeMux I__9906 (
            .O(N__43301),
            .I(\phase_controller_inst1.stoper_tr.time_passed11_cascade_ ));
    InMux I__9905 (
            .O(N__43298),
            .I(N__43293));
    InMux I__9904 (
            .O(N__43297),
            .I(N__43290));
    CascadeMux I__9903 (
            .O(N__43296),
            .I(N__43286));
    LocalMux I__9902 (
            .O(N__43293),
            .I(N__43283));
    LocalMux I__9901 (
            .O(N__43290),
            .I(N__43280));
    InMux I__9900 (
            .O(N__43289),
            .I(N__43275));
    InMux I__9899 (
            .O(N__43286),
            .I(N__43275));
    Span4Mux_h I__9898 (
            .O(N__43283),
            .I(N__43272));
    Span4Mux_v I__9897 (
            .O(N__43280),
            .I(N__43267));
    LocalMux I__9896 (
            .O(N__43275),
            .I(N__43267));
    Span4Mux_v I__9895 (
            .O(N__43272),
            .I(N__43264));
    Span4Mux_v I__9894 (
            .O(N__43267),
            .I(N__43261));
    Odrv4 I__9893 (
            .O(N__43264),
            .I(measured_delay_tr_17));
    Odrv4 I__9892 (
            .O(N__43261),
            .I(measured_delay_tr_17));
    InMux I__9891 (
            .O(N__43256),
            .I(N__43246));
    InMux I__9890 (
            .O(N__43255),
            .I(N__43246));
    InMux I__9889 (
            .O(N__43254),
            .I(N__43246));
    InMux I__9888 (
            .O(N__43253),
            .I(N__43243));
    LocalMux I__9887 (
            .O(N__43246),
            .I(N__43236));
    LocalMux I__9886 (
            .O(N__43243),
            .I(N__43233));
    InMux I__9885 (
            .O(N__43242),
            .I(N__43230));
    InMux I__9884 (
            .O(N__43241),
            .I(N__43225));
    InMux I__9883 (
            .O(N__43240),
            .I(N__43225));
    InMux I__9882 (
            .O(N__43239),
            .I(N__43222));
    Odrv4 I__9881 (
            .O(N__43236),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20 ));
    Odrv4 I__9880 (
            .O(N__43233),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20 ));
    LocalMux I__9879 (
            .O(N__43230),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20 ));
    LocalMux I__9878 (
            .O(N__43225),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20 ));
    LocalMux I__9877 (
            .O(N__43222),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20 ));
    InMux I__9876 (
            .O(N__43211),
            .I(N__43207));
    InMux I__9875 (
            .O(N__43210),
            .I(N__43202));
    LocalMux I__9874 (
            .O(N__43207),
            .I(N__43199));
    InMux I__9873 (
            .O(N__43206),
            .I(N__43194));
    InMux I__9872 (
            .O(N__43205),
            .I(N__43194));
    LocalMux I__9871 (
            .O(N__43202),
            .I(N__43191));
    Span4Mux_v I__9870 (
            .O(N__43199),
            .I(N__43186));
    LocalMux I__9869 (
            .O(N__43194),
            .I(N__43186));
    Span4Mux_v I__9868 (
            .O(N__43191),
            .I(N__43183));
    Span4Mux_v I__9867 (
            .O(N__43186),
            .I(N__43180));
    Odrv4 I__9866 (
            .O(N__43183),
            .I(measured_delay_tr_18));
    Odrv4 I__9865 (
            .O(N__43180),
            .I(measured_delay_tr_18));
    InMux I__9864 (
            .O(N__43175),
            .I(N__43172));
    LocalMux I__9863 (
            .O(N__43172),
            .I(N__43169));
    Span4Mux_v I__9862 (
            .O(N__43169),
            .I(N__43166));
    Span4Mux_h I__9861 (
            .O(N__43166),
            .I(N__43163));
    Odrv4 I__9860 (
            .O(N__43163),
            .I(\phase_controller_inst1.N_83 ));
    InMux I__9859 (
            .O(N__43160),
            .I(N__43157));
    LocalMux I__9858 (
            .O(N__43157),
            .I(N__43154));
    Span12Mux_h I__9857 (
            .O(N__43154),
            .I(N__43147));
    InMux I__9856 (
            .O(N__43153),
            .I(N__43144));
    InMux I__9855 (
            .O(N__43152),
            .I(N__43141));
    InMux I__9854 (
            .O(N__43151),
            .I(N__43136));
    InMux I__9853 (
            .O(N__43150),
            .I(N__43136));
    Odrv12 I__9852 (
            .O(N__43147),
            .I(\phase_controller_inst1.stateZ0Z_4 ));
    LocalMux I__9851 (
            .O(N__43144),
            .I(\phase_controller_inst1.stateZ0Z_4 ));
    LocalMux I__9850 (
            .O(N__43141),
            .I(\phase_controller_inst1.stateZ0Z_4 ));
    LocalMux I__9849 (
            .O(N__43136),
            .I(\phase_controller_inst1.stateZ0Z_4 ));
    CascadeMux I__9848 (
            .O(N__43127),
            .I(\phase_controller_inst1.N_83_cascade_ ));
    InMux I__9847 (
            .O(N__43124),
            .I(N__43121));
    LocalMux I__9846 (
            .O(N__43121),
            .I(N__43118));
    Span4Mux_v I__9845 (
            .O(N__43118),
            .I(N__43114));
    InMux I__9844 (
            .O(N__43117),
            .I(N__43111));
    Span4Mux_h I__9843 (
            .O(N__43114),
            .I(N__43106));
    LocalMux I__9842 (
            .O(N__43111),
            .I(N__43106));
    Odrv4 I__9841 (
            .O(N__43106),
            .I(\phase_controller_inst1.T01_0_sqmuxa ));
    CascadeMux I__9840 (
            .O(N__43103),
            .I(\phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa_cascade_ ));
    InMux I__9839 (
            .O(N__43100),
            .I(N__43097));
    LocalMux I__9838 (
            .O(N__43097),
            .I(N__43093));
    InMux I__9837 (
            .O(N__43096),
            .I(N__43090));
    Span4Mux_v I__9836 (
            .O(N__43093),
            .I(N__43087));
    LocalMux I__9835 (
            .O(N__43090),
            .I(N__43084));
    Span4Mux_v I__9834 (
            .O(N__43087),
            .I(N__43081));
    Span4Mux_v I__9833 (
            .O(N__43084),
            .I(N__43078));
    Span4Mux_v I__9832 (
            .O(N__43081),
            .I(N__43071));
    Span4Mux_h I__9831 (
            .O(N__43078),
            .I(N__43071));
    InMux I__9830 (
            .O(N__43077),
            .I(N__43068));
    InMux I__9829 (
            .O(N__43076),
            .I(N__43065));
    Span4Mux_v I__9828 (
            .O(N__43071),
            .I(N__43060));
    LocalMux I__9827 (
            .O(N__43068),
            .I(N__43060));
    LocalMux I__9826 (
            .O(N__43065),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv4 I__9825 (
            .O(N__43060),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    CascadeMux I__9824 (
            .O(N__43055),
            .I(N__43051));
    InMux I__9823 (
            .O(N__43054),
            .I(N__43043));
    InMux I__9822 (
            .O(N__43051),
            .I(N__43043));
    InMux I__9821 (
            .O(N__43050),
            .I(N__43043));
    LocalMux I__9820 (
            .O(N__43043),
            .I(\phase_controller_inst1.tr_time_passed ));
    InMux I__9819 (
            .O(N__43040),
            .I(N__43037));
    LocalMux I__9818 (
            .O(N__43037),
            .I(N__43034));
    Span4Mux_h I__9817 (
            .O(N__43034),
            .I(N__43030));
    InMux I__9816 (
            .O(N__43033),
            .I(N__43027));
    Span4Mux_h I__9815 (
            .O(N__43030),
            .I(N__43024));
    LocalMux I__9814 (
            .O(N__43027),
            .I(N__43020));
    Span4Mux_v I__9813 (
            .O(N__43024),
            .I(N__43017));
    InMux I__9812 (
            .O(N__43023),
            .I(N__43014));
    Span4Mux_h I__9811 (
            .O(N__43020),
            .I(N__43011));
    Odrv4 I__9810 (
            .O(N__43017),
            .I(il_min_comp1_D2));
    LocalMux I__9809 (
            .O(N__43014),
            .I(il_min_comp1_D2));
    Odrv4 I__9808 (
            .O(N__43011),
            .I(il_min_comp1_D2));
    InMux I__9807 (
            .O(N__43004),
            .I(N__42998));
    InMux I__9806 (
            .O(N__43003),
            .I(N__42998));
    LocalMux I__9805 (
            .O(N__42998),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    InMux I__9804 (
            .O(N__42995),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ));
    InMux I__9803 (
            .O(N__42992),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ));
    InMux I__9802 (
            .O(N__42989),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ));
    InMux I__9801 (
            .O(N__42986),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ));
    InMux I__9800 (
            .O(N__42983),
            .I(N__42971));
    InMux I__9799 (
            .O(N__42982),
            .I(N__42971));
    InMux I__9798 (
            .O(N__42981),
            .I(N__42971));
    InMux I__9797 (
            .O(N__42980),
            .I(N__42971));
    LocalMux I__9796 (
            .O(N__42971),
            .I(N__42942));
    InMux I__9795 (
            .O(N__42970),
            .I(N__42937));
    InMux I__9794 (
            .O(N__42969),
            .I(N__42937));
    InMux I__9793 (
            .O(N__42968),
            .I(N__42928));
    InMux I__9792 (
            .O(N__42967),
            .I(N__42928));
    InMux I__9791 (
            .O(N__42966),
            .I(N__42928));
    InMux I__9790 (
            .O(N__42965),
            .I(N__42928));
    InMux I__9789 (
            .O(N__42964),
            .I(N__42919));
    InMux I__9788 (
            .O(N__42963),
            .I(N__42919));
    InMux I__9787 (
            .O(N__42962),
            .I(N__42919));
    InMux I__9786 (
            .O(N__42961),
            .I(N__42919));
    InMux I__9785 (
            .O(N__42960),
            .I(N__42910));
    InMux I__9784 (
            .O(N__42959),
            .I(N__42910));
    InMux I__9783 (
            .O(N__42958),
            .I(N__42910));
    InMux I__9782 (
            .O(N__42957),
            .I(N__42910));
    InMux I__9781 (
            .O(N__42956),
            .I(N__42901));
    InMux I__9780 (
            .O(N__42955),
            .I(N__42901));
    InMux I__9779 (
            .O(N__42954),
            .I(N__42901));
    InMux I__9778 (
            .O(N__42953),
            .I(N__42901));
    InMux I__9777 (
            .O(N__42952),
            .I(N__42892));
    InMux I__9776 (
            .O(N__42951),
            .I(N__42892));
    InMux I__9775 (
            .O(N__42950),
            .I(N__42892));
    InMux I__9774 (
            .O(N__42949),
            .I(N__42892));
    InMux I__9773 (
            .O(N__42948),
            .I(N__42883));
    InMux I__9772 (
            .O(N__42947),
            .I(N__42883));
    InMux I__9771 (
            .O(N__42946),
            .I(N__42883));
    InMux I__9770 (
            .O(N__42945),
            .I(N__42883));
    Span4Mux_h I__9769 (
            .O(N__42942),
            .I(N__42878));
    LocalMux I__9768 (
            .O(N__42937),
            .I(N__42878));
    LocalMux I__9767 (
            .O(N__42928),
            .I(N__42873));
    LocalMux I__9766 (
            .O(N__42919),
            .I(N__42873));
    LocalMux I__9765 (
            .O(N__42910),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    LocalMux I__9764 (
            .O(N__42901),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    LocalMux I__9763 (
            .O(N__42892),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    LocalMux I__9762 (
            .O(N__42883),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    Odrv4 I__9761 (
            .O(N__42878),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    Odrv4 I__9760 (
            .O(N__42873),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    InMux I__9759 (
            .O(N__42860),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ));
    CEMux I__9758 (
            .O(N__42857),
            .I(N__42853));
    CEMux I__9757 (
            .O(N__42856),
            .I(N__42850));
    LocalMux I__9756 (
            .O(N__42853),
            .I(N__42846));
    LocalMux I__9755 (
            .O(N__42850),
            .I(N__42843));
    CEMux I__9754 (
            .O(N__42849),
            .I(N__42840));
    Span4Mux_v I__9753 (
            .O(N__42846),
            .I(N__42832));
    Span4Mux_v I__9752 (
            .O(N__42843),
            .I(N__42832));
    LocalMux I__9751 (
            .O(N__42840),
            .I(N__42832));
    CEMux I__9750 (
            .O(N__42839),
            .I(N__42829));
    Span4Mux_v I__9749 (
            .O(N__42832),
            .I(N__42826));
    LocalMux I__9748 (
            .O(N__42829),
            .I(N__42823));
    Span4Mux_h I__9747 (
            .O(N__42826),
            .I(N__42818));
    Span4Mux_v I__9746 (
            .O(N__42823),
            .I(N__42818));
    Span4Mux_v I__9745 (
            .O(N__42818),
            .I(N__42815));
    Odrv4 I__9744 (
            .O(N__42815),
            .I(\delay_measurement_inst.delay_tr_timer.N_324_i ));
    InMux I__9743 (
            .O(N__42812),
            .I(N__42809));
    LocalMux I__9742 (
            .O(N__42809),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_7_19 ));
    InMux I__9741 (
            .O(N__42806),
            .I(N__42803));
    LocalMux I__9740 (
            .O(N__42803),
            .I(N__42800));
    Odrv4 I__9739 (
            .O(N__42800),
            .I(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_4 ));
    InMux I__9738 (
            .O(N__42797),
            .I(N__42793));
    InMux I__9737 (
            .O(N__42796),
            .I(N__42790));
    LocalMux I__9736 (
            .O(N__42793),
            .I(N__42786));
    LocalMux I__9735 (
            .O(N__42790),
            .I(N__42783));
    InMux I__9734 (
            .O(N__42789),
            .I(N__42780));
    Span4Mux_v I__9733 (
            .O(N__42786),
            .I(N__42775));
    Span4Mux_v I__9732 (
            .O(N__42783),
            .I(N__42775));
    LocalMux I__9731 (
            .O(N__42780),
            .I(\delay_measurement_inst.elapsed_time_tr_2 ));
    Odrv4 I__9730 (
            .O(N__42775),
            .I(\delay_measurement_inst.elapsed_time_tr_2 ));
    InMux I__9729 (
            .O(N__42770),
            .I(N__42765));
    CascadeMux I__9728 (
            .O(N__42769),
            .I(N__42761));
    InMux I__9727 (
            .O(N__42768),
            .I(N__42758));
    LocalMux I__9726 (
            .O(N__42765),
            .I(N__42755));
    InMux I__9725 (
            .O(N__42764),
            .I(N__42752));
    InMux I__9724 (
            .O(N__42761),
            .I(N__42749));
    LocalMux I__9723 (
            .O(N__42758),
            .I(N__42744));
    Span4Mux_h I__9722 (
            .O(N__42755),
            .I(N__42744));
    LocalMux I__9721 (
            .O(N__42752),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16 ));
    LocalMux I__9720 (
            .O(N__42749),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16 ));
    Odrv4 I__9719 (
            .O(N__42744),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16 ));
    InMux I__9718 (
            .O(N__42737),
            .I(bfn_17_13_0_));
    InMux I__9717 (
            .O(N__42734),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ));
    InMux I__9716 (
            .O(N__42731),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ));
    InMux I__9715 (
            .O(N__42728),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ));
    InMux I__9714 (
            .O(N__42725),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ));
    InMux I__9713 (
            .O(N__42722),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ));
    InMux I__9712 (
            .O(N__42719),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ));
    InMux I__9711 (
            .O(N__42716),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ));
    InMux I__9710 (
            .O(N__42713),
            .I(bfn_17_14_0_));
    InMux I__9709 (
            .O(N__42710),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ));
    InMux I__9708 (
            .O(N__42707),
            .I(bfn_17_12_0_));
    InMux I__9707 (
            .O(N__42704),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ));
    InMux I__9706 (
            .O(N__42701),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ));
    InMux I__9705 (
            .O(N__42698),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ));
    InMux I__9704 (
            .O(N__42695),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ));
    InMux I__9703 (
            .O(N__42692),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ));
    InMux I__9702 (
            .O(N__42689),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ));
    InMux I__9701 (
            .O(N__42686),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ));
    CascadeMux I__9700 (
            .O(N__42683),
            .I(N__42679));
    CascadeMux I__9699 (
            .O(N__42682),
            .I(N__42676));
    InMux I__9698 (
            .O(N__42679),
            .I(N__42671));
    InMux I__9697 (
            .O(N__42676),
            .I(N__42671));
    LocalMux I__9696 (
            .O(N__42671),
            .I(N__42668));
    Span4Mux_v I__9695 (
            .O(N__42668),
            .I(N__42664));
    InMux I__9694 (
            .O(N__42667),
            .I(N__42661));
    Span4Mux_h I__9693 (
            .O(N__42664),
            .I(N__42658));
    LocalMux I__9692 (
            .O(N__42661),
            .I(measured_delay_hc_22));
    Odrv4 I__9691 (
            .O(N__42658),
            .I(measured_delay_hc_22));
    CascadeMux I__9690 (
            .O(N__42653),
            .I(N__42641));
    CascadeMux I__9689 (
            .O(N__42652),
            .I(N__42637));
    CascadeMux I__9688 (
            .O(N__42651),
            .I(N__42633));
    InMux I__9687 (
            .O(N__42650),
            .I(N__42615));
    InMux I__9686 (
            .O(N__42649),
            .I(N__42615));
    InMux I__9685 (
            .O(N__42648),
            .I(N__42612));
    InMux I__9684 (
            .O(N__42647),
            .I(N__42605));
    InMux I__9683 (
            .O(N__42646),
            .I(N__42605));
    InMux I__9682 (
            .O(N__42645),
            .I(N__42605));
    InMux I__9681 (
            .O(N__42644),
            .I(N__42594));
    InMux I__9680 (
            .O(N__42641),
            .I(N__42594));
    InMux I__9679 (
            .O(N__42640),
            .I(N__42594));
    InMux I__9678 (
            .O(N__42637),
            .I(N__42594));
    InMux I__9677 (
            .O(N__42636),
            .I(N__42594));
    InMux I__9676 (
            .O(N__42633),
            .I(N__42583));
    InMux I__9675 (
            .O(N__42632),
            .I(N__42583));
    InMux I__9674 (
            .O(N__42631),
            .I(N__42583));
    InMux I__9673 (
            .O(N__42630),
            .I(N__42583));
    InMux I__9672 (
            .O(N__42629),
            .I(N__42583));
    InMux I__9671 (
            .O(N__42628),
            .I(N__42574));
    InMux I__9670 (
            .O(N__42627),
            .I(N__42574));
    InMux I__9669 (
            .O(N__42626),
            .I(N__42574));
    InMux I__9668 (
            .O(N__42625),
            .I(N__42574));
    InMux I__9667 (
            .O(N__42624),
            .I(N__42571));
    InMux I__9666 (
            .O(N__42623),
            .I(N__42564));
    InMux I__9665 (
            .O(N__42622),
            .I(N__42564));
    InMux I__9664 (
            .O(N__42621),
            .I(N__42564));
    InMux I__9663 (
            .O(N__42620),
            .I(N__42561));
    LocalMux I__9662 (
            .O(N__42615),
            .I(N__42555));
    LocalMux I__9661 (
            .O(N__42612),
            .I(N__42552));
    LocalMux I__9660 (
            .O(N__42605),
            .I(N__42544));
    LocalMux I__9659 (
            .O(N__42594),
            .I(N__42544));
    LocalMux I__9658 (
            .O(N__42583),
            .I(N__42544));
    LocalMux I__9657 (
            .O(N__42574),
            .I(N__42535));
    LocalMux I__9656 (
            .O(N__42571),
            .I(N__42535));
    LocalMux I__9655 (
            .O(N__42564),
            .I(N__42535));
    LocalMux I__9654 (
            .O(N__42561),
            .I(N__42535));
    InMux I__9653 (
            .O(N__42560),
            .I(N__42528));
    InMux I__9652 (
            .O(N__42559),
            .I(N__42528));
    InMux I__9651 (
            .O(N__42558),
            .I(N__42528));
    Span4Mux_v I__9650 (
            .O(N__42555),
            .I(N__42522));
    Span4Mux_h I__9649 (
            .O(N__42552),
            .I(N__42519));
    InMux I__9648 (
            .O(N__42551),
            .I(N__42516));
    Span4Mux_v I__9647 (
            .O(N__42544),
            .I(N__42509));
    Span4Mux_v I__9646 (
            .O(N__42535),
            .I(N__42509));
    LocalMux I__9645 (
            .O(N__42528),
            .I(N__42509));
    InMux I__9644 (
            .O(N__42527),
            .I(N__42502));
    InMux I__9643 (
            .O(N__42526),
            .I(N__42502));
    InMux I__9642 (
            .O(N__42525),
            .I(N__42502));
    Odrv4 I__9641 (
            .O(N__42522),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    Odrv4 I__9640 (
            .O(N__42519),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    LocalMux I__9639 (
            .O(N__42516),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    Odrv4 I__9638 (
            .O(N__42509),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    LocalMux I__9637 (
            .O(N__42502),
            .I(\delay_measurement_inst.un1_elapsed_time_hc ));
    CascadeMux I__9636 (
            .O(N__42491),
            .I(N__42488));
    InMux I__9635 (
            .O(N__42488),
            .I(N__42485));
    LocalMux I__9634 (
            .O(N__42485),
            .I(N__42482));
    Span4Mux_h I__9633 (
            .O(N__42482),
            .I(N__42477));
    InMux I__9632 (
            .O(N__42481),
            .I(N__42472));
    InMux I__9631 (
            .O(N__42480),
            .I(N__42472));
    Odrv4 I__9630 (
            .O(N__42477),
            .I(\delay_measurement_inst.elapsed_time_hc_17 ));
    LocalMux I__9629 (
            .O(N__42472),
            .I(\delay_measurement_inst.elapsed_time_hc_17 ));
    InMux I__9628 (
            .O(N__42467),
            .I(N__42454));
    InMux I__9627 (
            .O(N__42466),
            .I(N__42454));
    InMux I__9626 (
            .O(N__42465),
            .I(N__42454));
    InMux I__9625 (
            .O(N__42464),
            .I(N__42447));
    InMux I__9624 (
            .O(N__42463),
            .I(N__42447));
    InMux I__9623 (
            .O(N__42462),
            .I(N__42447));
    InMux I__9622 (
            .O(N__42461),
            .I(N__42435));
    LocalMux I__9621 (
            .O(N__42454),
            .I(N__42432));
    LocalMux I__9620 (
            .O(N__42447),
            .I(N__42429));
    InMux I__9619 (
            .O(N__42446),
            .I(N__42422));
    InMux I__9618 (
            .O(N__42445),
            .I(N__42422));
    InMux I__9617 (
            .O(N__42444),
            .I(N__42422));
    InMux I__9616 (
            .O(N__42443),
            .I(N__42412));
    InMux I__9615 (
            .O(N__42442),
            .I(N__42412));
    InMux I__9614 (
            .O(N__42441),
            .I(N__42403));
    InMux I__9613 (
            .O(N__42440),
            .I(N__42403));
    InMux I__9612 (
            .O(N__42439),
            .I(N__42403));
    InMux I__9611 (
            .O(N__42438),
            .I(N__42403));
    LocalMux I__9610 (
            .O(N__42435),
            .I(N__42400));
    Span4Mux_v I__9609 (
            .O(N__42432),
            .I(N__42393));
    Span4Mux_v I__9608 (
            .O(N__42429),
            .I(N__42393));
    LocalMux I__9607 (
            .O(N__42422),
            .I(N__42393));
    InMux I__9606 (
            .O(N__42421),
            .I(N__42384));
    InMux I__9605 (
            .O(N__42420),
            .I(N__42384));
    InMux I__9604 (
            .O(N__42419),
            .I(N__42384));
    InMux I__9603 (
            .O(N__42418),
            .I(N__42384));
    InMux I__9602 (
            .O(N__42417),
            .I(N__42381));
    LocalMux I__9601 (
            .O(N__42412),
            .I(N__42375));
    LocalMux I__9600 (
            .O(N__42403),
            .I(N__42372));
    Span4Mux_v I__9599 (
            .O(N__42400),
            .I(N__42363));
    Span4Mux_h I__9598 (
            .O(N__42393),
            .I(N__42363));
    LocalMux I__9597 (
            .O(N__42384),
            .I(N__42363));
    LocalMux I__9596 (
            .O(N__42381),
            .I(N__42363));
    InMux I__9595 (
            .O(N__42380),
            .I(N__42356));
    InMux I__9594 (
            .O(N__42379),
            .I(N__42356));
    InMux I__9593 (
            .O(N__42378),
            .I(N__42356));
    Odrv4 I__9592 (
            .O(N__42375),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    Odrv12 I__9591 (
            .O(N__42372),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    Odrv4 I__9590 (
            .O(N__42363),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    LocalMux I__9589 (
            .O(N__42356),
            .I(\delay_measurement_inst.delay_hc_reg3 ));
    InMux I__9588 (
            .O(N__42347),
            .I(N__42343));
    InMux I__9587 (
            .O(N__42346),
            .I(N__42340));
    LocalMux I__9586 (
            .O(N__42343),
            .I(N__42336));
    LocalMux I__9585 (
            .O(N__42340),
            .I(N__42333));
    InMux I__9584 (
            .O(N__42339),
            .I(N__42330));
    Span4Mux_v I__9583 (
            .O(N__42336),
            .I(N__42326));
    Span4Mux_h I__9582 (
            .O(N__42333),
            .I(N__42323));
    LocalMux I__9581 (
            .O(N__42330),
            .I(N__42320));
    InMux I__9580 (
            .O(N__42329),
            .I(N__42316));
    Span4Mux_v I__9579 (
            .O(N__42326),
            .I(N__42311));
    Span4Mux_h I__9578 (
            .O(N__42323),
            .I(N__42311));
    Span4Mux_v I__9577 (
            .O(N__42320),
            .I(N__42308));
    InMux I__9576 (
            .O(N__42319),
            .I(N__42305));
    LocalMux I__9575 (
            .O(N__42316),
            .I(measured_delay_hc_17));
    Odrv4 I__9574 (
            .O(N__42311),
            .I(measured_delay_hc_17));
    Odrv4 I__9573 (
            .O(N__42308),
            .I(measured_delay_hc_17));
    LocalMux I__9572 (
            .O(N__42305),
            .I(measured_delay_hc_17));
    InMux I__9571 (
            .O(N__42296),
            .I(bfn_17_11_0_));
    InMux I__9570 (
            .O(N__42293),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ));
    InMux I__9569 (
            .O(N__42290),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ));
    InMux I__9568 (
            .O(N__42287),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ));
    InMux I__9567 (
            .O(N__42284),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ));
    InMux I__9566 (
            .O(N__42281),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ));
    InMux I__9565 (
            .O(N__42278),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ));
    CascadeMux I__9564 (
            .O(N__42275),
            .I(N__42271));
    InMux I__9563 (
            .O(N__42274),
            .I(N__42268));
    InMux I__9562 (
            .O(N__42271),
            .I(N__42265));
    LocalMux I__9561 (
            .O(N__42268),
            .I(measured_delay_hc_24));
    LocalMux I__9560 (
            .O(N__42265),
            .I(measured_delay_hc_24));
    CascadeMux I__9559 (
            .O(N__42260),
            .I(N__42256));
    CascadeMux I__9558 (
            .O(N__42259),
            .I(N__42253));
    InMux I__9557 (
            .O(N__42256),
            .I(N__42250));
    InMux I__9556 (
            .O(N__42253),
            .I(N__42247));
    LocalMux I__9555 (
            .O(N__42250),
            .I(N__42244));
    LocalMux I__9554 (
            .O(N__42247),
            .I(N__42240));
    Span4Mux_v I__9553 (
            .O(N__42244),
            .I(N__42237));
    InMux I__9552 (
            .O(N__42243),
            .I(N__42234));
    Span4Mux_v I__9551 (
            .O(N__42240),
            .I(N__42230));
    Span4Mux_h I__9550 (
            .O(N__42237),
            .I(N__42225));
    LocalMux I__9549 (
            .O(N__42234),
            .I(N__42225));
    InMux I__9548 (
            .O(N__42233),
            .I(N__42222));
    Span4Mux_v I__9547 (
            .O(N__42230),
            .I(N__42219));
    Span4Mux_h I__9546 (
            .O(N__42225),
            .I(N__42216));
    LocalMux I__9545 (
            .O(N__42222),
            .I(measured_delay_hc_0));
    Odrv4 I__9544 (
            .O(N__42219),
            .I(measured_delay_hc_0));
    Odrv4 I__9543 (
            .O(N__42216),
            .I(measured_delay_hc_0));
    InMux I__9542 (
            .O(N__42209),
            .I(N__42206));
    LocalMux I__9541 (
            .O(N__42206),
            .I(N__42201));
    InMux I__9540 (
            .O(N__42205),
            .I(N__42196));
    InMux I__9539 (
            .O(N__42204),
            .I(N__42196));
    Odrv4 I__9538 (
            .O(N__42201),
            .I(\delay_measurement_inst.elapsed_time_hc_18 ));
    LocalMux I__9537 (
            .O(N__42196),
            .I(\delay_measurement_inst.elapsed_time_hc_18 ));
    InMux I__9536 (
            .O(N__42191),
            .I(N__42187));
    InMux I__9535 (
            .O(N__42190),
            .I(N__42184));
    LocalMux I__9534 (
            .O(N__42187),
            .I(N__42178));
    LocalMux I__9533 (
            .O(N__42184),
            .I(N__42175));
    InMux I__9532 (
            .O(N__42183),
            .I(N__42172));
    CascadeMux I__9531 (
            .O(N__42182),
            .I(N__42169));
    CascadeMux I__9530 (
            .O(N__42181),
            .I(N__42166));
    Span4Mux_v I__9529 (
            .O(N__42178),
            .I(N__42163));
    Span4Mux_v I__9528 (
            .O(N__42175),
            .I(N__42160));
    LocalMux I__9527 (
            .O(N__42172),
            .I(N__42157));
    InMux I__9526 (
            .O(N__42169),
            .I(N__42154));
    InMux I__9525 (
            .O(N__42166),
            .I(N__42151));
    Span4Mux_h I__9524 (
            .O(N__42163),
            .I(N__42148));
    Span4Mux_v I__9523 (
            .O(N__42160),
            .I(N__42141));
    Span4Mux_h I__9522 (
            .O(N__42157),
            .I(N__42141));
    LocalMux I__9521 (
            .O(N__42154),
            .I(N__42141));
    LocalMux I__9520 (
            .O(N__42151),
            .I(measured_delay_hc_18));
    Odrv4 I__9519 (
            .O(N__42148),
            .I(measured_delay_hc_18));
    Odrv4 I__9518 (
            .O(N__42141),
            .I(measured_delay_hc_18));
    CascadeMux I__9517 (
            .O(N__42134),
            .I(N__42131));
    InMux I__9516 (
            .O(N__42131),
            .I(N__42126));
    InMux I__9515 (
            .O(N__42130),
            .I(N__42123));
    CascadeMux I__9514 (
            .O(N__42129),
            .I(N__42120));
    LocalMux I__9513 (
            .O(N__42126),
            .I(N__42117));
    LocalMux I__9512 (
            .O(N__42123),
            .I(N__42114));
    InMux I__9511 (
            .O(N__42120),
            .I(N__42111));
    Odrv4 I__9510 (
            .O(N__42117),
            .I(\delay_measurement_inst.elapsed_time_hc_19 ));
    Odrv4 I__9509 (
            .O(N__42114),
            .I(\delay_measurement_inst.elapsed_time_hc_19 ));
    LocalMux I__9508 (
            .O(N__42111),
            .I(\delay_measurement_inst.elapsed_time_hc_19 ));
    InMux I__9507 (
            .O(N__42104),
            .I(N__42094));
    InMux I__9506 (
            .O(N__42103),
            .I(N__42094));
    InMux I__9505 (
            .O(N__42102),
            .I(N__42089));
    InMux I__9504 (
            .O(N__42101),
            .I(N__42082));
    InMux I__9503 (
            .O(N__42100),
            .I(N__42082));
    InMux I__9502 (
            .O(N__42099),
            .I(N__42082));
    LocalMux I__9501 (
            .O(N__42094),
            .I(N__42079));
    InMux I__9500 (
            .O(N__42093),
            .I(N__42076));
    InMux I__9499 (
            .O(N__42092),
            .I(N__42073));
    LocalMux I__9498 (
            .O(N__42089),
            .I(N__42070));
    LocalMux I__9497 (
            .O(N__42082),
            .I(N__42067));
    Span4Mux_v I__9496 (
            .O(N__42079),
            .I(N__42062));
    LocalMux I__9495 (
            .O(N__42076),
            .I(N__42062));
    LocalMux I__9494 (
            .O(N__42073),
            .I(\delay_measurement_inst.delay_hc_reg3lto31_0_0 ));
    Odrv4 I__9493 (
            .O(N__42070),
            .I(\delay_measurement_inst.delay_hc_reg3lto31_0_0 ));
    Odrv4 I__9492 (
            .O(N__42067),
            .I(\delay_measurement_inst.delay_hc_reg3lto31_0_0 ));
    Odrv4 I__9491 (
            .O(N__42062),
            .I(\delay_measurement_inst.delay_hc_reg3lto31_0_0 ));
    CascadeMux I__9490 (
            .O(N__42053),
            .I(N__42050));
    InMux I__9489 (
            .O(N__42050),
            .I(N__42045));
    InMux I__9488 (
            .O(N__42049),
            .I(N__42042));
    InMux I__9487 (
            .O(N__42048),
            .I(N__42039));
    LocalMux I__9486 (
            .O(N__42045),
            .I(N__42036));
    LocalMux I__9485 (
            .O(N__42042),
            .I(N__42033));
    LocalMux I__9484 (
            .O(N__42039),
            .I(N__42028));
    Span4Mux_v I__9483 (
            .O(N__42036),
            .I(N__42028));
    Span4Mux_v I__9482 (
            .O(N__42033),
            .I(N__42025));
    Odrv4 I__9481 (
            .O(N__42028),
            .I(measured_delay_hc_19));
    Odrv4 I__9480 (
            .O(N__42025),
            .I(measured_delay_hc_19));
    InMux I__9479 (
            .O(N__42020),
            .I(N__42014));
    InMux I__9478 (
            .O(N__42019),
            .I(N__42014));
    LocalMux I__9477 (
            .O(N__42014),
            .I(N__42010));
    InMux I__9476 (
            .O(N__42013),
            .I(N__42007));
    Span4Mux_h I__9475 (
            .O(N__42010),
            .I(N__42004));
    LocalMux I__9474 (
            .O(N__42007),
            .I(measured_delay_hc_21));
    Odrv4 I__9473 (
            .O(N__42004),
            .I(measured_delay_hc_21));
    InMux I__9472 (
            .O(N__41999),
            .I(N__41995));
    InMux I__9471 (
            .O(N__41998),
            .I(N__41992));
    LocalMux I__9470 (
            .O(N__41995),
            .I(N__41988));
    LocalMux I__9469 (
            .O(N__41992),
            .I(N__41985));
    CascadeMux I__9468 (
            .O(N__41991),
            .I(N__41982));
    Span4Mux_v I__9467 (
            .O(N__41988),
            .I(N__41979));
    Span4Mux_v I__9466 (
            .O(N__41985),
            .I(N__41976));
    InMux I__9465 (
            .O(N__41982),
            .I(N__41973));
    Odrv4 I__9464 (
            .O(N__41979),
            .I(measured_delay_tr_13));
    Odrv4 I__9463 (
            .O(N__41976),
            .I(measured_delay_tr_13));
    LocalMux I__9462 (
            .O(N__41973),
            .I(measured_delay_tr_13));
    CascadeMux I__9461 (
            .O(N__41966),
            .I(N__41963));
    InMux I__9460 (
            .O(N__41963),
            .I(N__41960));
    LocalMux I__9459 (
            .O(N__41960),
            .I(N__41957));
    Odrv12 I__9458 (
            .O(N__41957),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ));
    InMux I__9457 (
            .O(N__41954),
            .I(N__41951));
    LocalMux I__9456 (
            .O(N__41951),
            .I(N__41948));
    Odrv12 I__9455 (
            .O(N__41948),
            .I(delay_hc_input_c));
    InMux I__9454 (
            .O(N__41945),
            .I(N__41942));
    LocalMux I__9453 (
            .O(N__41942),
            .I(delay_hc_d1));
    InMux I__9452 (
            .O(N__41939),
            .I(N__41936));
    LocalMux I__9451 (
            .O(N__41936),
            .I(N__41933));
    Span4Mux_v I__9450 (
            .O(N__41933),
            .I(N__41927));
    InMux I__9449 (
            .O(N__41932),
            .I(N__41922));
    InMux I__9448 (
            .O(N__41931),
            .I(N__41922));
    InMux I__9447 (
            .O(N__41930),
            .I(N__41919));
    Span4Mux_h I__9446 (
            .O(N__41927),
            .I(N__41916));
    LocalMux I__9445 (
            .O(N__41922),
            .I(N__41913));
    LocalMux I__9444 (
            .O(N__41919),
            .I(N__41910));
    Span4Mux_v I__9443 (
            .O(N__41916),
            .I(N__41907));
    Span12Mux_v I__9442 (
            .O(N__41913),
            .I(N__41904));
    Span4Mux_v I__9441 (
            .O(N__41910),
            .I(N__41901));
    Odrv4 I__9440 (
            .O(N__41907),
            .I(delay_hc_d2));
    Odrv12 I__9439 (
            .O(N__41904),
            .I(delay_hc_d2));
    Odrv4 I__9438 (
            .O(N__41901),
            .I(delay_hc_d2));
    InMux I__9437 (
            .O(N__41894),
            .I(N__41891));
    LocalMux I__9436 (
            .O(N__41891),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_3 ));
    InMux I__9435 (
            .O(N__41888),
            .I(N__41883));
    InMux I__9434 (
            .O(N__41887),
            .I(N__41880));
    InMux I__9433 (
            .O(N__41886),
            .I(N__41877));
    LocalMux I__9432 (
            .O(N__41883),
            .I(N__41873));
    LocalMux I__9431 (
            .O(N__41880),
            .I(N__41870));
    LocalMux I__9430 (
            .O(N__41877),
            .I(N__41867));
    InMux I__9429 (
            .O(N__41876),
            .I(N__41864));
    Span4Mux_v I__9428 (
            .O(N__41873),
            .I(N__41861));
    Sp12to4 I__9427 (
            .O(N__41870),
            .I(N__41856));
    Sp12to4 I__9426 (
            .O(N__41867),
            .I(N__41856));
    LocalMux I__9425 (
            .O(N__41864),
            .I(N__41853));
    Sp12to4 I__9424 (
            .O(N__41861),
            .I(N__41850));
    Span12Mux_v I__9423 (
            .O(N__41856),
            .I(N__41847));
    Span4Mux_v I__9422 (
            .O(N__41853),
            .I(N__41844));
    Odrv12 I__9421 (
            .O(N__41850),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_2 ));
    Odrv12 I__9420 (
            .O(N__41847),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_2 ));
    Odrv4 I__9419 (
            .O(N__41844),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_2 ));
    InMux I__9418 (
            .O(N__41837),
            .I(N__41833));
    InMux I__9417 (
            .O(N__41836),
            .I(N__41830));
    LocalMux I__9416 (
            .O(N__41833),
            .I(measured_delay_hc_25));
    LocalMux I__9415 (
            .O(N__41830),
            .I(measured_delay_hc_25));
    InMux I__9414 (
            .O(N__41825),
            .I(N__41821));
    InMux I__9413 (
            .O(N__41824),
            .I(N__41818));
    LocalMux I__9412 (
            .O(N__41821),
            .I(measured_delay_hc_26));
    LocalMux I__9411 (
            .O(N__41818),
            .I(measured_delay_hc_26));
    CascadeMux I__9410 (
            .O(N__41813),
            .I(N__41810));
    InMux I__9409 (
            .O(N__41810),
            .I(N__41804));
    InMux I__9408 (
            .O(N__41809),
            .I(N__41804));
    LocalMux I__9407 (
            .O(N__41804),
            .I(measured_delay_hc_23));
    InMux I__9406 (
            .O(N__41801),
            .I(N__41798));
    LocalMux I__9405 (
            .O(N__41798),
            .I(N__41794));
    CascadeMux I__9404 (
            .O(N__41797),
            .I(N__41789));
    Span4Mux_v I__9403 (
            .O(N__41794),
            .I(N__41786));
    InMux I__9402 (
            .O(N__41793),
            .I(N__41783));
    InMux I__9401 (
            .O(N__41792),
            .I(N__41780));
    InMux I__9400 (
            .O(N__41789),
            .I(N__41777));
    Odrv4 I__9399 (
            .O(N__41786),
            .I(\delay_measurement_inst.elapsed_time_hc_8 ));
    LocalMux I__9398 (
            .O(N__41783),
            .I(\delay_measurement_inst.elapsed_time_hc_8 ));
    LocalMux I__9397 (
            .O(N__41780),
            .I(\delay_measurement_inst.elapsed_time_hc_8 ));
    LocalMux I__9396 (
            .O(N__41777),
            .I(\delay_measurement_inst.elapsed_time_hc_8 ));
    InMux I__9395 (
            .O(N__41768),
            .I(N__41764));
    InMux I__9394 (
            .O(N__41767),
            .I(N__41760));
    LocalMux I__9393 (
            .O(N__41764),
            .I(N__41757));
    CascadeMux I__9392 (
            .O(N__41763),
            .I(N__41753));
    LocalMux I__9391 (
            .O(N__41760),
            .I(N__41750));
    Span4Mux_v I__9390 (
            .O(N__41757),
            .I(N__41747));
    InMux I__9389 (
            .O(N__41756),
            .I(N__41744));
    InMux I__9388 (
            .O(N__41753),
            .I(N__41741));
    Span4Mux_v I__9387 (
            .O(N__41750),
            .I(N__41737));
    Span4Mux_h I__9386 (
            .O(N__41747),
            .I(N__41734));
    LocalMux I__9385 (
            .O(N__41744),
            .I(N__41731));
    LocalMux I__9384 (
            .O(N__41741),
            .I(N__41728));
    InMux I__9383 (
            .O(N__41740),
            .I(N__41725));
    Span4Mux_v I__9382 (
            .O(N__41737),
            .I(N__41722));
    Span4Mux_h I__9381 (
            .O(N__41734),
            .I(N__41715));
    Span4Mux_v I__9380 (
            .O(N__41731),
            .I(N__41715));
    Span4Mux_v I__9379 (
            .O(N__41728),
            .I(N__41715));
    LocalMux I__9378 (
            .O(N__41725),
            .I(measured_delay_hc_8));
    Odrv4 I__9377 (
            .O(N__41722),
            .I(measured_delay_hc_8));
    Odrv4 I__9376 (
            .O(N__41715),
            .I(measured_delay_hc_8));
    CascadeMux I__9375 (
            .O(N__41708),
            .I(N__41705));
    InMux I__9374 (
            .O(N__41705),
            .I(N__41702));
    LocalMux I__9373 (
            .O(N__41702),
            .I(N__41699));
    Span4Mux_v I__9372 (
            .O(N__41699),
            .I(N__41693));
    InMux I__9371 (
            .O(N__41698),
            .I(N__41690));
    InMux I__9370 (
            .O(N__41697),
            .I(N__41687));
    InMux I__9369 (
            .O(N__41696),
            .I(N__41684));
    Odrv4 I__9368 (
            .O(N__41693),
            .I(\delay_measurement_inst.elapsed_time_hc_7 ));
    LocalMux I__9367 (
            .O(N__41690),
            .I(\delay_measurement_inst.elapsed_time_hc_7 ));
    LocalMux I__9366 (
            .O(N__41687),
            .I(\delay_measurement_inst.elapsed_time_hc_7 ));
    LocalMux I__9365 (
            .O(N__41684),
            .I(\delay_measurement_inst.elapsed_time_hc_7 ));
    InMux I__9364 (
            .O(N__41675),
            .I(N__41672));
    LocalMux I__9363 (
            .O(N__41672),
            .I(N__41667));
    InMux I__9362 (
            .O(N__41671),
            .I(N__41664));
    InMux I__9361 (
            .O(N__41670),
            .I(N__41661));
    Span4Mux_v I__9360 (
            .O(N__41667),
            .I(N__41655));
    LocalMux I__9359 (
            .O(N__41664),
            .I(N__41655));
    LocalMux I__9358 (
            .O(N__41661),
            .I(N__41652));
    InMux I__9357 (
            .O(N__41660),
            .I(N__41649));
    Span4Mux_v I__9356 (
            .O(N__41655),
            .I(N__41645));
    Span4Mux_h I__9355 (
            .O(N__41652),
            .I(N__41640));
    LocalMux I__9354 (
            .O(N__41649),
            .I(N__41640));
    InMux I__9353 (
            .O(N__41648),
            .I(N__41637));
    Span4Mux_h I__9352 (
            .O(N__41645),
            .I(N__41634));
    Span4Mux_h I__9351 (
            .O(N__41640),
            .I(N__41631));
    LocalMux I__9350 (
            .O(N__41637),
            .I(measured_delay_hc_7));
    Odrv4 I__9349 (
            .O(N__41634),
            .I(measured_delay_hc_7));
    Odrv4 I__9348 (
            .O(N__41631),
            .I(measured_delay_hc_7));
    InMux I__9347 (
            .O(N__41624),
            .I(N__41621));
    LocalMux I__9346 (
            .O(N__41621),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_16 ));
    CascadeMux I__9345 (
            .O(N__41618),
            .I(N__41615));
    InMux I__9344 (
            .O(N__41615),
            .I(N__41612));
    LocalMux I__9343 (
            .O(N__41612),
            .I(N__41609));
    Odrv4 I__9342 (
            .O(N__41609),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ));
    InMux I__9341 (
            .O(N__41606),
            .I(N__41603));
    LocalMux I__9340 (
            .O(N__41603),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_17 ));
    InMux I__9339 (
            .O(N__41600),
            .I(N__41597));
    LocalMux I__9338 (
            .O(N__41597),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_18 ));
    InMux I__9337 (
            .O(N__41594),
            .I(N__41591));
    LocalMux I__9336 (
            .O(N__41591),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_19 ));
    InMux I__9335 (
            .O(N__41588),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ));
    CascadeMux I__9334 (
            .O(N__41585),
            .I(N__41582));
    InMux I__9333 (
            .O(N__41582),
            .I(N__41579));
    LocalMux I__9332 (
            .O(N__41579),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ));
    InMux I__9331 (
            .O(N__41576),
            .I(N__41572));
    CascadeMux I__9330 (
            .O(N__41575),
            .I(N__41569));
    LocalMux I__9329 (
            .O(N__41572),
            .I(N__41564));
    InMux I__9328 (
            .O(N__41569),
            .I(N__41559));
    InMux I__9327 (
            .O(N__41568),
            .I(N__41559));
    InMux I__9326 (
            .O(N__41567),
            .I(N__41556));
    Span4Mux_v I__9325 (
            .O(N__41564),
            .I(N__41551));
    LocalMux I__9324 (
            .O(N__41559),
            .I(N__41551));
    LocalMux I__9323 (
            .O(N__41556),
            .I(N__41548));
    Span4Mux_v I__9322 (
            .O(N__41551),
            .I(N__41545));
    Odrv12 I__9321 (
            .O(N__41548),
            .I(measured_delay_tr_19));
    Odrv4 I__9320 (
            .O(N__41545),
            .I(measured_delay_tr_19));
    CascadeMux I__9319 (
            .O(N__41540),
            .I(N__41537));
    InMux I__9318 (
            .O(N__41537),
            .I(N__41534));
    LocalMux I__9317 (
            .O(N__41534),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ));
    InMux I__9316 (
            .O(N__41531),
            .I(N__41528));
    LocalMux I__9315 (
            .O(N__41528),
            .I(N__41524));
    InMux I__9314 (
            .O(N__41527),
            .I(N__41521));
    Span4Mux_h I__9313 (
            .O(N__41524),
            .I(N__41517));
    LocalMux I__9312 (
            .O(N__41521),
            .I(N__41514));
    InMux I__9311 (
            .O(N__41520),
            .I(N__41511));
    Odrv4 I__9310 (
            .O(N__41517),
            .I(measured_delay_tr_11));
    Odrv12 I__9309 (
            .O(N__41514),
            .I(measured_delay_tr_11));
    LocalMux I__9308 (
            .O(N__41511),
            .I(measured_delay_tr_11));
    CascadeMux I__9307 (
            .O(N__41504),
            .I(N__41501));
    InMux I__9306 (
            .O(N__41501),
            .I(N__41498));
    LocalMux I__9305 (
            .O(N__41498),
            .I(N__41495));
    Odrv4 I__9304 (
            .O(N__41495),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ));
    CascadeMux I__9303 (
            .O(N__41492),
            .I(N__41486));
    InMux I__9302 (
            .O(N__41491),
            .I(N__41476));
    InMux I__9301 (
            .O(N__41490),
            .I(N__41473));
    InMux I__9300 (
            .O(N__41489),
            .I(N__41470));
    InMux I__9299 (
            .O(N__41486),
            .I(N__41457));
    InMux I__9298 (
            .O(N__41485),
            .I(N__41457));
    InMux I__9297 (
            .O(N__41484),
            .I(N__41457));
    InMux I__9296 (
            .O(N__41483),
            .I(N__41457));
    InMux I__9295 (
            .O(N__41482),
            .I(N__41457));
    InMux I__9294 (
            .O(N__41481),
            .I(N__41457));
    CascadeMux I__9293 (
            .O(N__41480),
            .I(N__41454));
    CascadeMux I__9292 (
            .O(N__41479),
            .I(N__41448));
    LocalMux I__9291 (
            .O(N__41476),
            .I(N__41444));
    LocalMux I__9290 (
            .O(N__41473),
            .I(N__41441));
    LocalMux I__9289 (
            .O(N__41470),
            .I(N__41438));
    LocalMux I__9288 (
            .O(N__41457),
            .I(N__41434));
    InMux I__9287 (
            .O(N__41454),
            .I(N__41425));
    InMux I__9286 (
            .O(N__41453),
            .I(N__41425));
    InMux I__9285 (
            .O(N__41452),
            .I(N__41425));
    InMux I__9284 (
            .O(N__41451),
            .I(N__41425));
    InMux I__9283 (
            .O(N__41448),
            .I(N__41420));
    InMux I__9282 (
            .O(N__41447),
            .I(N__41420));
    Span4Mux_v I__9281 (
            .O(N__41444),
            .I(N__41415));
    Span4Mux_v I__9280 (
            .O(N__41441),
            .I(N__41415));
    Span12Mux_h I__9279 (
            .O(N__41438),
            .I(N__41412));
    InMux I__9278 (
            .O(N__41437),
            .I(N__41409));
    Span4Mux_h I__9277 (
            .O(N__41434),
            .I(N__41406));
    LocalMux I__9276 (
            .O(N__41425),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15 ));
    LocalMux I__9275 (
            .O(N__41420),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15 ));
    Odrv4 I__9274 (
            .O(N__41415),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15 ));
    Odrv12 I__9273 (
            .O(N__41412),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15 ));
    LocalMux I__9272 (
            .O(N__41409),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15 ));
    Odrv4 I__9271 (
            .O(N__41406),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15 ));
    CascadeMux I__9270 (
            .O(N__41393),
            .I(N__41390));
    InMux I__9269 (
            .O(N__41390),
            .I(N__41387));
    LocalMux I__9268 (
            .O(N__41387),
            .I(N__41384));
    Odrv4 I__9267 (
            .O(N__41384),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ));
    CascadeMux I__9266 (
            .O(N__41381),
            .I(N__41378));
    InMux I__9265 (
            .O(N__41378),
            .I(N__41375));
    LocalMux I__9264 (
            .O(N__41375),
            .I(N__41372));
    Odrv4 I__9263 (
            .O(N__41372),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ));
    InMux I__9262 (
            .O(N__41369),
            .I(N__41366));
    LocalMux I__9261 (
            .O(N__41366),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ));
    InMux I__9260 (
            .O(N__41363),
            .I(N__41360));
    LocalMux I__9259 (
            .O(N__41360),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ));
    CascadeMux I__9258 (
            .O(N__41357),
            .I(N__41354));
    InMux I__9257 (
            .O(N__41354),
            .I(N__41351));
    LocalMux I__9256 (
            .O(N__41351),
            .I(N__41348));
    Span4Mux_h I__9255 (
            .O(N__41348),
            .I(N__41345));
    Span4Mux_v I__9254 (
            .O(N__41345),
            .I(N__41342));
    Odrv4 I__9253 (
            .O(N__41342),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ));
    InMux I__9252 (
            .O(N__41339),
            .I(N__41336));
    LocalMux I__9251 (
            .O(N__41336),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ));
    InMux I__9250 (
            .O(N__41333),
            .I(N__41330));
    LocalMux I__9249 (
            .O(N__41330),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ));
    CascadeMux I__9248 (
            .O(N__41327),
            .I(N__41324));
    InMux I__9247 (
            .O(N__41324),
            .I(N__41321));
    LocalMux I__9246 (
            .O(N__41321),
            .I(N__41318));
    Span4Mux_h I__9245 (
            .O(N__41318),
            .I(N__41315));
    Span4Mux_v I__9244 (
            .O(N__41315),
            .I(N__41312));
    Odrv4 I__9243 (
            .O(N__41312),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ));
    InMux I__9242 (
            .O(N__41309),
            .I(N__41306));
    LocalMux I__9241 (
            .O(N__41306),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ));
    InMux I__9240 (
            .O(N__41303),
            .I(N__41300));
    LocalMux I__9239 (
            .O(N__41300),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ));
    CascadeMux I__9238 (
            .O(N__41297),
            .I(N__41294));
    InMux I__9237 (
            .O(N__41294),
            .I(N__41291));
    LocalMux I__9236 (
            .O(N__41291),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ));
    InMux I__9235 (
            .O(N__41288),
            .I(N__41285));
    LocalMux I__9234 (
            .O(N__41285),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ));
    InMux I__9233 (
            .O(N__41282),
            .I(N__41279));
    LocalMux I__9232 (
            .O(N__41279),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ));
    CascadeMux I__9231 (
            .O(N__41276),
            .I(N__41272));
    CascadeMux I__9230 (
            .O(N__41275),
            .I(N__41269));
    InMux I__9229 (
            .O(N__41272),
            .I(N__41266));
    InMux I__9228 (
            .O(N__41269),
            .I(N__41263));
    LocalMux I__9227 (
            .O(N__41266),
            .I(N__41260));
    LocalMux I__9226 (
            .O(N__41263),
            .I(N__41257));
    Span4Mux_v I__9225 (
            .O(N__41260),
            .I(N__41254));
    Span4Mux_h I__9224 (
            .O(N__41257),
            .I(N__41249));
    Span4Mux_h I__9223 (
            .O(N__41254),
            .I(N__41245));
    InMux I__9222 (
            .O(N__41253),
            .I(N__41242));
    CascadeMux I__9221 (
            .O(N__41252),
            .I(N__41239));
    Span4Mux_v I__9220 (
            .O(N__41249),
            .I(N__41236));
    InMux I__9219 (
            .O(N__41248),
            .I(N__41233));
    Span4Mux_h I__9218 (
            .O(N__41245),
            .I(N__41228));
    LocalMux I__9217 (
            .O(N__41242),
            .I(N__41228));
    InMux I__9216 (
            .O(N__41239),
            .I(N__41225));
    Span4Mux_v I__9215 (
            .O(N__41236),
            .I(N__41220));
    LocalMux I__9214 (
            .O(N__41233),
            .I(N__41220));
    Span4Mux_v I__9213 (
            .O(N__41228),
            .I(N__41217));
    LocalMux I__9212 (
            .O(N__41225),
            .I(measured_delay_hc_1));
    Odrv4 I__9211 (
            .O(N__41220),
            .I(measured_delay_hc_1));
    Odrv4 I__9210 (
            .O(N__41217),
            .I(measured_delay_hc_1));
    CascadeMux I__9209 (
            .O(N__41210),
            .I(N__41207));
    InMux I__9208 (
            .O(N__41207),
            .I(N__41204));
    LocalMux I__9207 (
            .O(N__41204),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_1 ));
    CascadeMux I__9206 (
            .O(N__41201),
            .I(N__41198));
    InMux I__9205 (
            .O(N__41198),
            .I(N__41195));
    LocalMux I__9204 (
            .O(N__41195),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ));
    InMux I__9203 (
            .O(N__41192),
            .I(N__41189));
    LocalMux I__9202 (
            .O(N__41189),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ));
    InMux I__9201 (
            .O(N__41186),
            .I(N__41183));
    LocalMux I__9200 (
            .O(N__41183),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ));
    CascadeMux I__9199 (
            .O(N__41180),
            .I(N__41177));
    InMux I__9198 (
            .O(N__41177),
            .I(N__41174));
    LocalMux I__9197 (
            .O(N__41174),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ));
    CascadeMux I__9196 (
            .O(N__41171),
            .I(N__41168));
    InMux I__9195 (
            .O(N__41168),
            .I(N__41165));
    LocalMux I__9194 (
            .O(N__41165),
            .I(N__41162));
    Span4Mux_h I__9193 (
            .O(N__41162),
            .I(N__41159));
    Odrv4 I__9192 (
            .O(N__41159),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ));
    InMux I__9191 (
            .O(N__41156),
            .I(N__41153));
    LocalMux I__9190 (
            .O(N__41153),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ));
    CascadeMux I__9189 (
            .O(N__41150),
            .I(N__41147));
    InMux I__9188 (
            .O(N__41147),
            .I(N__41144));
    LocalMux I__9187 (
            .O(N__41144),
            .I(N__41141));
    Odrv4 I__9186 (
            .O(N__41141),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ));
    InMux I__9185 (
            .O(N__41138),
            .I(N__41135));
    LocalMux I__9184 (
            .O(N__41135),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ));
    CascadeMux I__9183 (
            .O(N__41132),
            .I(N__41129));
    InMux I__9182 (
            .O(N__41129),
            .I(N__41126));
    LocalMux I__9181 (
            .O(N__41126),
            .I(N__41123));
    Span4Mux_h I__9180 (
            .O(N__41123),
            .I(N__41120));
    Odrv4 I__9179 (
            .O(N__41120),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ));
    InMux I__9178 (
            .O(N__41117),
            .I(N__41114));
    LocalMux I__9177 (
            .O(N__41114),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ));
    CascadeMux I__9176 (
            .O(N__41111),
            .I(N__41108));
    InMux I__9175 (
            .O(N__41108),
            .I(N__41105));
    LocalMux I__9174 (
            .O(N__41105),
            .I(N__41102));
    Span4Mux_h I__9173 (
            .O(N__41102),
            .I(N__41099));
    Odrv4 I__9172 (
            .O(N__41099),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ));
    InMux I__9171 (
            .O(N__41096),
            .I(N__41093));
    LocalMux I__9170 (
            .O(N__41093),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ));
    CascadeMux I__9169 (
            .O(N__41090),
            .I(N__41087));
    InMux I__9168 (
            .O(N__41087),
            .I(N__41084));
    LocalMux I__9167 (
            .O(N__41084),
            .I(N__41081));
    Span4Mux_v I__9166 (
            .O(N__41081),
            .I(N__41078));
    Odrv4 I__9165 (
            .O(N__41078),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ));
    InMux I__9164 (
            .O(N__41075),
            .I(N__41072));
    LocalMux I__9163 (
            .O(N__41072),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ));
    CascadeMux I__9162 (
            .O(N__41069),
            .I(N__41055));
    InMux I__9161 (
            .O(N__41068),
            .I(N__41046));
    InMux I__9160 (
            .O(N__41067),
            .I(N__41046));
    InMux I__9159 (
            .O(N__41066),
            .I(N__41046));
    InMux I__9158 (
            .O(N__41065),
            .I(N__41037));
    InMux I__9157 (
            .O(N__41064),
            .I(N__41037));
    InMux I__9156 (
            .O(N__41063),
            .I(N__41037));
    InMux I__9155 (
            .O(N__41062),
            .I(N__41037));
    InMux I__9154 (
            .O(N__41061),
            .I(N__41030));
    InMux I__9153 (
            .O(N__41060),
            .I(N__41030));
    InMux I__9152 (
            .O(N__41059),
            .I(N__41030));
    InMux I__9151 (
            .O(N__41058),
            .I(N__41023));
    InMux I__9150 (
            .O(N__41055),
            .I(N__41018));
    InMux I__9149 (
            .O(N__41054),
            .I(N__41015));
    InMux I__9148 (
            .O(N__41053),
            .I(N__41012));
    LocalMux I__9147 (
            .O(N__41046),
            .I(N__41009));
    LocalMux I__9146 (
            .O(N__41037),
            .I(N__41004));
    LocalMux I__9145 (
            .O(N__41030),
            .I(N__41004));
    CascadeMux I__9144 (
            .O(N__41029),
            .I(N__41001));
    InMux I__9143 (
            .O(N__41028),
            .I(N__40991));
    InMux I__9142 (
            .O(N__41027),
            .I(N__40991));
    InMux I__9141 (
            .O(N__41026),
            .I(N__40991));
    LocalMux I__9140 (
            .O(N__41023),
            .I(N__40988));
    InMux I__9139 (
            .O(N__41022),
            .I(N__40985));
    InMux I__9138 (
            .O(N__41021),
            .I(N__40982));
    LocalMux I__9137 (
            .O(N__41018),
            .I(N__40970));
    LocalMux I__9136 (
            .O(N__41015),
            .I(N__40970));
    LocalMux I__9135 (
            .O(N__41012),
            .I(N__40970));
    Span4Mux_v I__9134 (
            .O(N__41009),
            .I(N__40970));
    Span4Mux_v I__9133 (
            .O(N__41004),
            .I(N__40970));
    InMux I__9132 (
            .O(N__41001),
            .I(N__40961));
    InMux I__9131 (
            .O(N__41000),
            .I(N__40961));
    InMux I__9130 (
            .O(N__40999),
            .I(N__40961));
    InMux I__9129 (
            .O(N__40998),
            .I(N__40961));
    LocalMux I__9128 (
            .O(N__40991),
            .I(N__40956));
    Span4Mux_v I__9127 (
            .O(N__40988),
            .I(N__40956));
    LocalMux I__9126 (
            .O(N__40985),
            .I(N__40953));
    LocalMux I__9125 (
            .O(N__40982),
            .I(N__40950));
    InMux I__9124 (
            .O(N__40981),
            .I(N__40947));
    Span4Mux_v I__9123 (
            .O(N__40970),
            .I(N__40942));
    LocalMux I__9122 (
            .O(N__40961),
            .I(N__40942));
    Span4Mux_v I__9121 (
            .O(N__40956),
            .I(N__40937));
    Span4Mux_h I__9120 (
            .O(N__40953),
            .I(N__40937));
    Span4Mux_v I__9119 (
            .O(N__40950),
            .I(N__40934));
    LocalMux I__9118 (
            .O(N__40947),
            .I(N__40929));
    Span4Mux_v I__9117 (
            .O(N__40942),
            .I(N__40929));
    Span4Mux_v I__9116 (
            .O(N__40937),
            .I(N__40926));
    Odrv4 I__9115 (
            .O(N__40934),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__9114 (
            .O(N__40929),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__9113 (
            .O(N__40926),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ));
    CascadeMux I__9112 (
            .O(N__40919),
            .I(N__40911));
    CascadeMux I__9111 (
            .O(N__40918),
            .I(N__40906));
    CascadeMux I__9110 (
            .O(N__40917),
            .I(N__40903));
    CascadeMux I__9109 (
            .O(N__40916),
            .I(N__40896));
    CascadeMux I__9108 (
            .O(N__40915),
            .I(N__40891));
    CascadeMux I__9107 (
            .O(N__40914),
            .I(N__40888));
    InMux I__9106 (
            .O(N__40911),
            .I(N__40885));
    CascadeMux I__9105 (
            .O(N__40910),
            .I(N__40882));
    CascadeMux I__9104 (
            .O(N__40909),
            .I(N__40879));
    InMux I__9103 (
            .O(N__40906),
            .I(N__40876));
    InMux I__9102 (
            .O(N__40903),
            .I(N__40873));
    CascadeMux I__9101 (
            .O(N__40902),
            .I(N__40869));
    CascadeMux I__9100 (
            .O(N__40901),
            .I(N__40866));
    CascadeMux I__9099 (
            .O(N__40900),
            .I(N__40863));
    CascadeMux I__9098 (
            .O(N__40899),
            .I(N__40854));
    InMux I__9097 (
            .O(N__40896),
            .I(N__40849));
    InMux I__9096 (
            .O(N__40895),
            .I(N__40842));
    InMux I__9095 (
            .O(N__40894),
            .I(N__40842));
    InMux I__9094 (
            .O(N__40891),
            .I(N__40842));
    InMux I__9093 (
            .O(N__40888),
            .I(N__40839));
    LocalMux I__9092 (
            .O(N__40885),
            .I(N__40836));
    InMux I__9091 (
            .O(N__40882),
            .I(N__40831));
    InMux I__9090 (
            .O(N__40879),
            .I(N__40831));
    LocalMux I__9089 (
            .O(N__40876),
            .I(N__40826));
    LocalMux I__9088 (
            .O(N__40873),
            .I(N__40826));
    InMux I__9087 (
            .O(N__40872),
            .I(N__40821));
    InMux I__9086 (
            .O(N__40869),
            .I(N__40821));
    InMux I__9085 (
            .O(N__40866),
            .I(N__40812));
    InMux I__9084 (
            .O(N__40863),
            .I(N__40812));
    InMux I__9083 (
            .O(N__40862),
            .I(N__40812));
    InMux I__9082 (
            .O(N__40861),
            .I(N__40812));
    InMux I__9081 (
            .O(N__40860),
            .I(N__40803));
    InMux I__9080 (
            .O(N__40859),
            .I(N__40803));
    InMux I__9079 (
            .O(N__40858),
            .I(N__40803));
    InMux I__9078 (
            .O(N__40857),
            .I(N__40803));
    InMux I__9077 (
            .O(N__40854),
            .I(N__40795));
    InMux I__9076 (
            .O(N__40853),
            .I(N__40795));
    InMux I__9075 (
            .O(N__40852),
            .I(N__40795));
    LocalMux I__9074 (
            .O(N__40849),
            .I(N__40792));
    LocalMux I__9073 (
            .O(N__40842),
            .I(N__40789));
    LocalMux I__9072 (
            .O(N__40839),
            .I(N__40784));
    Span4Mux_h I__9071 (
            .O(N__40836),
            .I(N__40784));
    LocalMux I__9070 (
            .O(N__40831),
            .I(N__40775));
    Span4Mux_h I__9069 (
            .O(N__40826),
            .I(N__40775));
    LocalMux I__9068 (
            .O(N__40821),
            .I(N__40775));
    LocalMux I__9067 (
            .O(N__40812),
            .I(N__40775));
    LocalMux I__9066 (
            .O(N__40803),
            .I(N__40772));
    InMux I__9065 (
            .O(N__40802),
            .I(N__40769));
    LocalMux I__9064 (
            .O(N__40795),
            .I(N__40766));
    Span4Mux_v I__9063 (
            .O(N__40792),
            .I(N__40763));
    Span4Mux_h I__9062 (
            .O(N__40789),
            .I(N__40760));
    Span4Mux_v I__9061 (
            .O(N__40784),
            .I(N__40755));
    Span4Mux_v I__9060 (
            .O(N__40775),
            .I(N__40755));
    Span4Mux_h I__9059 (
            .O(N__40772),
            .I(N__40752));
    LocalMux I__9058 (
            .O(N__40769),
            .I(\phase_controller_slave.start_timer_hcZ0 ));
    Odrv12 I__9057 (
            .O(N__40766),
            .I(\phase_controller_slave.start_timer_hcZ0 ));
    Odrv4 I__9056 (
            .O(N__40763),
            .I(\phase_controller_slave.start_timer_hcZ0 ));
    Odrv4 I__9055 (
            .O(N__40760),
            .I(\phase_controller_slave.start_timer_hcZ0 ));
    Odrv4 I__9054 (
            .O(N__40755),
            .I(\phase_controller_slave.start_timer_hcZ0 ));
    Odrv4 I__9053 (
            .O(N__40752),
            .I(\phase_controller_slave.start_timer_hcZ0 ));
    InMux I__9052 (
            .O(N__40739),
            .I(N__40735));
    InMux I__9051 (
            .O(N__40738),
            .I(N__40732));
    LocalMux I__9050 (
            .O(N__40735),
            .I(N__40729));
    LocalMux I__9049 (
            .O(N__40732),
            .I(N__40725));
    Span4Mux_v I__9048 (
            .O(N__40729),
            .I(N__40722));
    InMux I__9047 (
            .O(N__40728),
            .I(N__40719));
    Span4Mux_h I__9046 (
            .O(N__40725),
            .I(N__40713));
    Span4Mux_h I__9045 (
            .O(N__40722),
            .I(N__40708));
    LocalMux I__9044 (
            .O(N__40719),
            .I(N__40708));
    InMux I__9043 (
            .O(N__40718),
            .I(N__40705));
    InMux I__9042 (
            .O(N__40717),
            .I(N__40700));
    InMux I__9041 (
            .O(N__40716),
            .I(N__40700));
    Odrv4 I__9040 (
            .O(N__40713),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__9039 (
            .O(N__40708),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__9038 (
            .O(N__40705),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__9037 (
            .O(N__40700),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    CascadeMux I__9036 (
            .O(N__40691),
            .I(N__40687));
    CascadeMux I__9035 (
            .O(N__40690),
            .I(N__40684));
    InMux I__9034 (
            .O(N__40687),
            .I(N__40674));
    InMux I__9033 (
            .O(N__40684),
            .I(N__40674));
    InMux I__9032 (
            .O(N__40683),
            .I(N__40671));
    InMux I__9031 (
            .O(N__40682),
            .I(N__40668));
    InMux I__9030 (
            .O(N__40681),
            .I(N__40656));
    InMux I__9029 (
            .O(N__40680),
            .I(N__40656));
    InMux I__9028 (
            .O(N__40679),
            .I(N__40656));
    LocalMux I__9027 (
            .O(N__40674),
            .I(N__40650));
    LocalMux I__9026 (
            .O(N__40671),
            .I(N__40650));
    LocalMux I__9025 (
            .O(N__40668),
            .I(N__40647));
    CascadeMux I__9024 (
            .O(N__40667),
            .I(N__40644));
    CascadeMux I__9023 (
            .O(N__40666),
            .I(N__40641));
    CascadeMux I__9022 (
            .O(N__40665),
            .I(N__40637));
    InMux I__9021 (
            .O(N__40664),
            .I(N__40625));
    InMux I__9020 (
            .O(N__40663),
            .I(N__40622));
    LocalMux I__9019 (
            .O(N__40656),
            .I(N__40619));
    InMux I__9018 (
            .O(N__40655),
            .I(N__40616));
    Span4Mux_v I__9017 (
            .O(N__40650),
            .I(N__40611));
    Span4Mux_v I__9016 (
            .O(N__40647),
            .I(N__40611));
    InMux I__9015 (
            .O(N__40644),
            .I(N__40604));
    InMux I__9014 (
            .O(N__40641),
            .I(N__40604));
    InMux I__9013 (
            .O(N__40640),
            .I(N__40604));
    InMux I__9012 (
            .O(N__40637),
            .I(N__40595));
    InMux I__9011 (
            .O(N__40636),
            .I(N__40595));
    InMux I__9010 (
            .O(N__40635),
            .I(N__40595));
    InMux I__9009 (
            .O(N__40634),
            .I(N__40595));
    InMux I__9008 (
            .O(N__40633),
            .I(N__40588));
    InMux I__9007 (
            .O(N__40632),
            .I(N__40588));
    InMux I__9006 (
            .O(N__40631),
            .I(N__40588));
    InMux I__9005 (
            .O(N__40630),
            .I(N__40583));
    InMux I__9004 (
            .O(N__40629),
            .I(N__40583));
    InMux I__9003 (
            .O(N__40628),
            .I(N__40580));
    LocalMux I__9002 (
            .O(N__40625),
            .I(N__40572));
    LocalMux I__9001 (
            .O(N__40622),
            .I(N__40572));
    Span4Mux_v I__9000 (
            .O(N__40619),
            .I(N__40572));
    LocalMux I__8999 (
            .O(N__40616),
            .I(N__40569));
    Span4Mux_v I__8998 (
            .O(N__40611),
            .I(N__40564));
    LocalMux I__8997 (
            .O(N__40604),
            .I(N__40564));
    LocalMux I__8996 (
            .O(N__40595),
            .I(N__40557));
    LocalMux I__8995 (
            .O(N__40588),
            .I(N__40557));
    LocalMux I__8994 (
            .O(N__40583),
            .I(N__40557));
    LocalMux I__8993 (
            .O(N__40580),
            .I(N__40554));
    InMux I__8992 (
            .O(N__40579),
            .I(N__40551));
    Span4Mux_v I__8991 (
            .O(N__40572),
            .I(N__40548));
    Span4Mux_h I__8990 (
            .O(N__40569),
            .I(N__40543));
    Span4Mux_h I__8989 (
            .O(N__40564),
            .I(N__40543));
    Span4Mux_v I__8988 (
            .O(N__40557),
            .I(N__40538));
    Span4Mux_h I__8987 (
            .O(N__40554),
            .I(N__40538));
    LocalMux I__8986 (
            .O(N__40551),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__8985 (
            .O(N__40548),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__8984 (
            .O(N__40543),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__8983 (
            .O(N__40538),
            .I(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ));
    IoInMux I__8982 (
            .O(N__40529),
            .I(N__40526));
    LocalMux I__8981 (
            .O(N__40526),
            .I(N__40523));
    Span4Mux_s2_v I__8980 (
            .O(N__40523),
            .I(N__40519));
    CEMux I__8979 (
            .O(N__40522),
            .I(N__40515));
    Span4Mux_h I__8978 (
            .O(N__40519),
            .I(N__40511));
    CEMux I__8977 (
            .O(N__40518),
            .I(N__40508));
    LocalMux I__8976 (
            .O(N__40515),
            .I(N__40505));
    CEMux I__8975 (
            .O(N__40514),
            .I(N__40502));
    Span4Mux_v I__8974 (
            .O(N__40511),
            .I(N__40499));
    LocalMux I__8973 (
            .O(N__40508),
            .I(N__40496));
    Span4Mux_v I__8972 (
            .O(N__40505),
            .I(N__40491));
    LocalMux I__8971 (
            .O(N__40502),
            .I(N__40491));
    Span4Mux_v I__8970 (
            .O(N__40499),
            .I(N__40488));
    Sp12to4 I__8969 (
            .O(N__40496),
            .I(N__40485));
    Span4Mux_v I__8968 (
            .O(N__40491),
            .I(N__40482));
    Odrv4 I__8967 (
            .O(N__40488),
            .I(red_c_i));
    Odrv12 I__8966 (
            .O(N__40485),
            .I(red_c_i));
    Odrv4 I__8965 (
            .O(N__40482),
            .I(red_c_i));
    CascadeMux I__8964 (
            .O(N__40475),
            .I(N__40472));
    InMux I__8963 (
            .O(N__40472),
            .I(N__40469));
    LocalMux I__8962 (
            .O(N__40469),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_17 ));
    CascadeMux I__8961 (
            .O(N__40466),
            .I(N__40463));
    InMux I__8960 (
            .O(N__40463),
            .I(N__40460));
    LocalMux I__8959 (
            .O(N__40460),
            .I(N__40457));
    Odrv4 I__8958 (
            .O(N__40457),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_8 ));
    InMux I__8957 (
            .O(N__40454),
            .I(N__40450));
    InMux I__8956 (
            .O(N__40453),
            .I(N__40447));
    LocalMux I__8955 (
            .O(N__40450),
            .I(N__40444));
    LocalMux I__8954 (
            .O(N__40447),
            .I(N__40441));
    Span4Mux_v I__8953 (
            .O(N__40444),
            .I(N__40436));
    Span4Mux_v I__8952 (
            .O(N__40441),
            .I(N__40433));
    InMux I__8951 (
            .O(N__40440),
            .I(N__40430));
    CascadeMux I__8950 (
            .O(N__40439),
            .I(N__40426));
    Span4Mux_v I__8949 (
            .O(N__40436),
            .I(N__40419));
    Span4Mux_h I__8948 (
            .O(N__40433),
            .I(N__40419));
    LocalMux I__8947 (
            .O(N__40430),
            .I(N__40419));
    InMux I__8946 (
            .O(N__40429),
            .I(N__40414));
    InMux I__8945 (
            .O(N__40426),
            .I(N__40414));
    Odrv4 I__8944 (
            .O(N__40419),
            .I(measured_delay_hc_16));
    LocalMux I__8943 (
            .O(N__40414),
            .I(measured_delay_hc_16));
    CascadeMux I__8942 (
            .O(N__40409),
            .I(N__40406));
    InMux I__8941 (
            .O(N__40406),
            .I(N__40403));
    LocalMux I__8940 (
            .O(N__40403),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_16 ));
    InMux I__8939 (
            .O(N__40400),
            .I(N__40397));
    LocalMux I__8938 (
            .O(N__40397),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_18 ));
    InMux I__8937 (
            .O(N__40394),
            .I(N__40390));
    InMux I__8936 (
            .O(N__40393),
            .I(N__40386));
    LocalMux I__8935 (
            .O(N__40390),
            .I(N__40383));
    InMux I__8934 (
            .O(N__40389),
            .I(N__40380));
    LocalMux I__8933 (
            .O(N__40386),
            .I(N__40377));
    Span4Mux_h I__8932 (
            .O(N__40383),
            .I(N__40374));
    LocalMux I__8931 (
            .O(N__40380),
            .I(N__40371));
    Span4Mux_h I__8930 (
            .O(N__40377),
            .I(N__40368));
    Span4Mux_v I__8929 (
            .O(N__40374),
            .I(N__40365));
    Span4Mux_h I__8928 (
            .O(N__40371),
            .I(N__40360));
    Span4Mux_v I__8927 (
            .O(N__40368),
            .I(N__40360));
    Odrv4 I__8926 (
            .O(N__40365),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1 ));
    Odrv4 I__8925 (
            .O(N__40360),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1 ));
    CascadeMux I__8924 (
            .O(N__40355),
            .I(N__40352));
    InMux I__8923 (
            .O(N__40352),
            .I(N__40349));
    LocalMux I__8922 (
            .O(N__40349),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_19 ));
    InMux I__8921 (
            .O(N__40346),
            .I(N__40337));
    InMux I__8920 (
            .O(N__40345),
            .I(N__40337));
    InMux I__8919 (
            .O(N__40344),
            .I(N__40332));
    CascadeMux I__8918 (
            .O(N__40343),
            .I(N__40329));
    InMux I__8917 (
            .O(N__40342),
            .I(N__40323));
    LocalMux I__8916 (
            .O(N__40337),
            .I(N__40320));
    InMux I__8915 (
            .O(N__40336),
            .I(N__40311));
    InMux I__8914 (
            .O(N__40335),
            .I(N__40311));
    LocalMux I__8913 (
            .O(N__40332),
            .I(N__40308));
    InMux I__8912 (
            .O(N__40329),
            .I(N__40299));
    InMux I__8911 (
            .O(N__40328),
            .I(N__40299));
    InMux I__8910 (
            .O(N__40327),
            .I(N__40299));
    InMux I__8909 (
            .O(N__40326),
            .I(N__40299));
    LocalMux I__8908 (
            .O(N__40323),
            .I(N__40296));
    Span4Mux_h I__8907 (
            .O(N__40320),
            .I(N__40293));
    InMux I__8906 (
            .O(N__40319),
            .I(N__40284));
    InMux I__8905 (
            .O(N__40318),
            .I(N__40284));
    InMux I__8904 (
            .O(N__40317),
            .I(N__40284));
    InMux I__8903 (
            .O(N__40316),
            .I(N__40284));
    LocalMux I__8902 (
            .O(N__40311),
            .I(N__40281));
    Span4Mux_v I__8901 (
            .O(N__40308),
            .I(N__40278));
    LocalMux I__8900 (
            .O(N__40299),
            .I(N__40275));
    Span4Mux_v I__8899 (
            .O(N__40296),
            .I(N__40272));
    Span4Mux_v I__8898 (
            .O(N__40293),
            .I(N__40269));
    LocalMux I__8897 (
            .O(N__40284),
            .I(N__40262));
    Span4Mux_v I__8896 (
            .O(N__40281),
            .I(N__40262));
    Span4Mux_v I__8895 (
            .O(N__40278),
            .I(N__40262));
    Span12Mux_h I__8894 (
            .O(N__40275),
            .I(N__40259));
    Odrv4 I__8893 (
            .O(N__40272),
            .I(\phase_controller_inst1.stoper_hc.un2_startlt31 ));
    Odrv4 I__8892 (
            .O(N__40269),
            .I(\phase_controller_inst1.stoper_hc.un2_startlt31 ));
    Odrv4 I__8891 (
            .O(N__40262),
            .I(\phase_controller_inst1.stoper_hc.un2_startlt31 ));
    Odrv12 I__8890 (
            .O(N__40259),
            .I(\phase_controller_inst1.stoper_hc.un2_startlt31 ));
    InMux I__8889 (
            .O(N__40250),
            .I(N__40245));
    InMux I__8888 (
            .O(N__40249),
            .I(N__40242));
    InMux I__8887 (
            .O(N__40248),
            .I(N__40239));
    LocalMux I__8886 (
            .O(N__40245),
            .I(N__40236));
    LocalMux I__8885 (
            .O(N__40242),
            .I(N__40233));
    LocalMux I__8884 (
            .O(N__40239),
            .I(N__40230));
    Span4Mux_v I__8883 (
            .O(N__40236),
            .I(N__40225));
    Span4Mux_h I__8882 (
            .O(N__40233),
            .I(N__40225));
    Span12Mux_v I__8881 (
            .O(N__40230),
            .I(N__40222));
    Odrv4 I__8880 (
            .O(N__40225),
            .I(measured_delay_tr_6));
    Odrv12 I__8879 (
            .O(N__40222),
            .I(measured_delay_tr_6));
    InMux I__8878 (
            .O(N__40217),
            .I(N__40210));
    InMux I__8877 (
            .O(N__40216),
            .I(N__40210));
    CascadeMux I__8876 (
            .O(N__40215),
            .I(N__40207));
    LocalMux I__8875 (
            .O(N__40210),
            .I(N__40202));
    InMux I__8874 (
            .O(N__40207),
            .I(N__40195));
    InMux I__8873 (
            .O(N__40206),
            .I(N__40195));
    InMux I__8872 (
            .O(N__40205),
            .I(N__40195));
    Span4Mux_v I__8871 (
            .O(N__40202),
            .I(N__40192));
    LocalMux I__8870 (
            .O(N__40195),
            .I(N__40189));
    Span4Mux_h I__8869 (
            .O(N__40192),
            .I(N__40186));
    Span4Mux_v I__8868 (
            .O(N__40189),
            .I(N__40183));
    Odrv4 I__8867 (
            .O(N__40186),
            .I(measured_delay_tr_3));
    Odrv4 I__8866 (
            .O(N__40183),
            .I(measured_delay_tr_3));
    InMux I__8865 (
            .O(N__40178),
            .I(N__40174));
    CascadeMux I__8864 (
            .O(N__40177),
            .I(N__40171));
    LocalMux I__8863 (
            .O(N__40174),
            .I(N__40168));
    InMux I__8862 (
            .O(N__40171),
            .I(N__40165));
    Span4Mux_v I__8861 (
            .O(N__40168),
            .I(N__40161));
    LocalMux I__8860 (
            .O(N__40165),
            .I(N__40158));
    InMux I__8859 (
            .O(N__40164),
            .I(N__40155));
    Span4Mux_h I__8858 (
            .O(N__40161),
            .I(N__40150));
    Span4Mux_v I__8857 (
            .O(N__40158),
            .I(N__40150));
    LocalMux I__8856 (
            .O(N__40155),
            .I(N__40147));
    Sp12to4 I__8855 (
            .O(N__40150),
            .I(N__40142));
    Span12Mux_h I__8854 (
            .O(N__40147),
            .I(N__40142));
    Odrv12 I__8853 (
            .O(N__40142),
            .I(measured_delay_tr_5));
    InMux I__8852 (
            .O(N__40139),
            .I(N__40135));
    InMux I__8851 (
            .O(N__40138),
            .I(N__40132));
    LocalMux I__8850 (
            .O(N__40135),
            .I(N__40129));
    LocalMux I__8849 (
            .O(N__40132),
            .I(N__40126));
    Odrv12 I__8848 (
            .O(N__40129),
            .I(\delay_measurement_inst.elapsed_time_tr_1 ));
    Odrv4 I__8847 (
            .O(N__40126),
            .I(\delay_measurement_inst.elapsed_time_tr_1 ));
    CascadeMux I__8846 (
            .O(N__40121),
            .I(N__40118));
    InMux I__8845 (
            .O(N__40118),
            .I(N__40114));
    InMux I__8844 (
            .O(N__40117),
            .I(N__40111));
    LocalMux I__8843 (
            .O(N__40114),
            .I(N__40108));
    LocalMux I__8842 (
            .O(N__40111),
            .I(N__40105));
    Span4Mux_v I__8841 (
            .O(N__40108),
            .I(N__40102));
    Span4Mux_v I__8840 (
            .O(N__40105),
            .I(N__40099));
    Odrv4 I__8839 (
            .O(N__40102),
            .I(measured_delay_tr_1));
    Odrv4 I__8838 (
            .O(N__40099),
            .I(measured_delay_tr_1));
    InMux I__8837 (
            .O(N__40094),
            .I(N__40089));
    InMux I__8836 (
            .O(N__40093),
            .I(N__40084));
    InMux I__8835 (
            .O(N__40092),
            .I(N__40084));
    LocalMux I__8834 (
            .O(N__40089),
            .I(N__40081));
    LocalMux I__8833 (
            .O(N__40084),
            .I(N__40078));
    Span4Mux_h I__8832 (
            .O(N__40081),
            .I(N__40075));
    Span4Mux_v I__8831 (
            .O(N__40078),
            .I(N__40072));
    Odrv4 I__8830 (
            .O(N__40075),
            .I(measured_delay_tr_2));
    Odrv4 I__8829 (
            .O(N__40072),
            .I(measured_delay_tr_2));
    InMux I__8828 (
            .O(N__40067),
            .I(N__40061));
    InMux I__8827 (
            .O(N__40066),
            .I(N__40056));
    InMux I__8826 (
            .O(N__40065),
            .I(N__40056));
    InMux I__8825 (
            .O(N__40064),
            .I(N__40053));
    LocalMux I__8824 (
            .O(N__40061),
            .I(N__40050));
    LocalMux I__8823 (
            .O(N__40056),
            .I(N__40047));
    LocalMux I__8822 (
            .O(N__40053),
            .I(N__40044));
    Span4Mux_h I__8821 (
            .O(N__40050),
            .I(N__40041));
    Span12Mux_h I__8820 (
            .O(N__40047),
            .I(N__40036));
    Span4Mux_h I__8819 (
            .O(N__40044),
            .I(N__40031));
    Span4Mux_v I__8818 (
            .O(N__40041),
            .I(N__40031));
    InMux I__8817 (
            .O(N__40040),
            .I(N__40026));
    InMux I__8816 (
            .O(N__40039),
            .I(N__40026));
    Odrv12 I__8815 (
            .O(N__40036),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__8814 (
            .O(N__40031),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__8813 (
            .O(N__40026),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    CascadeMux I__8812 (
            .O(N__40019),
            .I(N__40008));
    CascadeMux I__8811 (
            .O(N__40018),
            .I(N__40003));
    CascadeMux I__8810 (
            .O(N__40017),
            .I(N__39998));
    CascadeMux I__8809 (
            .O(N__40016),
            .I(N__39995));
    CascadeMux I__8808 (
            .O(N__40015),
            .I(N__39991));
    CascadeMux I__8807 (
            .O(N__40014),
            .I(N__39985));
    CascadeMux I__8806 (
            .O(N__40013),
            .I(N__39982));
    CascadeMux I__8805 (
            .O(N__40012),
            .I(N__39979));
    InMux I__8804 (
            .O(N__40011),
            .I(N__39972));
    InMux I__8803 (
            .O(N__40008),
            .I(N__39972));
    CascadeMux I__8802 (
            .O(N__40007),
            .I(N__39969));
    CascadeMux I__8801 (
            .O(N__40006),
            .I(N__39966));
    InMux I__8800 (
            .O(N__40003),
            .I(N__39963));
    InMux I__8799 (
            .O(N__40002),
            .I(N__39946));
    InMux I__8798 (
            .O(N__40001),
            .I(N__39946));
    InMux I__8797 (
            .O(N__39998),
            .I(N__39946));
    InMux I__8796 (
            .O(N__39995),
            .I(N__39946));
    InMux I__8795 (
            .O(N__39994),
            .I(N__39946));
    InMux I__8794 (
            .O(N__39991),
            .I(N__39946));
    InMux I__8793 (
            .O(N__39990),
            .I(N__39946));
    InMux I__8792 (
            .O(N__39989),
            .I(N__39933));
    InMux I__8791 (
            .O(N__39988),
            .I(N__39933));
    InMux I__8790 (
            .O(N__39985),
            .I(N__39933));
    InMux I__8789 (
            .O(N__39982),
            .I(N__39933));
    InMux I__8788 (
            .O(N__39979),
            .I(N__39933));
    InMux I__8787 (
            .O(N__39978),
            .I(N__39933));
    CascadeMux I__8786 (
            .O(N__39977),
            .I(N__39929));
    LocalMux I__8785 (
            .O(N__39972),
            .I(N__39925));
    InMux I__8784 (
            .O(N__39969),
            .I(N__39920));
    InMux I__8783 (
            .O(N__39966),
            .I(N__39920));
    LocalMux I__8782 (
            .O(N__39963),
            .I(N__39917));
    InMux I__8781 (
            .O(N__39962),
            .I(N__39914));
    InMux I__8780 (
            .O(N__39961),
            .I(N__39911));
    LocalMux I__8779 (
            .O(N__39946),
            .I(N__39907));
    LocalMux I__8778 (
            .O(N__39933),
            .I(N__39904));
    InMux I__8777 (
            .O(N__39932),
            .I(N__39899));
    InMux I__8776 (
            .O(N__39929),
            .I(N__39899));
    CascadeMux I__8775 (
            .O(N__39928),
            .I(N__39896));
    Span4Mux_v I__8774 (
            .O(N__39925),
            .I(N__39893));
    LocalMux I__8773 (
            .O(N__39920),
            .I(N__39890));
    Span4Mux_v I__8772 (
            .O(N__39917),
            .I(N__39883));
    LocalMux I__8771 (
            .O(N__39914),
            .I(N__39883));
    LocalMux I__8770 (
            .O(N__39911),
            .I(N__39883));
    InMux I__8769 (
            .O(N__39910),
            .I(N__39880));
    Span4Mux_v I__8768 (
            .O(N__39907),
            .I(N__39873));
    Span4Mux_v I__8767 (
            .O(N__39904),
            .I(N__39873));
    LocalMux I__8766 (
            .O(N__39899),
            .I(N__39873));
    InMux I__8765 (
            .O(N__39896),
            .I(N__39870));
    Span4Mux_h I__8764 (
            .O(N__39893),
            .I(N__39863));
    Span4Mux_h I__8763 (
            .O(N__39890),
            .I(N__39863));
    Span4Mux_h I__8762 (
            .O(N__39883),
            .I(N__39863));
    LocalMux I__8761 (
            .O(N__39880),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__8760 (
            .O(N__39873),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    LocalMux I__8759 (
            .O(N__39870),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__8758 (
            .O(N__39863),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    CascadeMux I__8757 (
            .O(N__39854),
            .I(N__39842));
    CascadeMux I__8756 (
            .O(N__39853),
            .I(N__39839));
    CascadeMux I__8755 (
            .O(N__39852),
            .I(N__39836));
    CascadeMux I__8754 (
            .O(N__39851),
            .I(N__39833));
    CascadeMux I__8753 (
            .O(N__39850),
            .I(N__39830));
    CascadeMux I__8752 (
            .O(N__39849),
            .I(N__39827));
    CascadeMux I__8751 (
            .O(N__39848),
            .I(N__39824));
    InMux I__8750 (
            .O(N__39847),
            .I(N__39813));
    InMux I__8749 (
            .O(N__39846),
            .I(N__39813));
    InMux I__8748 (
            .O(N__39845),
            .I(N__39808));
    InMux I__8747 (
            .O(N__39842),
            .I(N__39799));
    InMux I__8746 (
            .O(N__39839),
            .I(N__39799));
    InMux I__8745 (
            .O(N__39836),
            .I(N__39799));
    InMux I__8744 (
            .O(N__39833),
            .I(N__39799));
    InMux I__8743 (
            .O(N__39830),
            .I(N__39792));
    InMux I__8742 (
            .O(N__39827),
            .I(N__39792));
    InMux I__8741 (
            .O(N__39824),
            .I(N__39792));
    InMux I__8740 (
            .O(N__39823),
            .I(N__39785));
    InMux I__8739 (
            .O(N__39822),
            .I(N__39785));
    InMux I__8738 (
            .O(N__39821),
            .I(N__39785));
    InMux I__8737 (
            .O(N__39820),
            .I(N__39778));
    InMux I__8736 (
            .O(N__39819),
            .I(N__39778));
    InMux I__8735 (
            .O(N__39818),
            .I(N__39778));
    LocalMux I__8734 (
            .O(N__39813),
            .I(N__39775));
    InMux I__8733 (
            .O(N__39812),
            .I(N__39770));
    InMux I__8732 (
            .O(N__39811),
            .I(N__39770));
    LocalMux I__8731 (
            .O(N__39808),
            .I(N__39755));
    LocalMux I__8730 (
            .O(N__39799),
            .I(N__39755));
    LocalMux I__8729 (
            .O(N__39792),
            .I(N__39755));
    LocalMux I__8728 (
            .O(N__39785),
            .I(N__39755));
    LocalMux I__8727 (
            .O(N__39778),
            .I(N__39755));
    Span4Mux_v I__8726 (
            .O(N__39775),
            .I(N__39750));
    LocalMux I__8725 (
            .O(N__39770),
            .I(N__39750));
    InMux I__8724 (
            .O(N__39769),
            .I(N__39747));
    InMux I__8723 (
            .O(N__39768),
            .I(N__39744));
    InMux I__8722 (
            .O(N__39767),
            .I(N__39739));
    InMux I__8721 (
            .O(N__39766),
            .I(N__39739));
    Span4Mux_h I__8720 (
            .O(N__39755),
            .I(N__39735));
    Span4Mux_h I__8719 (
            .O(N__39750),
            .I(N__39732));
    LocalMux I__8718 (
            .O(N__39747),
            .I(N__39729));
    LocalMux I__8717 (
            .O(N__39744),
            .I(N__39726));
    LocalMux I__8716 (
            .O(N__39739),
            .I(N__39723));
    CascadeMux I__8715 (
            .O(N__39738),
            .I(N__39720));
    Span4Mux_v I__8714 (
            .O(N__39735),
            .I(N__39716));
    Span4Mux_v I__8713 (
            .O(N__39732),
            .I(N__39713));
    Span4Mux_h I__8712 (
            .O(N__39729),
            .I(N__39710));
    Span4Mux_v I__8711 (
            .O(N__39726),
            .I(N__39705));
    Span4Mux_h I__8710 (
            .O(N__39723),
            .I(N__39705));
    InMux I__8709 (
            .O(N__39720),
            .I(N__39700));
    InMux I__8708 (
            .O(N__39719),
            .I(N__39700));
    Span4Mux_h I__8707 (
            .O(N__39716),
            .I(N__39697));
    Span4Mux_h I__8706 (
            .O(N__39713),
            .I(N__39694));
    Span4Mux_h I__8705 (
            .O(N__39710),
            .I(N__39689));
    Span4Mux_h I__8704 (
            .O(N__39705),
            .I(N__39689));
    LocalMux I__8703 (
            .O(N__39700),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__8702 (
            .O(N__39697),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__8701 (
            .O(N__39694),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__8700 (
            .O(N__39689),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    CascadeMux I__8699 (
            .O(N__39680),
            .I(N__39675));
    InMux I__8698 (
            .O(N__39679),
            .I(N__39670));
    InMux I__8697 (
            .O(N__39678),
            .I(N__39670));
    InMux I__8696 (
            .O(N__39675),
            .I(N__39651));
    LocalMux I__8695 (
            .O(N__39670),
            .I(N__39648));
    InMux I__8694 (
            .O(N__39669),
            .I(N__39645));
    InMux I__8693 (
            .O(N__39668),
            .I(N__39642));
    InMux I__8692 (
            .O(N__39667),
            .I(N__39629));
    InMux I__8691 (
            .O(N__39666),
            .I(N__39629));
    InMux I__8690 (
            .O(N__39665),
            .I(N__39629));
    InMux I__8689 (
            .O(N__39664),
            .I(N__39629));
    InMux I__8688 (
            .O(N__39663),
            .I(N__39629));
    InMux I__8687 (
            .O(N__39662),
            .I(N__39629));
    InMux I__8686 (
            .O(N__39661),
            .I(N__39614));
    InMux I__8685 (
            .O(N__39660),
            .I(N__39614));
    InMux I__8684 (
            .O(N__39659),
            .I(N__39614));
    InMux I__8683 (
            .O(N__39658),
            .I(N__39614));
    InMux I__8682 (
            .O(N__39657),
            .I(N__39614));
    InMux I__8681 (
            .O(N__39656),
            .I(N__39614));
    InMux I__8680 (
            .O(N__39655),
            .I(N__39614));
    InMux I__8679 (
            .O(N__39654),
            .I(N__39611));
    LocalMux I__8678 (
            .O(N__39651),
            .I(N__39601));
    Span4Mux_v I__8677 (
            .O(N__39648),
            .I(N__39601));
    LocalMux I__8676 (
            .O(N__39645),
            .I(N__39601));
    LocalMux I__8675 (
            .O(N__39642),
            .I(N__39594));
    LocalMux I__8674 (
            .O(N__39629),
            .I(N__39594));
    LocalMux I__8673 (
            .O(N__39614),
            .I(N__39594));
    LocalMux I__8672 (
            .O(N__39611),
            .I(N__39591));
    InMux I__8671 (
            .O(N__39610),
            .I(N__39588));
    InMux I__8670 (
            .O(N__39609),
            .I(N__39583));
    InMux I__8669 (
            .O(N__39608),
            .I(N__39583));
    Span4Mux_h I__8668 (
            .O(N__39601),
            .I(N__39580));
    Span4Mux_h I__8667 (
            .O(N__39594),
            .I(N__39577));
    Span4Mux_v I__8666 (
            .O(N__39591),
            .I(N__39570));
    LocalMux I__8665 (
            .O(N__39588),
            .I(N__39570));
    LocalMux I__8664 (
            .O(N__39583),
            .I(N__39570));
    Span4Mux_v I__8663 (
            .O(N__39580),
            .I(N__39565));
    Span4Mux_v I__8662 (
            .O(N__39577),
            .I(N__39562));
    Span4Mux_h I__8661 (
            .O(N__39570),
            .I(N__39559));
    InMux I__8660 (
            .O(N__39569),
            .I(N__39554));
    InMux I__8659 (
            .O(N__39568),
            .I(N__39554));
    Span4Mux_h I__8658 (
            .O(N__39565),
            .I(N__39551));
    Span4Mux_h I__8657 (
            .O(N__39562),
            .I(N__39548));
    Span4Mux_h I__8656 (
            .O(N__39559),
            .I(N__39545));
    LocalMux I__8655 (
            .O(N__39554),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__8654 (
            .O(N__39551),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__8653 (
            .O(N__39548),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__8652 (
            .O(N__39545),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    InMux I__8651 (
            .O(N__39536),
            .I(N__39532));
    InMux I__8650 (
            .O(N__39535),
            .I(N__39529));
    LocalMux I__8649 (
            .O(N__39532),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10 ));
    LocalMux I__8648 (
            .O(N__39529),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10 ));
    CascadeMux I__8647 (
            .O(N__39524),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10_cascade_ ));
    CascadeMux I__8646 (
            .O(N__39521),
            .I(\delay_measurement_inst.delay_tr_timer.N_400_cascade_ ));
    CascadeMux I__8645 (
            .O(N__39518),
            .I(\delay_measurement_inst.N_394_1_cascade_ ));
    InMux I__8644 (
            .O(N__39515),
            .I(N__39503));
    InMux I__8643 (
            .O(N__39514),
            .I(N__39503));
    InMux I__8642 (
            .O(N__39513),
            .I(N__39503));
    InMux I__8641 (
            .O(N__39512),
            .I(N__39503));
    LocalMux I__8640 (
            .O(N__39503),
            .I(\delay_measurement_inst.N_394_1 ));
    InMux I__8639 (
            .O(N__39500),
            .I(N__39497));
    LocalMux I__8638 (
            .O(N__39497),
            .I(N__39493));
    InMux I__8637 (
            .O(N__39496),
            .I(N__39490));
    Span4Mux_v I__8636 (
            .O(N__39493),
            .I(N__39486));
    LocalMux I__8635 (
            .O(N__39490),
            .I(N__39483));
    InMux I__8634 (
            .O(N__39489),
            .I(N__39480));
    Odrv4 I__8633 (
            .O(N__39486),
            .I(measured_delay_tr_12));
    Odrv4 I__8632 (
            .O(N__39483),
            .I(measured_delay_tr_12));
    LocalMux I__8631 (
            .O(N__39480),
            .I(measured_delay_tr_12));
    InMux I__8630 (
            .O(N__39473),
            .I(N__39470));
    LocalMux I__8629 (
            .O(N__39470),
            .I(N__39466));
    InMux I__8628 (
            .O(N__39469),
            .I(N__39463));
    Span4Mux_h I__8627 (
            .O(N__39466),
            .I(N__39459));
    LocalMux I__8626 (
            .O(N__39463),
            .I(N__39456));
    InMux I__8625 (
            .O(N__39462),
            .I(N__39453));
    Odrv4 I__8624 (
            .O(N__39459),
            .I(measured_delay_tr_10));
    Odrv4 I__8623 (
            .O(N__39456),
            .I(measured_delay_tr_10));
    LocalMux I__8622 (
            .O(N__39453),
            .I(measured_delay_tr_10));
    InMux I__8621 (
            .O(N__39446),
            .I(N__39443));
    LocalMux I__8620 (
            .O(N__39443),
            .I(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_4 ));
    CascadeMux I__8619 (
            .O(N__39440),
            .I(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_6_cascade_ ));
    InMux I__8618 (
            .O(N__39437),
            .I(N__39434));
    LocalMux I__8617 (
            .O(N__39434),
            .I(\delay_measurement_inst.delay_tr_timer.N_364 ));
    InMux I__8616 (
            .O(N__39431),
            .I(N__39428));
    LocalMux I__8615 (
            .O(N__39428),
            .I(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_5 ));
    CascadeMux I__8614 (
            .O(N__39425),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_6_19_cascade_ ));
    InMux I__8613 (
            .O(N__39422),
            .I(N__39419));
    LocalMux I__8612 (
            .O(N__39419),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_0_19 ));
    CascadeMux I__8611 (
            .O(N__39416),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20_cascade_ ));
    InMux I__8610 (
            .O(N__39413),
            .I(N__39410));
    LocalMux I__8609 (
            .O(N__39410),
            .I(\delay_measurement_inst.delay_tr_timer.N_409 ));
    InMux I__8608 (
            .O(N__39407),
            .I(N__39402));
    InMux I__8607 (
            .O(N__39406),
            .I(N__39398));
    CascadeMux I__8606 (
            .O(N__39405),
            .I(N__39395));
    LocalMux I__8605 (
            .O(N__39402),
            .I(N__39392));
    InMux I__8604 (
            .O(N__39401),
            .I(N__39389));
    LocalMux I__8603 (
            .O(N__39398),
            .I(N__39386));
    InMux I__8602 (
            .O(N__39395),
            .I(N__39383));
    Span4Mux_v I__8601 (
            .O(N__39392),
            .I(N__39380));
    LocalMux I__8600 (
            .O(N__39389),
            .I(N__39376));
    Span4Mux_v I__8599 (
            .O(N__39386),
            .I(N__39373));
    LocalMux I__8598 (
            .O(N__39383),
            .I(N__39368));
    Span4Mux_h I__8597 (
            .O(N__39380),
            .I(N__39368));
    InMux I__8596 (
            .O(N__39379),
            .I(N__39365));
    Span4Mux_v I__8595 (
            .O(N__39376),
            .I(N__39362));
    Odrv4 I__8594 (
            .O(N__39373),
            .I(measured_delay_hc_12));
    Odrv4 I__8593 (
            .O(N__39368),
            .I(measured_delay_hc_12));
    LocalMux I__8592 (
            .O(N__39365),
            .I(measured_delay_hc_12));
    Odrv4 I__8591 (
            .O(N__39362),
            .I(measured_delay_hc_12));
    InMux I__8590 (
            .O(N__39353),
            .I(N__39347));
    InMux I__8589 (
            .O(N__39352),
            .I(N__39344));
    InMux I__8588 (
            .O(N__39351),
            .I(N__39341));
    CascadeMux I__8587 (
            .O(N__39350),
            .I(N__39338));
    LocalMux I__8586 (
            .O(N__39347),
            .I(N__39335));
    LocalMux I__8585 (
            .O(N__39344),
            .I(N__39332));
    LocalMux I__8584 (
            .O(N__39341),
            .I(N__39328));
    InMux I__8583 (
            .O(N__39338),
            .I(N__39325));
    Span4Mux_v I__8582 (
            .O(N__39335),
            .I(N__39322));
    Span4Mux_h I__8581 (
            .O(N__39332),
            .I(N__39319));
    InMux I__8580 (
            .O(N__39331),
            .I(N__39316));
    Span4Mux_v I__8579 (
            .O(N__39328),
            .I(N__39313));
    LocalMux I__8578 (
            .O(N__39325),
            .I(measured_delay_hc_11));
    Odrv4 I__8577 (
            .O(N__39322),
            .I(measured_delay_hc_11));
    Odrv4 I__8576 (
            .O(N__39319),
            .I(measured_delay_hc_11));
    LocalMux I__8575 (
            .O(N__39316),
            .I(measured_delay_hc_11));
    Odrv4 I__8574 (
            .O(N__39313),
            .I(measured_delay_hc_11));
    InMux I__8573 (
            .O(N__39302),
            .I(N__39299));
    LocalMux I__8572 (
            .O(N__39299),
            .I(N__39296));
    Odrv4 I__8571 (
            .O(N__39296),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9 ));
    InMux I__8570 (
            .O(N__39293),
            .I(N__39290));
    LocalMux I__8569 (
            .O(N__39290),
            .I(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_5 ));
    CascadeMux I__8568 (
            .O(N__39287),
            .I(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_6_cascade_ ));
    InMux I__8567 (
            .O(N__39284),
            .I(N__39281));
    LocalMux I__8566 (
            .O(N__39281),
            .I(N__39278));
    Span4Mux_h I__8565 (
            .O(N__39278),
            .I(N__39275));
    Odrv4 I__8564 (
            .O(N__39275),
            .I(\delay_measurement_inst.tr_state_RNIMR6LZ0Z_0 ));
    CascadeMux I__8563 (
            .O(N__39272),
            .I(\delay_measurement_inst.delay_tr_timer.N_375_cascade_ ));
    CascadeMux I__8562 (
            .O(N__39269),
            .I(\delay_measurement_inst.N_265_i_cascade_ ));
    InMux I__8561 (
            .O(N__39266),
            .I(N__39263));
    LocalMux I__8560 (
            .O(N__39263),
            .I(N__39260));
    Span4Mux_v I__8559 (
            .O(N__39260),
            .I(N__39256));
    InMux I__8558 (
            .O(N__39259),
            .I(N__39251));
    Span4Mux_v I__8557 (
            .O(N__39256),
            .I(N__39248));
    InMux I__8556 (
            .O(N__39255),
            .I(N__39243));
    InMux I__8555 (
            .O(N__39254),
            .I(N__39243));
    LocalMux I__8554 (
            .O(N__39251),
            .I(N__39240));
    Odrv4 I__8553 (
            .O(N__39248),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    LocalMux I__8552 (
            .O(N__39243),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    Odrv4 I__8551 (
            .O(N__39240),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    CascadeMux I__8550 (
            .O(N__39233),
            .I(N__39228));
    CascadeMux I__8549 (
            .O(N__39232),
            .I(N__39225));
    InMux I__8548 (
            .O(N__39231),
            .I(N__39222));
    InMux I__8547 (
            .O(N__39228),
            .I(N__39217));
    InMux I__8546 (
            .O(N__39225),
            .I(N__39217));
    LocalMux I__8545 (
            .O(N__39222),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    LocalMux I__8544 (
            .O(N__39217),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    InMux I__8543 (
            .O(N__39212),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ));
    CascadeMux I__8542 (
            .O(N__39209),
            .I(N__39204));
    CascadeMux I__8541 (
            .O(N__39208),
            .I(N__39201));
    InMux I__8540 (
            .O(N__39207),
            .I(N__39198));
    InMux I__8539 (
            .O(N__39204),
            .I(N__39193));
    InMux I__8538 (
            .O(N__39201),
            .I(N__39193));
    LocalMux I__8537 (
            .O(N__39198),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    LocalMux I__8536 (
            .O(N__39193),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    InMux I__8535 (
            .O(N__39188),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ));
    InMux I__8534 (
            .O(N__39185),
            .I(N__39180));
    InMux I__8533 (
            .O(N__39184),
            .I(N__39177));
    InMux I__8532 (
            .O(N__39183),
            .I(N__39174));
    LocalMux I__8531 (
            .O(N__39180),
            .I(N__39171));
    LocalMux I__8530 (
            .O(N__39177),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    LocalMux I__8529 (
            .O(N__39174),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    Odrv4 I__8528 (
            .O(N__39171),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    InMux I__8527 (
            .O(N__39164),
            .I(bfn_16_10_0_));
    InMux I__8526 (
            .O(N__39161),
            .I(N__39156));
    InMux I__8525 (
            .O(N__39160),
            .I(N__39153));
    InMux I__8524 (
            .O(N__39159),
            .I(N__39150));
    LocalMux I__8523 (
            .O(N__39156),
            .I(N__39147));
    LocalMux I__8522 (
            .O(N__39153),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    LocalMux I__8521 (
            .O(N__39150),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    Odrv4 I__8520 (
            .O(N__39147),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    InMux I__8519 (
            .O(N__39140),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ));
    CascadeMux I__8518 (
            .O(N__39137),
            .I(N__39132));
    CascadeMux I__8517 (
            .O(N__39136),
            .I(N__39129));
    InMux I__8516 (
            .O(N__39135),
            .I(N__39126));
    InMux I__8515 (
            .O(N__39132),
            .I(N__39121));
    InMux I__8514 (
            .O(N__39129),
            .I(N__39121));
    LocalMux I__8513 (
            .O(N__39126),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    LocalMux I__8512 (
            .O(N__39121),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    InMux I__8511 (
            .O(N__39116),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ));
    CascadeMux I__8510 (
            .O(N__39113),
            .I(N__39108));
    CascadeMux I__8509 (
            .O(N__39112),
            .I(N__39105));
    InMux I__8508 (
            .O(N__39111),
            .I(N__39102));
    InMux I__8507 (
            .O(N__39108),
            .I(N__39097));
    InMux I__8506 (
            .O(N__39105),
            .I(N__39097));
    LocalMux I__8505 (
            .O(N__39102),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    LocalMux I__8504 (
            .O(N__39097),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    InMux I__8503 (
            .O(N__39092),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ));
    InMux I__8502 (
            .O(N__39089),
            .I(N__39085));
    InMux I__8501 (
            .O(N__39088),
            .I(N__39082));
    LocalMux I__8500 (
            .O(N__39085),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    LocalMux I__8499 (
            .O(N__39082),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    InMux I__8498 (
            .O(N__39077),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ));
    InMux I__8497 (
            .O(N__39074),
            .I(N__39044));
    InMux I__8496 (
            .O(N__39073),
            .I(N__39044));
    InMux I__8495 (
            .O(N__39072),
            .I(N__39035));
    InMux I__8494 (
            .O(N__39071),
            .I(N__39035));
    InMux I__8493 (
            .O(N__39070),
            .I(N__39035));
    InMux I__8492 (
            .O(N__39069),
            .I(N__39035));
    InMux I__8491 (
            .O(N__39068),
            .I(N__39022));
    InMux I__8490 (
            .O(N__39067),
            .I(N__39022));
    InMux I__8489 (
            .O(N__39066),
            .I(N__39022));
    InMux I__8488 (
            .O(N__39065),
            .I(N__39022));
    InMux I__8487 (
            .O(N__39064),
            .I(N__39013));
    InMux I__8486 (
            .O(N__39063),
            .I(N__39013));
    InMux I__8485 (
            .O(N__39062),
            .I(N__39013));
    InMux I__8484 (
            .O(N__39061),
            .I(N__39013));
    InMux I__8483 (
            .O(N__39060),
            .I(N__39004));
    InMux I__8482 (
            .O(N__39059),
            .I(N__39004));
    InMux I__8481 (
            .O(N__39058),
            .I(N__39004));
    InMux I__8480 (
            .O(N__39057),
            .I(N__39004));
    InMux I__8479 (
            .O(N__39056),
            .I(N__38995));
    InMux I__8478 (
            .O(N__39055),
            .I(N__38995));
    InMux I__8477 (
            .O(N__39054),
            .I(N__38995));
    InMux I__8476 (
            .O(N__39053),
            .I(N__38995));
    InMux I__8475 (
            .O(N__39052),
            .I(N__38986));
    InMux I__8474 (
            .O(N__39051),
            .I(N__38986));
    InMux I__8473 (
            .O(N__39050),
            .I(N__38986));
    InMux I__8472 (
            .O(N__39049),
            .I(N__38986));
    LocalMux I__8471 (
            .O(N__39044),
            .I(N__38983));
    LocalMux I__8470 (
            .O(N__39035),
            .I(N__38980));
    InMux I__8469 (
            .O(N__39034),
            .I(N__38971));
    InMux I__8468 (
            .O(N__39033),
            .I(N__38971));
    InMux I__8467 (
            .O(N__39032),
            .I(N__38971));
    InMux I__8466 (
            .O(N__39031),
            .I(N__38971));
    LocalMux I__8465 (
            .O(N__39022),
            .I(N__38962));
    LocalMux I__8464 (
            .O(N__39013),
            .I(N__38962));
    LocalMux I__8463 (
            .O(N__39004),
            .I(N__38962));
    LocalMux I__8462 (
            .O(N__38995),
            .I(N__38962));
    LocalMux I__8461 (
            .O(N__38986),
            .I(N__38959));
    Span4Mux_h I__8460 (
            .O(N__38983),
            .I(N__38956));
    Span4Mux_h I__8459 (
            .O(N__38980),
            .I(N__38953));
    LocalMux I__8458 (
            .O(N__38971),
            .I(N__38948));
    Span4Mux_v I__8457 (
            .O(N__38962),
            .I(N__38948));
    Odrv12 I__8456 (
            .O(N__38959),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__8455 (
            .O(N__38956),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__8454 (
            .O(N__38953),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__8453 (
            .O(N__38948),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    InMux I__8452 (
            .O(N__38939),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ));
    InMux I__8451 (
            .O(N__38936),
            .I(N__38932));
    InMux I__8450 (
            .O(N__38935),
            .I(N__38929));
    LocalMux I__8449 (
            .O(N__38932),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    LocalMux I__8448 (
            .O(N__38929),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    CEMux I__8447 (
            .O(N__38924),
            .I(N__38921));
    LocalMux I__8446 (
            .O(N__38921),
            .I(N__38918));
    Span4Mux_v I__8445 (
            .O(N__38918),
            .I(N__38913));
    CEMux I__8444 (
            .O(N__38917),
            .I(N__38910));
    CEMux I__8443 (
            .O(N__38916),
            .I(N__38906));
    Span4Mux_h I__8442 (
            .O(N__38913),
            .I(N__38901));
    LocalMux I__8441 (
            .O(N__38910),
            .I(N__38901));
    CEMux I__8440 (
            .O(N__38909),
            .I(N__38898));
    LocalMux I__8439 (
            .O(N__38906),
            .I(N__38895));
    Span4Mux_v I__8438 (
            .O(N__38901),
            .I(N__38890));
    LocalMux I__8437 (
            .O(N__38898),
            .I(N__38890));
    Span4Mux_h I__8436 (
            .O(N__38895),
            .I(N__38887));
    Span4Mux_v I__8435 (
            .O(N__38890),
            .I(N__38884));
    Odrv4 I__8434 (
            .O(N__38887),
            .I(\delay_measurement_inst.delay_hc_timer.N_322_i ));
    Odrv4 I__8433 (
            .O(N__38884),
            .I(\delay_measurement_inst.delay_hc_timer.N_322_i ));
    CascadeMux I__8432 (
            .O(N__38879),
            .I(N__38874));
    CascadeMux I__8431 (
            .O(N__38878),
            .I(N__38871));
    InMux I__8430 (
            .O(N__38877),
            .I(N__38868));
    InMux I__8429 (
            .O(N__38874),
            .I(N__38863));
    InMux I__8428 (
            .O(N__38871),
            .I(N__38863));
    LocalMux I__8427 (
            .O(N__38868),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    LocalMux I__8426 (
            .O(N__38863),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    InMux I__8425 (
            .O(N__38858),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ));
    CascadeMux I__8424 (
            .O(N__38855),
            .I(N__38850));
    CascadeMux I__8423 (
            .O(N__38854),
            .I(N__38847));
    InMux I__8422 (
            .O(N__38853),
            .I(N__38844));
    InMux I__8421 (
            .O(N__38850),
            .I(N__38839));
    InMux I__8420 (
            .O(N__38847),
            .I(N__38839));
    LocalMux I__8419 (
            .O(N__38844),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    LocalMux I__8418 (
            .O(N__38839),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    InMux I__8417 (
            .O(N__38834),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ));
    InMux I__8416 (
            .O(N__38831),
            .I(N__38826));
    InMux I__8415 (
            .O(N__38830),
            .I(N__38823));
    InMux I__8414 (
            .O(N__38829),
            .I(N__38820));
    LocalMux I__8413 (
            .O(N__38826),
            .I(N__38817));
    LocalMux I__8412 (
            .O(N__38823),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    LocalMux I__8411 (
            .O(N__38820),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    Odrv4 I__8410 (
            .O(N__38817),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    InMux I__8409 (
            .O(N__38810),
            .I(bfn_16_9_0_));
    InMux I__8408 (
            .O(N__38807),
            .I(N__38802));
    InMux I__8407 (
            .O(N__38806),
            .I(N__38799));
    InMux I__8406 (
            .O(N__38805),
            .I(N__38796));
    LocalMux I__8405 (
            .O(N__38802),
            .I(N__38793));
    LocalMux I__8404 (
            .O(N__38799),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    LocalMux I__8403 (
            .O(N__38796),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    Odrv4 I__8402 (
            .O(N__38793),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    InMux I__8401 (
            .O(N__38786),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ));
    CascadeMux I__8400 (
            .O(N__38783),
            .I(N__38778));
    CascadeMux I__8399 (
            .O(N__38782),
            .I(N__38775));
    InMux I__8398 (
            .O(N__38781),
            .I(N__38772));
    InMux I__8397 (
            .O(N__38778),
            .I(N__38767));
    InMux I__8396 (
            .O(N__38775),
            .I(N__38767));
    LocalMux I__8395 (
            .O(N__38772),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    LocalMux I__8394 (
            .O(N__38767),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    InMux I__8393 (
            .O(N__38762),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ));
    CascadeMux I__8392 (
            .O(N__38759),
            .I(N__38754));
    CascadeMux I__8391 (
            .O(N__38758),
            .I(N__38751));
    InMux I__8390 (
            .O(N__38757),
            .I(N__38748));
    InMux I__8389 (
            .O(N__38754),
            .I(N__38743));
    InMux I__8388 (
            .O(N__38751),
            .I(N__38743));
    LocalMux I__8387 (
            .O(N__38748),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    LocalMux I__8386 (
            .O(N__38743),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    InMux I__8385 (
            .O(N__38738),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ));
    InMux I__8384 (
            .O(N__38735),
            .I(N__38730));
    InMux I__8383 (
            .O(N__38734),
            .I(N__38725));
    InMux I__8382 (
            .O(N__38733),
            .I(N__38725));
    LocalMux I__8381 (
            .O(N__38730),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    LocalMux I__8380 (
            .O(N__38725),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    InMux I__8379 (
            .O(N__38720),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ));
    InMux I__8378 (
            .O(N__38717),
            .I(N__38712));
    InMux I__8377 (
            .O(N__38716),
            .I(N__38707));
    InMux I__8376 (
            .O(N__38715),
            .I(N__38707));
    LocalMux I__8375 (
            .O(N__38712),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    LocalMux I__8374 (
            .O(N__38707),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    InMux I__8373 (
            .O(N__38702),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ));
    CascadeMux I__8372 (
            .O(N__38699),
            .I(N__38694));
    CascadeMux I__8371 (
            .O(N__38698),
            .I(N__38691));
    InMux I__8370 (
            .O(N__38697),
            .I(N__38688));
    InMux I__8369 (
            .O(N__38694),
            .I(N__38683));
    InMux I__8368 (
            .O(N__38691),
            .I(N__38683));
    LocalMux I__8367 (
            .O(N__38688),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    LocalMux I__8366 (
            .O(N__38683),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    InMux I__8365 (
            .O(N__38678),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ));
    CascadeMux I__8364 (
            .O(N__38675),
            .I(N__38670));
    CascadeMux I__8363 (
            .O(N__38674),
            .I(N__38667));
    InMux I__8362 (
            .O(N__38673),
            .I(N__38664));
    InMux I__8361 (
            .O(N__38670),
            .I(N__38659));
    InMux I__8360 (
            .O(N__38667),
            .I(N__38659));
    LocalMux I__8359 (
            .O(N__38664),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    LocalMux I__8358 (
            .O(N__38659),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    InMux I__8357 (
            .O(N__38654),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ));
    InMux I__8356 (
            .O(N__38651),
            .I(N__38646));
    InMux I__8355 (
            .O(N__38650),
            .I(N__38643));
    InMux I__8354 (
            .O(N__38649),
            .I(N__38640));
    LocalMux I__8353 (
            .O(N__38646),
            .I(N__38637));
    LocalMux I__8352 (
            .O(N__38643),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    LocalMux I__8351 (
            .O(N__38640),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    Odrv4 I__8350 (
            .O(N__38637),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    InMux I__8349 (
            .O(N__38630),
            .I(bfn_16_8_0_));
    InMux I__8348 (
            .O(N__38627),
            .I(N__38622));
    InMux I__8347 (
            .O(N__38626),
            .I(N__38619));
    InMux I__8346 (
            .O(N__38625),
            .I(N__38616));
    LocalMux I__8345 (
            .O(N__38622),
            .I(N__38613));
    LocalMux I__8344 (
            .O(N__38619),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    LocalMux I__8343 (
            .O(N__38616),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    Odrv4 I__8342 (
            .O(N__38613),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    InMux I__8341 (
            .O(N__38606),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ));
    CascadeMux I__8340 (
            .O(N__38603),
            .I(N__38598));
    CascadeMux I__8339 (
            .O(N__38602),
            .I(N__38595));
    InMux I__8338 (
            .O(N__38601),
            .I(N__38592));
    InMux I__8337 (
            .O(N__38598),
            .I(N__38587));
    InMux I__8336 (
            .O(N__38595),
            .I(N__38587));
    LocalMux I__8335 (
            .O(N__38592),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    LocalMux I__8334 (
            .O(N__38587),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    InMux I__8333 (
            .O(N__38582),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ));
    CascadeMux I__8332 (
            .O(N__38579),
            .I(N__38574));
    CascadeMux I__8331 (
            .O(N__38578),
            .I(N__38571));
    InMux I__8330 (
            .O(N__38577),
            .I(N__38568));
    InMux I__8329 (
            .O(N__38574),
            .I(N__38563));
    InMux I__8328 (
            .O(N__38571),
            .I(N__38563));
    LocalMux I__8327 (
            .O(N__38568),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    LocalMux I__8326 (
            .O(N__38563),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    InMux I__8325 (
            .O(N__38558),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ));
    InMux I__8324 (
            .O(N__38555),
            .I(N__38550));
    InMux I__8323 (
            .O(N__38554),
            .I(N__38545));
    InMux I__8322 (
            .O(N__38553),
            .I(N__38545));
    LocalMux I__8321 (
            .O(N__38550),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    LocalMux I__8320 (
            .O(N__38545),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    InMux I__8319 (
            .O(N__38540),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ));
    InMux I__8318 (
            .O(N__38537),
            .I(N__38532));
    InMux I__8317 (
            .O(N__38536),
            .I(N__38527));
    InMux I__8316 (
            .O(N__38535),
            .I(N__38527));
    LocalMux I__8315 (
            .O(N__38532),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    LocalMux I__8314 (
            .O(N__38527),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    InMux I__8313 (
            .O(N__38522),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ));
    InMux I__8312 (
            .O(N__38519),
            .I(N__38516));
    LocalMux I__8311 (
            .O(N__38516),
            .I(N__38513));
    Odrv4 I__8310 (
            .O(N__38513),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9 ));
    InMux I__8309 (
            .O(N__38510),
            .I(N__38506));
    InMux I__8308 (
            .O(N__38509),
            .I(N__38503));
    LocalMux I__8307 (
            .O(N__38506),
            .I(N__38500));
    LocalMux I__8306 (
            .O(N__38503),
            .I(N__38497));
    Span4Mux_v I__8305 (
            .O(N__38500),
            .I(N__38494));
    Odrv4 I__8304 (
            .O(N__38497),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9 ));
    Odrv4 I__8303 (
            .O(N__38494),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9 ));
    CascadeMux I__8302 (
            .O(N__38489),
            .I(N__38486));
    InMux I__8301 (
            .O(N__38486),
            .I(N__38483));
    LocalMux I__8300 (
            .O(N__38483),
            .I(N__38480));
    Odrv12 I__8299 (
            .O(N__38480),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15 ));
    InMux I__8298 (
            .O(N__38477),
            .I(N__38473));
    InMux I__8297 (
            .O(N__38476),
            .I(N__38470));
    LocalMux I__8296 (
            .O(N__38473),
            .I(N__38467));
    LocalMux I__8295 (
            .O(N__38470),
            .I(N__38464));
    Span4Mux_v I__8294 (
            .O(N__38467),
            .I(N__38461));
    Odrv12 I__8293 (
            .O(N__38464),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15 ));
    Odrv4 I__8292 (
            .O(N__38461),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__8291 (
            .O(N__38456),
            .I(N__38451));
    InMux I__8290 (
            .O(N__38455),
            .I(N__38448));
    InMux I__8289 (
            .O(N__38454),
            .I(N__38445));
    LocalMux I__8288 (
            .O(N__38451),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__8287 (
            .O(N__38448),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__8286 (
            .O(N__38445),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    InMux I__8285 (
            .O(N__38438),
            .I(bfn_16_7_0_));
    InMux I__8284 (
            .O(N__38435),
            .I(N__38430));
    InMux I__8283 (
            .O(N__38434),
            .I(N__38427));
    InMux I__8282 (
            .O(N__38433),
            .I(N__38424));
    LocalMux I__8281 (
            .O(N__38430),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    LocalMux I__8280 (
            .O(N__38427),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    LocalMux I__8279 (
            .O(N__38424),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    InMux I__8278 (
            .O(N__38417),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ));
    CascadeMux I__8277 (
            .O(N__38414),
            .I(N__38409));
    CascadeMux I__8276 (
            .O(N__38413),
            .I(N__38406));
    InMux I__8275 (
            .O(N__38412),
            .I(N__38403));
    InMux I__8274 (
            .O(N__38409),
            .I(N__38398));
    InMux I__8273 (
            .O(N__38406),
            .I(N__38398));
    LocalMux I__8272 (
            .O(N__38403),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    LocalMux I__8271 (
            .O(N__38398),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    InMux I__8270 (
            .O(N__38393),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ));
    CascadeMux I__8269 (
            .O(N__38390),
            .I(N__38385));
    CascadeMux I__8268 (
            .O(N__38389),
            .I(N__38382));
    InMux I__8267 (
            .O(N__38388),
            .I(N__38379));
    InMux I__8266 (
            .O(N__38385),
            .I(N__38374));
    InMux I__8265 (
            .O(N__38382),
            .I(N__38374));
    LocalMux I__8264 (
            .O(N__38379),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    LocalMux I__8263 (
            .O(N__38374),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    InMux I__8262 (
            .O(N__38369),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ));
    InMux I__8261 (
            .O(N__38366),
            .I(N__38361));
    InMux I__8260 (
            .O(N__38365),
            .I(N__38356));
    InMux I__8259 (
            .O(N__38364),
            .I(N__38356));
    LocalMux I__8258 (
            .O(N__38361),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    LocalMux I__8257 (
            .O(N__38356),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    InMux I__8256 (
            .O(N__38351),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ));
    InMux I__8255 (
            .O(N__38348),
            .I(N__38343));
    InMux I__8254 (
            .O(N__38347),
            .I(N__38338));
    InMux I__8253 (
            .O(N__38346),
            .I(N__38338));
    LocalMux I__8252 (
            .O(N__38343),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    LocalMux I__8251 (
            .O(N__38338),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    InMux I__8250 (
            .O(N__38333),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ));
    InMux I__8249 (
            .O(N__38330),
            .I(N__38327));
    LocalMux I__8248 (
            .O(N__38327),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14 ));
    InMux I__8247 (
            .O(N__38324),
            .I(N__38321));
    LocalMux I__8246 (
            .O(N__38321),
            .I(N__38317));
    InMux I__8245 (
            .O(N__38320),
            .I(N__38314));
    Span4Mux_h I__8244 (
            .O(N__38317),
            .I(N__38311));
    LocalMux I__8243 (
            .O(N__38314),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14 ));
    Odrv4 I__8242 (
            .O(N__38311),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14 ));
    CascadeMux I__8241 (
            .O(N__38306),
            .I(N__38303));
    InMux I__8240 (
            .O(N__38303),
            .I(N__38300));
    LocalMux I__8239 (
            .O(N__38300),
            .I(N__38297));
    Span4Mux_v I__8238 (
            .O(N__38297),
            .I(N__38294));
    Odrv4 I__8237 (
            .O(N__38294),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0 ));
    CascadeMux I__8236 (
            .O(N__38291),
            .I(N__38288));
    InMux I__8235 (
            .O(N__38288),
            .I(N__38283));
    InMux I__8234 (
            .O(N__38287),
            .I(N__38280));
    InMux I__8233 (
            .O(N__38286),
            .I(N__38277));
    LocalMux I__8232 (
            .O(N__38283),
            .I(N__38274));
    LocalMux I__8231 (
            .O(N__38280),
            .I(N__38269));
    LocalMux I__8230 (
            .O(N__38277),
            .I(N__38269));
    Odrv4 I__8229 (
            .O(N__38274),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv12 I__8228 (
            .O(N__38269),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1 ));
    InMux I__8227 (
            .O(N__38264),
            .I(N__38261));
    LocalMux I__8226 (
            .O(N__38261),
            .I(N__38258));
    Span4Mux_h I__8225 (
            .O(N__38258),
            .I(N__38255));
    Odrv4 I__8224 (
            .O(N__38255),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2 ));
    InMux I__8223 (
            .O(N__38252),
            .I(N__38248));
    InMux I__8222 (
            .O(N__38251),
            .I(N__38245));
    LocalMux I__8221 (
            .O(N__38248),
            .I(N__38242));
    LocalMux I__8220 (
            .O(N__38245),
            .I(N__38239));
    Odrv4 I__8219 (
            .O(N__38242),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2 ));
    Odrv12 I__8218 (
            .O(N__38239),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2 ));
    CascadeMux I__8217 (
            .O(N__38234),
            .I(N__38231));
    InMux I__8216 (
            .O(N__38231),
            .I(N__38228));
    LocalMux I__8215 (
            .O(N__38228),
            .I(N__38225));
    Odrv4 I__8214 (
            .O(N__38225),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17 ));
    InMux I__8213 (
            .O(N__38222),
            .I(N__38219));
    LocalMux I__8212 (
            .O(N__38219),
            .I(N__38215));
    InMux I__8211 (
            .O(N__38218),
            .I(N__38212));
    Span4Mux_h I__8210 (
            .O(N__38215),
            .I(N__38209));
    LocalMux I__8209 (
            .O(N__38212),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17 ));
    Odrv4 I__8208 (
            .O(N__38209),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__8207 (
            .O(N__38204),
            .I(N__38201));
    LocalMux I__8206 (
            .O(N__38201),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18 ));
    InMux I__8205 (
            .O(N__38198),
            .I(N__38195));
    LocalMux I__8204 (
            .O(N__38195),
            .I(N__38191));
    InMux I__8203 (
            .O(N__38194),
            .I(N__38188));
    Span4Mux_h I__8202 (
            .O(N__38191),
            .I(N__38185));
    LocalMux I__8201 (
            .O(N__38188),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18 ));
    Odrv4 I__8200 (
            .O(N__38185),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18 ));
    CascadeMux I__8199 (
            .O(N__38180),
            .I(N__38170));
    CascadeMux I__8198 (
            .O(N__38179),
            .I(N__38167));
    InMux I__8197 (
            .O(N__38178),
            .I(N__38148));
    InMux I__8196 (
            .O(N__38177),
            .I(N__38148));
    InMux I__8195 (
            .O(N__38176),
            .I(N__38148));
    InMux I__8194 (
            .O(N__38175),
            .I(N__38148));
    InMux I__8193 (
            .O(N__38174),
            .I(N__38148));
    InMux I__8192 (
            .O(N__38173),
            .I(N__38127));
    InMux I__8191 (
            .O(N__38170),
            .I(N__38127));
    InMux I__8190 (
            .O(N__38167),
            .I(N__38127));
    InMux I__8189 (
            .O(N__38166),
            .I(N__38127));
    InMux I__8188 (
            .O(N__38165),
            .I(N__38127));
    InMux I__8187 (
            .O(N__38164),
            .I(N__38127));
    InMux I__8186 (
            .O(N__38163),
            .I(N__38127));
    InMux I__8185 (
            .O(N__38162),
            .I(N__38118));
    InMux I__8184 (
            .O(N__38161),
            .I(N__38118));
    InMux I__8183 (
            .O(N__38160),
            .I(N__38118));
    InMux I__8182 (
            .O(N__38159),
            .I(N__38118));
    LocalMux I__8181 (
            .O(N__38148),
            .I(N__38114));
    InMux I__8180 (
            .O(N__38147),
            .I(N__38107));
    InMux I__8179 (
            .O(N__38146),
            .I(N__38107));
    InMux I__8178 (
            .O(N__38145),
            .I(N__38107));
    CascadeMux I__8177 (
            .O(N__38144),
            .I(N__38104));
    InMux I__8176 (
            .O(N__38143),
            .I(N__38098));
    InMux I__8175 (
            .O(N__38142),
            .I(N__38098));
    LocalMux I__8174 (
            .O(N__38127),
            .I(N__38093));
    LocalMux I__8173 (
            .O(N__38118),
            .I(N__38093));
    InMux I__8172 (
            .O(N__38117),
            .I(N__38090));
    Span4Mux_h I__8171 (
            .O(N__38114),
            .I(N__38085));
    LocalMux I__8170 (
            .O(N__38107),
            .I(N__38085));
    InMux I__8169 (
            .O(N__38104),
            .I(N__38080));
    InMux I__8168 (
            .O(N__38103),
            .I(N__38080));
    LocalMux I__8167 (
            .O(N__38098),
            .I(N__38075));
    Span4Mux_v I__8166 (
            .O(N__38093),
            .I(N__38075));
    LocalMux I__8165 (
            .O(N__38090),
            .I(N__38072));
    Span4Mux_v I__8164 (
            .O(N__38085),
            .I(N__38069));
    LocalMux I__8163 (
            .O(N__38080),
            .I(N__38064));
    Span4Mux_v I__8162 (
            .O(N__38075),
            .I(N__38064));
    Span4Mux_h I__8161 (
            .O(N__38072),
            .I(N__38061));
    Span4Mux_v I__8160 (
            .O(N__38069),
            .I(N__38058));
    Odrv4 I__8159 (
            .O(N__38064),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__8158 (
            .O(N__38061),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__8157 (
            .O(N__38058),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ));
    CascadeMux I__8156 (
            .O(N__38051),
            .I(N__38040));
    CascadeMux I__8155 (
            .O(N__38050),
            .I(N__38034));
    CascadeMux I__8154 (
            .O(N__38049),
            .I(N__38031));
    CascadeMux I__8153 (
            .O(N__38048),
            .I(N__38028));
    CascadeMux I__8152 (
            .O(N__38047),
            .I(N__38025));
    CascadeMux I__8151 (
            .O(N__38046),
            .I(N__38019));
    InMux I__8150 (
            .O(N__38045),
            .I(N__38012));
    CascadeMux I__8149 (
            .O(N__38044),
            .I(N__38009));
    CascadeMux I__8148 (
            .O(N__38043),
            .I(N__38006));
    InMux I__8147 (
            .O(N__38040),
            .I(N__37999));
    InMux I__8146 (
            .O(N__38039),
            .I(N__37999));
    InMux I__8145 (
            .O(N__38038),
            .I(N__37987));
    InMux I__8144 (
            .O(N__38037),
            .I(N__37987));
    InMux I__8143 (
            .O(N__38034),
            .I(N__37987));
    InMux I__8142 (
            .O(N__38031),
            .I(N__37987));
    InMux I__8141 (
            .O(N__38028),
            .I(N__37987));
    InMux I__8140 (
            .O(N__38025),
            .I(N__37982));
    InMux I__8139 (
            .O(N__38024),
            .I(N__37982));
    InMux I__8138 (
            .O(N__38023),
            .I(N__37967));
    InMux I__8137 (
            .O(N__38022),
            .I(N__37967));
    InMux I__8136 (
            .O(N__38019),
            .I(N__37967));
    InMux I__8135 (
            .O(N__38018),
            .I(N__37967));
    InMux I__8134 (
            .O(N__38017),
            .I(N__37967));
    InMux I__8133 (
            .O(N__38016),
            .I(N__37967));
    InMux I__8132 (
            .O(N__38015),
            .I(N__37967));
    LocalMux I__8131 (
            .O(N__38012),
            .I(N__37964));
    InMux I__8130 (
            .O(N__38009),
            .I(N__37955));
    InMux I__8129 (
            .O(N__38006),
            .I(N__37955));
    InMux I__8128 (
            .O(N__38005),
            .I(N__37955));
    InMux I__8127 (
            .O(N__38004),
            .I(N__37955));
    LocalMux I__8126 (
            .O(N__37999),
            .I(N__37952));
    CascadeMux I__8125 (
            .O(N__37998),
            .I(N__37948));
    LocalMux I__8124 (
            .O(N__37987),
            .I(N__37944));
    LocalMux I__8123 (
            .O(N__37982),
            .I(N__37937));
    LocalMux I__8122 (
            .O(N__37967),
            .I(N__37937));
    Span4Mux_v I__8121 (
            .O(N__37964),
            .I(N__37937));
    LocalMux I__8120 (
            .O(N__37955),
            .I(N__37934));
    Sp12to4 I__8119 (
            .O(N__37952),
            .I(N__37931));
    InMux I__8118 (
            .O(N__37951),
            .I(N__37924));
    InMux I__8117 (
            .O(N__37948),
            .I(N__37924));
    InMux I__8116 (
            .O(N__37947),
            .I(N__37924));
    Span4Mux_h I__8115 (
            .O(N__37944),
            .I(N__37919));
    Span4Mux_v I__8114 (
            .O(N__37937),
            .I(N__37919));
    Odrv4 I__8113 (
            .O(N__37934),
            .I(\phase_controller_slave.start_timer_trZ0 ));
    Odrv12 I__8112 (
            .O(N__37931),
            .I(\phase_controller_slave.start_timer_trZ0 ));
    LocalMux I__8111 (
            .O(N__37924),
            .I(\phase_controller_slave.start_timer_trZ0 ));
    Odrv4 I__8110 (
            .O(N__37919),
            .I(\phase_controller_slave.start_timer_trZ0 ));
    CascadeMux I__8109 (
            .O(N__37910),
            .I(N__37907));
    InMux I__8108 (
            .O(N__37907),
            .I(N__37904));
    LocalMux I__8107 (
            .O(N__37904),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19 ));
    CascadeMux I__8106 (
            .O(N__37901),
            .I(N__37889));
    CascadeMux I__8105 (
            .O(N__37900),
            .I(N__37886));
    CascadeMux I__8104 (
            .O(N__37899),
            .I(N__37881));
    CascadeMux I__8103 (
            .O(N__37898),
            .I(N__37878));
    InMux I__8102 (
            .O(N__37897),
            .I(N__37862));
    InMux I__8101 (
            .O(N__37896),
            .I(N__37862));
    InMux I__8100 (
            .O(N__37895),
            .I(N__37862));
    InMux I__8099 (
            .O(N__37894),
            .I(N__37862));
    InMux I__8098 (
            .O(N__37893),
            .I(N__37862));
    InMux I__8097 (
            .O(N__37892),
            .I(N__37855));
    InMux I__8096 (
            .O(N__37889),
            .I(N__37850));
    InMux I__8095 (
            .O(N__37886),
            .I(N__37850));
    InMux I__8094 (
            .O(N__37885),
            .I(N__37845));
    InMux I__8093 (
            .O(N__37884),
            .I(N__37845));
    InMux I__8092 (
            .O(N__37881),
            .I(N__37830));
    InMux I__8091 (
            .O(N__37878),
            .I(N__37830));
    InMux I__8090 (
            .O(N__37877),
            .I(N__37830));
    InMux I__8089 (
            .O(N__37876),
            .I(N__37830));
    InMux I__8088 (
            .O(N__37875),
            .I(N__37830));
    InMux I__8087 (
            .O(N__37874),
            .I(N__37830));
    InMux I__8086 (
            .O(N__37873),
            .I(N__37830));
    LocalMux I__8085 (
            .O(N__37862),
            .I(N__37827));
    InMux I__8084 (
            .O(N__37861),
            .I(N__37823));
    InMux I__8083 (
            .O(N__37860),
            .I(N__37818));
    InMux I__8082 (
            .O(N__37859),
            .I(N__37818));
    InMux I__8081 (
            .O(N__37858),
            .I(N__37815));
    LocalMux I__8080 (
            .O(N__37855),
            .I(N__37812));
    LocalMux I__8079 (
            .O(N__37850),
            .I(N__37803));
    LocalMux I__8078 (
            .O(N__37845),
            .I(N__37803));
    LocalMux I__8077 (
            .O(N__37830),
            .I(N__37803));
    Span4Mux_v I__8076 (
            .O(N__37827),
            .I(N__37803));
    InMux I__8075 (
            .O(N__37826),
            .I(N__37800));
    LocalMux I__8074 (
            .O(N__37823),
            .I(N__37795));
    LocalMux I__8073 (
            .O(N__37818),
            .I(N__37795));
    LocalMux I__8072 (
            .O(N__37815),
            .I(N__37786));
    Span4Mux_h I__8071 (
            .O(N__37812),
            .I(N__37786));
    Span4Mux_v I__8070 (
            .O(N__37803),
            .I(N__37786));
    LocalMux I__8069 (
            .O(N__37800),
            .I(N__37783));
    Span4Mux_v I__8068 (
            .O(N__37795),
            .I(N__37780));
    InMux I__8067 (
            .O(N__37794),
            .I(N__37775));
    InMux I__8066 (
            .O(N__37793),
            .I(N__37775));
    Span4Mux_v I__8065 (
            .O(N__37786),
            .I(N__37770));
    Span4Mux_v I__8064 (
            .O(N__37783),
            .I(N__37770));
    Span4Mux_v I__8063 (
            .O(N__37780),
            .I(N__37767));
    LocalMux I__8062 (
            .O(N__37775),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__8061 (
            .O(N__37770),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__8060 (
            .O(N__37767),
            .I(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ));
    InMux I__8059 (
            .O(N__37760),
            .I(N__37757));
    LocalMux I__8058 (
            .O(N__37757),
            .I(N__37753));
    InMux I__8057 (
            .O(N__37756),
            .I(N__37750));
    Span4Mux_h I__8056 (
            .O(N__37753),
            .I(N__37747));
    LocalMux I__8055 (
            .O(N__37750),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19 ));
    Odrv4 I__8054 (
            .O(N__37747),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__8053 (
            .O(N__37742),
            .I(N__37739));
    LocalMux I__8052 (
            .O(N__37739),
            .I(N__37736));
    Odrv4 I__8051 (
            .O(N__37736),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10 ));
    InMux I__8050 (
            .O(N__37733),
            .I(N__37729));
    InMux I__8049 (
            .O(N__37732),
            .I(N__37726));
    LocalMux I__8048 (
            .O(N__37729),
            .I(N__37723));
    LocalMux I__8047 (
            .O(N__37726),
            .I(N__37720));
    Odrv12 I__8046 (
            .O(N__37723),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10 ));
    Odrv12 I__8045 (
            .O(N__37720),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10 ));
    InMux I__8044 (
            .O(N__37715),
            .I(N__37712));
    LocalMux I__8043 (
            .O(N__37712),
            .I(N__37709));
    Odrv4 I__8042 (
            .O(N__37709),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11 ));
    InMux I__8041 (
            .O(N__37706),
            .I(N__37702));
    InMux I__8040 (
            .O(N__37705),
            .I(N__37699));
    LocalMux I__8039 (
            .O(N__37702),
            .I(N__37696));
    LocalMux I__8038 (
            .O(N__37699),
            .I(N__37693));
    Span4Mux_v I__8037 (
            .O(N__37696),
            .I(N__37690));
    Odrv4 I__8036 (
            .O(N__37693),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11 ));
    Odrv4 I__8035 (
            .O(N__37690),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11 ));
    InMux I__8034 (
            .O(N__37685),
            .I(N__37682));
    LocalMux I__8033 (
            .O(N__37682),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15 ));
    InMux I__8032 (
            .O(N__37679),
            .I(N__37676));
    LocalMux I__8031 (
            .O(N__37676),
            .I(N__37672));
    InMux I__8030 (
            .O(N__37675),
            .I(N__37669));
    Span4Mux_h I__8029 (
            .O(N__37672),
            .I(N__37666));
    LocalMux I__8028 (
            .O(N__37669),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15 ));
    Odrv4 I__8027 (
            .O(N__37666),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__8026 (
            .O(N__37661),
            .I(N__37658));
    LocalMux I__8025 (
            .O(N__37658),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12 ));
    InMux I__8024 (
            .O(N__37655),
            .I(N__37652));
    LocalMux I__8023 (
            .O(N__37652),
            .I(N__37648));
    InMux I__8022 (
            .O(N__37651),
            .I(N__37645));
    Span4Mux_v I__8021 (
            .O(N__37648),
            .I(N__37642));
    LocalMux I__8020 (
            .O(N__37645),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12 ));
    Odrv4 I__8019 (
            .O(N__37642),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__8018 (
            .O(N__37637),
            .I(N__37634));
    LocalMux I__8017 (
            .O(N__37634),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16 ));
    InMux I__8016 (
            .O(N__37631),
            .I(N__37628));
    LocalMux I__8015 (
            .O(N__37628),
            .I(N__37624));
    InMux I__8014 (
            .O(N__37627),
            .I(N__37621));
    Span4Mux_v I__8013 (
            .O(N__37624),
            .I(N__37618));
    LocalMux I__8012 (
            .O(N__37621),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv4 I__8011 (
            .O(N__37618),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16 ));
    InMux I__8010 (
            .O(N__37613),
            .I(N__37610));
    LocalMux I__8009 (
            .O(N__37610),
            .I(N__37607));
    Span4Mux_h I__8008 (
            .O(N__37607),
            .I(N__37604));
    Odrv4 I__8007 (
            .O(N__37604),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4 ));
    InMux I__8006 (
            .O(N__37601),
            .I(N__37598));
    LocalMux I__8005 (
            .O(N__37598),
            .I(N__37594));
    InMux I__8004 (
            .O(N__37597),
            .I(N__37591));
    Span4Mux_v I__8003 (
            .O(N__37594),
            .I(N__37588));
    LocalMux I__8002 (
            .O(N__37591),
            .I(N__37585));
    Odrv4 I__8001 (
            .O(N__37588),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4 ));
    Odrv12 I__8000 (
            .O(N__37585),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4 ));
    InMux I__7999 (
            .O(N__37580),
            .I(N__37577));
    LocalMux I__7998 (
            .O(N__37577),
            .I(N__37574));
    Span4Mux_h I__7997 (
            .O(N__37574),
            .I(N__37571));
    Odrv4 I__7996 (
            .O(N__37571),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5 ));
    InMux I__7995 (
            .O(N__37568),
            .I(N__37565));
    LocalMux I__7994 (
            .O(N__37565),
            .I(N__37561));
    InMux I__7993 (
            .O(N__37564),
            .I(N__37558));
    Span4Mux_h I__7992 (
            .O(N__37561),
            .I(N__37555));
    LocalMux I__7991 (
            .O(N__37558),
            .I(N__37552));
    Odrv4 I__7990 (
            .O(N__37555),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5 ));
    Odrv12 I__7989 (
            .O(N__37552),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5 ));
    InMux I__7988 (
            .O(N__37547),
            .I(N__37544));
    LocalMux I__7987 (
            .O(N__37544),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13 ));
    InMux I__7986 (
            .O(N__37541),
            .I(N__37538));
    LocalMux I__7985 (
            .O(N__37538),
            .I(N__37534));
    InMux I__7984 (
            .O(N__37537),
            .I(N__37531));
    Span4Mux_h I__7983 (
            .O(N__37534),
            .I(N__37528));
    LocalMux I__7982 (
            .O(N__37531),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13 ));
    Odrv4 I__7981 (
            .O(N__37528),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__7980 (
            .O(N__37523),
            .I(N__37520));
    LocalMux I__7979 (
            .O(N__37520),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9 ));
    InMux I__7978 (
            .O(N__37517),
            .I(N__37514));
    LocalMux I__7977 (
            .O(N__37514),
            .I(N__37510));
    InMux I__7976 (
            .O(N__37513),
            .I(N__37507));
    Span4Mux_h I__7975 (
            .O(N__37510),
            .I(N__37504));
    LocalMux I__7974 (
            .O(N__37507),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9 ));
    Odrv4 I__7973 (
            .O(N__37504),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9 ));
    CascadeMux I__7972 (
            .O(N__37499),
            .I(N__37496));
    InMux I__7971 (
            .O(N__37496),
            .I(N__37493));
    LocalMux I__7970 (
            .O(N__37493),
            .I(N__37490));
    Odrv12 I__7969 (
            .O(N__37490),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6 ));
    InMux I__7968 (
            .O(N__37487),
            .I(N__37483));
    InMux I__7967 (
            .O(N__37486),
            .I(N__37480));
    LocalMux I__7966 (
            .O(N__37483),
            .I(N__37477));
    LocalMux I__7965 (
            .O(N__37480),
            .I(N__37474));
    Odrv4 I__7964 (
            .O(N__37477),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6 ));
    Odrv12 I__7963 (
            .O(N__37474),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6 ));
    CascadeMux I__7962 (
            .O(N__37469),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1_cascade_ ));
    InMux I__7961 (
            .O(N__37466),
            .I(N__37457));
    InMux I__7960 (
            .O(N__37465),
            .I(N__37457));
    InMux I__7959 (
            .O(N__37464),
            .I(N__37457));
    LocalMux I__7958 (
            .O(N__37457),
            .I(N__37451));
    InMux I__7957 (
            .O(N__37456),
            .I(N__37444));
    InMux I__7956 (
            .O(N__37455),
            .I(N__37444));
    InMux I__7955 (
            .O(N__37454),
            .I(N__37444));
    Odrv4 I__7954 (
            .O(N__37451),
            .I(\phase_controller_inst1.stoper_tr.N_20_li ));
    LocalMux I__7953 (
            .O(N__37444),
            .I(\phase_controller_inst1.stoper_tr.N_20_li ));
    InMux I__7952 (
            .O(N__37439),
            .I(N__37434));
    InMux I__7951 (
            .O(N__37438),
            .I(N__37429));
    InMux I__7950 (
            .O(N__37437),
            .I(N__37429));
    LocalMux I__7949 (
            .O(N__37434),
            .I(N__37424));
    LocalMux I__7948 (
            .O(N__37429),
            .I(N__37424));
    Span4Mux_h I__7947 (
            .O(N__37424),
            .I(N__37419));
    InMux I__7946 (
            .O(N__37423),
            .I(N__37414));
    InMux I__7945 (
            .O(N__37422),
            .I(N__37414));
    Odrv4 I__7944 (
            .O(N__37419),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3 ));
    LocalMux I__7943 (
            .O(N__37414),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3 ));
    InMux I__7942 (
            .O(N__37409),
            .I(N__37406));
    LocalMux I__7941 (
            .O(N__37406),
            .I(N__37402));
    CascadeMux I__7940 (
            .O(N__37405),
            .I(N__37399));
    Span4Mux_v I__7939 (
            .O(N__37402),
            .I(N__37395));
    InMux I__7938 (
            .O(N__37399),
            .I(N__37390));
    InMux I__7937 (
            .O(N__37398),
            .I(N__37390));
    Odrv4 I__7936 (
            .O(N__37395),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    LocalMux I__7935 (
            .O(N__37390),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    InMux I__7934 (
            .O(N__37385),
            .I(N__37382));
    LocalMux I__7933 (
            .O(N__37382),
            .I(N__37379));
    Span4Mux_v I__7932 (
            .O(N__37379),
            .I(N__37375));
    InMux I__7931 (
            .O(N__37378),
            .I(N__37372));
    Span4Mux_v I__7930 (
            .O(N__37375),
            .I(N__37369));
    LocalMux I__7929 (
            .O(N__37372),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    Odrv4 I__7928 (
            .O(N__37369),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    InMux I__7927 (
            .O(N__37364),
            .I(N__37354));
    InMux I__7926 (
            .O(N__37363),
            .I(N__37354));
    InMux I__7925 (
            .O(N__37362),
            .I(N__37354));
    InMux I__7924 (
            .O(N__37361),
            .I(N__37351));
    LocalMux I__7923 (
            .O(N__37354),
            .I(N__37346));
    LocalMux I__7922 (
            .O(N__37351),
            .I(N__37343));
    InMux I__7921 (
            .O(N__37350),
            .I(N__37338));
    InMux I__7920 (
            .O(N__37349),
            .I(N__37338));
    Span4Mux_v I__7919 (
            .O(N__37346),
            .I(N__37333));
    Span4Mux_h I__7918 (
            .O(N__37343),
            .I(N__37333));
    LocalMux I__7917 (
            .O(N__37338),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6 ));
    Odrv4 I__7916 (
            .O(N__37333),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6 ));
    InMux I__7915 (
            .O(N__37328),
            .I(N__37323));
    InMux I__7914 (
            .O(N__37327),
            .I(N__37320));
    InMux I__7913 (
            .O(N__37326),
            .I(N__37317));
    LocalMux I__7912 (
            .O(N__37323),
            .I(N__37314));
    LocalMux I__7911 (
            .O(N__37320),
            .I(N__37310));
    LocalMux I__7910 (
            .O(N__37317),
            .I(N__37307));
    Span4Mux_v I__7909 (
            .O(N__37314),
            .I(N__37304));
    CascadeMux I__7908 (
            .O(N__37313),
            .I(N__37301));
    Span4Mux_v I__7907 (
            .O(N__37310),
            .I(N__37296));
    Span4Mux_h I__7906 (
            .O(N__37307),
            .I(N__37296));
    Span4Mux_v I__7905 (
            .O(N__37304),
            .I(N__37293));
    InMux I__7904 (
            .O(N__37301),
            .I(N__37290));
    Span4Mux_v I__7903 (
            .O(N__37296),
            .I(N__37287));
    Odrv4 I__7902 (
            .O(N__37293),
            .I(measured_delay_tr_7));
    LocalMux I__7901 (
            .O(N__37290),
            .I(measured_delay_tr_7));
    Odrv4 I__7900 (
            .O(N__37287),
            .I(measured_delay_tr_7));
    InMux I__7899 (
            .O(N__37280),
            .I(N__37264));
    InMux I__7898 (
            .O(N__37279),
            .I(N__37264));
    InMux I__7897 (
            .O(N__37278),
            .I(N__37264));
    InMux I__7896 (
            .O(N__37277),
            .I(N__37264));
    InMux I__7895 (
            .O(N__37276),
            .I(N__37264));
    InMux I__7894 (
            .O(N__37275),
            .I(N__37261));
    LocalMux I__7893 (
            .O(N__37264),
            .I(N__37257));
    LocalMux I__7892 (
            .O(N__37261),
            .I(N__37251));
    InMux I__7891 (
            .O(N__37260),
            .I(N__37248));
    Span4Mux_h I__7890 (
            .O(N__37257),
            .I(N__37245));
    InMux I__7889 (
            .O(N__37256),
            .I(N__37238));
    InMux I__7888 (
            .O(N__37255),
            .I(N__37238));
    InMux I__7887 (
            .O(N__37254),
            .I(N__37238));
    Span4Mux_h I__7886 (
            .O(N__37251),
            .I(N__37235));
    LocalMux I__7885 (
            .O(N__37248),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6 ));
    Odrv4 I__7884 (
            .O(N__37245),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6 ));
    LocalMux I__7883 (
            .O(N__37238),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6 ));
    Odrv4 I__7882 (
            .O(N__37235),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6 ));
    InMux I__7881 (
            .O(N__37226),
            .I(N__37221));
    InMux I__7880 (
            .O(N__37225),
            .I(N__37218));
    InMux I__7879 (
            .O(N__37224),
            .I(N__37215));
    LocalMux I__7878 (
            .O(N__37221),
            .I(N__37212));
    LocalMux I__7877 (
            .O(N__37218),
            .I(N__37209));
    LocalMux I__7876 (
            .O(N__37215),
            .I(N__37206));
    Span4Mux_h I__7875 (
            .O(N__37212),
            .I(N__37203));
    Span4Mux_v I__7874 (
            .O(N__37209),
            .I(N__37197));
    Span4Mux_h I__7873 (
            .O(N__37206),
            .I(N__37197));
    Span4Mux_v I__7872 (
            .O(N__37203),
            .I(N__37194));
    InMux I__7871 (
            .O(N__37202),
            .I(N__37191));
    Span4Mux_v I__7870 (
            .O(N__37197),
            .I(N__37188));
    Odrv4 I__7869 (
            .O(N__37194),
            .I(measured_delay_tr_8));
    LocalMux I__7868 (
            .O(N__37191),
            .I(measured_delay_tr_8));
    Odrv4 I__7867 (
            .O(N__37188),
            .I(measured_delay_tr_8));
    InMux I__7866 (
            .O(N__37181),
            .I(N__37178));
    LocalMux I__7865 (
            .O(N__37178),
            .I(N__37175));
    Span4Mux_v I__7864 (
            .O(N__37175),
            .I(N__37171));
    InMux I__7863 (
            .O(N__37174),
            .I(N__37168));
    Span4Mux_h I__7862 (
            .O(N__37171),
            .I(N__37165));
    LocalMux I__7861 (
            .O(N__37168),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16 ));
    Odrv4 I__7860 (
            .O(N__37165),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16 ));
    InMux I__7859 (
            .O(N__37160),
            .I(N__37157));
    LocalMux I__7858 (
            .O(N__37157),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_16 ));
    InMux I__7857 (
            .O(N__37154),
            .I(N__37151));
    LocalMux I__7856 (
            .O(N__37151),
            .I(N__37147));
    InMux I__7855 (
            .O(N__37150),
            .I(N__37144));
    Span4Mux_v I__7854 (
            .O(N__37147),
            .I(N__37141));
    LocalMux I__7853 (
            .O(N__37144),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17 ));
    Odrv4 I__7852 (
            .O(N__37141),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17 ));
    InMux I__7851 (
            .O(N__37136),
            .I(N__37133));
    LocalMux I__7850 (
            .O(N__37133),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_17 ));
    InMux I__7849 (
            .O(N__37130),
            .I(N__37127));
    LocalMux I__7848 (
            .O(N__37127),
            .I(N__37123));
    InMux I__7847 (
            .O(N__37126),
            .I(N__37120));
    Span4Mux_v I__7846 (
            .O(N__37123),
            .I(N__37117));
    LocalMux I__7845 (
            .O(N__37120),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18 ));
    Odrv4 I__7844 (
            .O(N__37117),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18 ));
    CascadeMux I__7843 (
            .O(N__37112),
            .I(N__37109));
    InMux I__7842 (
            .O(N__37109),
            .I(N__37106));
    LocalMux I__7841 (
            .O(N__37106),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_18 ));
    InMux I__7840 (
            .O(N__37103),
            .I(N__37100));
    LocalMux I__7839 (
            .O(N__37100),
            .I(N__37096));
    InMux I__7838 (
            .O(N__37099),
            .I(N__37093));
    Span12Mux_v I__7837 (
            .O(N__37096),
            .I(N__37090));
    LocalMux I__7836 (
            .O(N__37093),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19 ));
    Odrv12 I__7835 (
            .O(N__37090),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__7834 (
            .O(N__37085),
            .I(N__37082));
    LocalMux I__7833 (
            .O(N__37082),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_19 ));
    InMux I__7832 (
            .O(N__37079),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19 ));
    InMux I__7831 (
            .O(N__37076),
            .I(N__37072));
    InMux I__7830 (
            .O(N__37075),
            .I(N__37069));
    LocalMux I__7829 (
            .O(N__37072),
            .I(N__37066));
    LocalMux I__7828 (
            .O(N__37069),
            .I(N__37063));
    Span4Mux_v I__7827 (
            .O(N__37066),
            .I(N__37059));
    Span4Mux_h I__7826 (
            .O(N__37063),
            .I(N__37056));
    InMux I__7825 (
            .O(N__37062),
            .I(N__37053));
    Odrv4 I__7824 (
            .O(N__37059),
            .I(\phase_controller_slave.stoper_hc.time_passed11 ));
    Odrv4 I__7823 (
            .O(N__37056),
            .I(\phase_controller_slave.stoper_hc.time_passed11 ));
    LocalMux I__7822 (
            .O(N__37053),
            .I(\phase_controller_slave.stoper_hc.time_passed11 ));
    InMux I__7821 (
            .O(N__37046),
            .I(N__37043));
    LocalMux I__7820 (
            .O(N__37043),
            .I(N__37040));
    Span4Mux_v I__7819 (
            .O(N__37040),
            .I(N__37037));
    Odrv4 I__7818 (
            .O(N__37037),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1 ));
    InMux I__7817 (
            .O(N__37034),
            .I(N__37031));
    LocalMux I__7816 (
            .O(N__37031),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_9 ));
    CascadeMux I__7815 (
            .O(N__37028),
            .I(N__37025));
    InMux I__7814 (
            .O(N__37025),
            .I(N__37022));
    LocalMux I__7813 (
            .O(N__37022),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_9 ));
    CascadeMux I__7812 (
            .O(N__37019),
            .I(N__37016));
    InMux I__7811 (
            .O(N__37016),
            .I(N__37013));
    LocalMux I__7810 (
            .O(N__37013),
            .I(N__37010));
    Span4Mux_h I__7809 (
            .O(N__37010),
            .I(N__37007));
    Odrv4 I__7808 (
            .O(N__37007),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_10 ));
    InMux I__7807 (
            .O(N__37004),
            .I(N__37001));
    LocalMux I__7806 (
            .O(N__37001),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_10 ));
    CascadeMux I__7805 (
            .O(N__36998),
            .I(N__36995));
    InMux I__7804 (
            .O(N__36995),
            .I(N__36992));
    LocalMux I__7803 (
            .O(N__36992),
            .I(N__36989));
    Odrv4 I__7802 (
            .O(N__36989),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_11 ));
    InMux I__7801 (
            .O(N__36986),
            .I(N__36983));
    LocalMux I__7800 (
            .O(N__36983),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_11 ));
    CascadeMux I__7799 (
            .O(N__36980),
            .I(N__36977));
    InMux I__7798 (
            .O(N__36977),
            .I(N__36974));
    LocalMux I__7797 (
            .O(N__36974),
            .I(N__36971));
    Odrv4 I__7796 (
            .O(N__36971),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_12 ));
    InMux I__7795 (
            .O(N__36968),
            .I(N__36965));
    LocalMux I__7794 (
            .O(N__36965),
            .I(N__36962));
    Span4Mux_h I__7793 (
            .O(N__36962),
            .I(N__36958));
    InMux I__7792 (
            .O(N__36961),
            .I(N__36955));
    Span4Mux_v I__7791 (
            .O(N__36958),
            .I(N__36952));
    LocalMux I__7790 (
            .O(N__36955),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12 ));
    Odrv4 I__7789 (
            .O(N__36952),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__7788 (
            .O(N__36947),
            .I(N__36944));
    LocalMux I__7787 (
            .O(N__36944),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_12 ));
    InMux I__7786 (
            .O(N__36941),
            .I(N__36938));
    LocalMux I__7785 (
            .O(N__36938),
            .I(N__36935));
    Span4Mux_h I__7784 (
            .O(N__36935),
            .I(N__36931));
    InMux I__7783 (
            .O(N__36934),
            .I(N__36928));
    Span4Mux_v I__7782 (
            .O(N__36931),
            .I(N__36925));
    LocalMux I__7781 (
            .O(N__36928),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13 ));
    Odrv4 I__7780 (
            .O(N__36925),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__7779 (
            .O(N__36920),
            .I(N__36917));
    LocalMux I__7778 (
            .O(N__36917),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_13 ));
    CascadeMux I__7777 (
            .O(N__36914),
            .I(N__36911));
    InMux I__7776 (
            .O(N__36911),
            .I(N__36908));
    LocalMux I__7775 (
            .O(N__36908),
            .I(N__36905));
    Span4Mux_v I__7774 (
            .O(N__36905),
            .I(N__36902));
    Odrv4 I__7773 (
            .O(N__36902),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_14 ));
    InMux I__7772 (
            .O(N__36899),
            .I(N__36896));
    LocalMux I__7771 (
            .O(N__36896),
            .I(N__36892));
    InMux I__7770 (
            .O(N__36895),
            .I(N__36889));
    Span12Mux_h I__7769 (
            .O(N__36892),
            .I(N__36886));
    LocalMux I__7768 (
            .O(N__36889),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14 ));
    Odrv12 I__7767 (
            .O(N__36886),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14 ));
    InMux I__7766 (
            .O(N__36881),
            .I(N__36878));
    LocalMux I__7765 (
            .O(N__36878),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_14 ));
    CascadeMux I__7764 (
            .O(N__36875),
            .I(N__36872));
    InMux I__7763 (
            .O(N__36872),
            .I(N__36869));
    LocalMux I__7762 (
            .O(N__36869),
            .I(N__36866));
    Span4Mux_h I__7761 (
            .O(N__36866),
            .I(N__36863));
    Odrv4 I__7760 (
            .O(N__36863),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_15 ));
    InMux I__7759 (
            .O(N__36860),
            .I(N__36857));
    LocalMux I__7758 (
            .O(N__36857),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_15 ));
    InMux I__7757 (
            .O(N__36854),
            .I(N__36851));
    LocalMux I__7756 (
            .O(N__36851),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_1 ));
    CascadeMux I__7755 (
            .O(N__36848),
            .I(N__36845));
    InMux I__7754 (
            .O(N__36845),
            .I(N__36842));
    LocalMux I__7753 (
            .O(N__36842),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_2 ));
    InMux I__7752 (
            .O(N__36839),
            .I(N__36836));
    LocalMux I__7751 (
            .O(N__36836),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_2 ));
    CascadeMux I__7750 (
            .O(N__36833),
            .I(N__36830));
    InMux I__7749 (
            .O(N__36830),
            .I(N__36827));
    LocalMux I__7748 (
            .O(N__36827),
            .I(N__36823));
    InMux I__7747 (
            .O(N__36826),
            .I(N__36820));
    Span4Mux_v I__7746 (
            .O(N__36823),
            .I(N__36817));
    LocalMux I__7745 (
            .O(N__36820),
            .I(N__36814));
    Odrv4 I__7744 (
            .O(N__36817),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3 ));
    Odrv4 I__7743 (
            .O(N__36814),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3 ));
    CascadeMux I__7742 (
            .O(N__36809),
            .I(N__36806));
    InMux I__7741 (
            .O(N__36806),
            .I(N__36803));
    LocalMux I__7740 (
            .O(N__36803),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_3 ));
    InMux I__7739 (
            .O(N__36800),
            .I(N__36797));
    LocalMux I__7738 (
            .O(N__36797),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_3 ));
    CascadeMux I__7737 (
            .O(N__36794),
            .I(N__36791));
    InMux I__7736 (
            .O(N__36791),
            .I(N__36788));
    LocalMux I__7735 (
            .O(N__36788),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_4 ));
    InMux I__7734 (
            .O(N__36785),
            .I(N__36782));
    LocalMux I__7733 (
            .O(N__36782),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_4 ));
    InMux I__7732 (
            .O(N__36779),
            .I(N__36776));
    LocalMux I__7731 (
            .O(N__36776),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_5 ));
    CascadeMux I__7730 (
            .O(N__36773),
            .I(N__36770));
    InMux I__7729 (
            .O(N__36770),
            .I(N__36767));
    LocalMux I__7728 (
            .O(N__36767),
            .I(\phase_controller_slave.stoper_hc.target_timeZ1Z_6 ));
    InMux I__7727 (
            .O(N__36764),
            .I(N__36761));
    LocalMux I__7726 (
            .O(N__36761),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_6 ));
    CascadeMux I__7725 (
            .O(N__36758),
            .I(N__36755));
    InMux I__7724 (
            .O(N__36755),
            .I(N__36752));
    LocalMux I__7723 (
            .O(N__36752),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_7 ));
    InMux I__7722 (
            .O(N__36749),
            .I(N__36746));
    LocalMux I__7721 (
            .O(N__36746),
            .I(N__36743));
    Sp12to4 I__7720 (
            .O(N__36743),
            .I(N__36739));
    InMux I__7719 (
            .O(N__36742),
            .I(N__36736));
    Odrv12 I__7718 (
            .O(N__36739),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7 ));
    LocalMux I__7717 (
            .O(N__36736),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7 ));
    InMux I__7716 (
            .O(N__36731),
            .I(N__36728));
    LocalMux I__7715 (
            .O(N__36728),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_7 ));
    InMux I__7714 (
            .O(N__36725),
            .I(N__36722));
    LocalMux I__7713 (
            .O(N__36722),
            .I(N__36719));
    Span4Mux_v I__7712 (
            .O(N__36719),
            .I(N__36715));
    InMux I__7711 (
            .O(N__36718),
            .I(N__36712));
    Odrv4 I__7710 (
            .O(N__36715),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8 ));
    LocalMux I__7709 (
            .O(N__36712),
            .I(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8 ));
    InMux I__7708 (
            .O(N__36707),
            .I(N__36704));
    LocalMux I__7707 (
            .O(N__36704),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_i_8 ));
    CascadeMux I__7706 (
            .O(N__36701),
            .I(N__36697));
    CascadeMux I__7705 (
            .O(N__36700),
            .I(N__36694));
    InMux I__7704 (
            .O(N__36697),
            .I(N__36688));
    InMux I__7703 (
            .O(N__36694),
            .I(N__36688));
    InMux I__7702 (
            .O(N__36693),
            .I(N__36685));
    LocalMux I__7701 (
            .O(N__36688),
            .I(N__36682));
    LocalMux I__7700 (
            .O(N__36685),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    Odrv12 I__7699 (
            .O(N__36682),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    InMux I__7698 (
            .O(N__36677),
            .I(\current_shift_inst.timer_s1.counter_cry_22 ));
    InMux I__7697 (
            .O(N__36674),
            .I(N__36670));
    InMux I__7696 (
            .O(N__36673),
            .I(N__36666));
    LocalMux I__7695 (
            .O(N__36670),
            .I(N__36663));
    InMux I__7694 (
            .O(N__36669),
            .I(N__36660));
    LocalMux I__7693 (
            .O(N__36666),
            .I(N__36655));
    Span4Mux_v I__7692 (
            .O(N__36663),
            .I(N__36655));
    LocalMux I__7691 (
            .O(N__36660),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    Odrv4 I__7690 (
            .O(N__36655),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    InMux I__7689 (
            .O(N__36650),
            .I(bfn_15_16_0_));
    InMux I__7688 (
            .O(N__36647),
            .I(N__36643));
    InMux I__7687 (
            .O(N__36646),
            .I(N__36639));
    LocalMux I__7686 (
            .O(N__36643),
            .I(N__36636));
    InMux I__7685 (
            .O(N__36642),
            .I(N__36633));
    LocalMux I__7684 (
            .O(N__36639),
            .I(N__36628));
    Span4Mux_v I__7683 (
            .O(N__36636),
            .I(N__36628));
    LocalMux I__7682 (
            .O(N__36633),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    Odrv4 I__7681 (
            .O(N__36628),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    InMux I__7680 (
            .O(N__36623),
            .I(\current_shift_inst.timer_s1.counter_cry_24 ));
    CascadeMux I__7679 (
            .O(N__36620),
            .I(N__36616));
    CascadeMux I__7678 (
            .O(N__36619),
            .I(N__36613));
    InMux I__7677 (
            .O(N__36616),
            .I(N__36607));
    InMux I__7676 (
            .O(N__36613),
            .I(N__36607));
    InMux I__7675 (
            .O(N__36612),
            .I(N__36604));
    LocalMux I__7674 (
            .O(N__36607),
            .I(N__36601));
    LocalMux I__7673 (
            .O(N__36604),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    Odrv4 I__7672 (
            .O(N__36601),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    InMux I__7671 (
            .O(N__36596),
            .I(\current_shift_inst.timer_s1.counter_cry_25 ));
    CascadeMux I__7670 (
            .O(N__36593),
            .I(N__36589));
    CascadeMux I__7669 (
            .O(N__36592),
            .I(N__36586));
    InMux I__7668 (
            .O(N__36589),
            .I(N__36580));
    InMux I__7667 (
            .O(N__36586),
            .I(N__36580));
    InMux I__7666 (
            .O(N__36585),
            .I(N__36577));
    LocalMux I__7665 (
            .O(N__36580),
            .I(N__36574));
    LocalMux I__7664 (
            .O(N__36577),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    Odrv4 I__7663 (
            .O(N__36574),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    InMux I__7662 (
            .O(N__36569),
            .I(\current_shift_inst.timer_s1.counter_cry_26 ));
    InMux I__7661 (
            .O(N__36566),
            .I(N__36562));
    InMux I__7660 (
            .O(N__36565),
            .I(N__36559));
    LocalMux I__7659 (
            .O(N__36562),
            .I(N__36556));
    LocalMux I__7658 (
            .O(N__36559),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    Odrv12 I__7657 (
            .O(N__36556),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    InMux I__7656 (
            .O(N__36551),
            .I(\current_shift_inst.timer_s1.counter_cry_27 ));
    InMux I__7655 (
            .O(N__36548),
            .I(N__36510));
    InMux I__7654 (
            .O(N__36547),
            .I(N__36510));
    InMux I__7653 (
            .O(N__36546),
            .I(N__36510));
    InMux I__7652 (
            .O(N__36545),
            .I(N__36510));
    InMux I__7651 (
            .O(N__36544),
            .I(N__36501));
    InMux I__7650 (
            .O(N__36543),
            .I(N__36501));
    InMux I__7649 (
            .O(N__36542),
            .I(N__36501));
    InMux I__7648 (
            .O(N__36541),
            .I(N__36501));
    InMux I__7647 (
            .O(N__36540),
            .I(N__36492));
    InMux I__7646 (
            .O(N__36539),
            .I(N__36492));
    InMux I__7645 (
            .O(N__36538),
            .I(N__36492));
    InMux I__7644 (
            .O(N__36537),
            .I(N__36492));
    InMux I__7643 (
            .O(N__36536),
            .I(N__36483));
    InMux I__7642 (
            .O(N__36535),
            .I(N__36483));
    InMux I__7641 (
            .O(N__36534),
            .I(N__36483));
    InMux I__7640 (
            .O(N__36533),
            .I(N__36483));
    InMux I__7639 (
            .O(N__36532),
            .I(N__36478));
    InMux I__7638 (
            .O(N__36531),
            .I(N__36478));
    InMux I__7637 (
            .O(N__36530),
            .I(N__36469));
    InMux I__7636 (
            .O(N__36529),
            .I(N__36469));
    InMux I__7635 (
            .O(N__36528),
            .I(N__36469));
    InMux I__7634 (
            .O(N__36527),
            .I(N__36469));
    InMux I__7633 (
            .O(N__36526),
            .I(N__36460));
    InMux I__7632 (
            .O(N__36525),
            .I(N__36460));
    InMux I__7631 (
            .O(N__36524),
            .I(N__36460));
    InMux I__7630 (
            .O(N__36523),
            .I(N__36460));
    InMux I__7629 (
            .O(N__36522),
            .I(N__36451));
    InMux I__7628 (
            .O(N__36521),
            .I(N__36451));
    InMux I__7627 (
            .O(N__36520),
            .I(N__36451));
    InMux I__7626 (
            .O(N__36519),
            .I(N__36451));
    LocalMux I__7625 (
            .O(N__36510),
            .I(N__36448));
    LocalMux I__7624 (
            .O(N__36501),
            .I(N__36433));
    LocalMux I__7623 (
            .O(N__36492),
            .I(N__36433));
    LocalMux I__7622 (
            .O(N__36483),
            .I(N__36433));
    LocalMux I__7621 (
            .O(N__36478),
            .I(N__36433));
    LocalMux I__7620 (
            .O(N__36469),
            .I(N__36433));
    LocalMux I__7619 (
            .O(N__36460),
            .I(N__36433));
    LocalMux I__7618 (
            .O(N__36451),
            .I(N__36433));
    Odrv4 I__7617 (
            .O(N__36448),
            .I(\current_shift_inst.timer_s1.running_i ));
    Odrv12 I__7616 (
            .O(N__36433),
            .I(\current_shift_inst.timer_s1.running_i ));
    InMux I__7615 (
            .O(N__36428),
            .I(\current_shift_inst.timer_s1.counter_cry_28 ));
    InMux I__7614 (
            .O(N__36425),
            .I(N__36421));
    InMux I__7613 (
            .O(N__36424),
            .I(N__36418));
    LocalMux I__7612 (
            .O(N__36421),
            .I(N__36415));
    LocalMux I__7611 (
            .O(N__36418),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    Odrv12 I__7610 (
            .O(N__36415),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    CEMux I__7609 (
            .O(N__36410),
            .I(N__36404));
    CEMux I__7608 (
            .O(N__36409),
            .I(N__36401));
    CEMux I__7607 (
            .O(N__36408),
            .I(N__36398));
    CEMux I__7606 (
            .O(N__36407),
            .I(N__36395));
    LocalMux I__7605 (
            .O(N__36404),
            .I(N__36390));
    LocalMux I__7604 (
            .O(N__36401),
            .I(N__36390));
    LocalMux I__7603 (
            .O(N__36398),
            .I(N__36385));
    LocalMux I__7602 (
            .O(N__36395),
            .I(N__36385));
    Span4Mux_v I__7601 (
            .O(N__36390),
            .I(N__36382));
    Span4Mux_v I__7600 (
            .O(N__36385),
            .I(N__36377));
    Span4Mux_h I__7599 (
            .O(N__36382),
            .I(N__36377));
    Span4Mux_v I__7598 (
            .O(N__36377),
            .I(N__36374));
    Odrv4 I__7597 (
            .O(N__36374),
            .I(\current_shift_inst.timer_s1.N_191_i ));
    InMux I__7596 (
            .O(N__36371),
            .I(N__36368));
    LocalMux I__7595 (
            .O(N__36368),
            .I(\phase_controller_slave.stoper_hc.target_timeZ0Z_0 ));
    CascadeMux I__7594 (
            .O(N__36365),
            .I(N__36361));
    CascadeMux I__7593 (
            .O(N__36364),
            .I(N__36358));
    InMux I__7592 (
            .O(N__36361),
            .I(N__36352));
    InMux I__7591 (
            .O(N__36358),
            .I(N__36352));
    InMux I__7590 (
            .O(N__36357),
            .I(N__36349));
    LocalMux I__7589 (
            .O(N__36352),
            .I(N__36346));
    LocalMux I__7588 (
            .O(N__36349),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    Odrv12 I__7587 (
            .O(N__36346),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    InMux I__7586 (
            .O(N__36341),
            .I(\current_shift_inst.timer_s1.counter_cry_13 ));
    CascadeMux I__7585 (
            .O(N__36338),
            .I(N__36334));
    CascadeMux I__7584 (
            .O(N__36337),
            .I(N__36331));
    InMux I__7583 (
            .O(N__36334),
            .I(N__36325));
    InMux I__7582 (
            .O(N__36331),
            .I(N__36325));
    InMux I__7581 (
            .O(N__36330),
            .I(N__36322));
    LocalMux I__7580 (
            .O(N__36325),
            .I(N__36319));
    LocalMux I__7579 (
            .O(N__36322),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    Odrv4 I__7578 (
            .O(N__36319),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    InMux I__7577 (
            .O(N__36314),
            .I(\current_shift_inst.timer_s1.counter_cry_14 ));
    InMux I__7576 (
            .O(N__36311),
            .I(N__36307));
    InMux I__7575 (
            .O(N__36310),
            .I(N__36304));
    LocalMux I__7574 (
            .O(N__36307),
            .I(N__36300));
    LocalMux I__7573 (
            .O(N__36304),
            .I(N__36297));
    InMux I__7572 (
            .O(N__36303),
            .I(N__36294));
    Span4Mux_h I__7571 (
            .O(N__36300),
            .I(N__36289));
    Span4Mux_v I__7570 (
            .O(N__36297),
            .I(N__36289));
    LocalMux I__7569 (
            .O(N__36294),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    Odrv4 I__7568 (
            .O(N__36289),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    InMux I__7567 (
            .O(N__36284),
            .I(bfn_15_15_0_));
    InMux I__7566 (
            .O(N__36281),
            .I(N__36277));
    InMux I__7565 (
            .O(N__36280),
            .I(N__36273));
    LocalMux I__7564 (
            .O(N__36277),
            .I(N__36270));
    InMux I__7563 (
            .O(N__36276),
            .I(N__36267));
    LocalMux I__7562 (
            .O(N__36273),
            .I(N__36262));
    Span4Mux_v I__7561 (
            .O(N__36270),
            .I(N__36262));
    LocalMux I__7560 (
            .O(N__36267),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    Odrv4 I__7559 (
            .O(N__36262),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    InMux I__7558 (
            .O(N__36257),
            .I(\current_shift_inst.timer_s1.counter_cry_16 ));
    CascadeMux I__7557 (
            .O(N__36254),
            .I(N__36250));
    CascadeMux I__7556 (
            .O(N__36253),
            .I(N__36247));
    InMux I__7555 (
            .O(N__36250),
            .I(N__36241));
    InMux I__7554 (
            .O(N__36247),
            .I(N__36241));
    InMux I__7553 (
            .O(N__36246),
            .I(N__36238));
    LocalMux I__7552 (
            .O(N__36241),
            .I(N__36235));
    LocalMux I__7551 (
            .O(N__36238),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    Odrv4 I__7550 (
            .O(N__36235),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    InMux I__7549 (
            .O(N__36230),
            .I(\current_shift_inst.timer_s1.counter_cry_17 ));
    CascadeMux I__7548 (
            .O(N__36227),
            .I(N__36223));
    CascadeMux I__7547 (
            .O(N__36226),
            .I(N__36220));
    InMux I__7546 (
            .O(N__36223),
            .I(N__36214));
    InMux I__7545 (
            .O(N__36220),
            .I(N__36214));
    InMux I__7544 (
            .O(N__36219),
            .I(N__36211));
    LocalMux I__7543 (
            .O(N__36214),
            .I(N__36208));
    LocalMux I__7542 (
            .O(N__36211),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    Odrv4 I__7541 (
            .O(N__36208),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    InMux I__7540 (
            .O(N__36203),
            .I(\current_shift_inst.timer_s1.counter_cry_18 ));
    InMux I__7539 (
            .O(N__36200),
            .I(N__36193));
    InMux I__7538 (
            .O(N__36199),
            .I(N__36193));
    InMux I__7537 (
            .O(N__36198),
            .I(N__36190));
    LocalMux I__7536 (
            .O(N__36193),
            .I(N__36187));
    LocalMux I__7535 (
            .O(N__36190),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    Odrv4 I__7534 (
            .O(N__36187),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    InMux I__7533 (
            .O(N__36182),
            .I(\current_shift_inst.timer_s1.counter_cry_19 ));
    InMux I__7532 (
            .O(N__36179),
            .I(N__36172));
    InMux I__7531 (
            .O(N__36178),
            .I(N__36172));
    InMux I__7530 (
            .O(N__36177),
            .I(N__36169));
    LocalMux I__7529 (
            .O(N__36172),
            .I(N__36166));
    LocalMux I__7528 (
            .O(N__36169),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    Odrv12 I__7527 (
            .O(N__36166),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    InMux I__7526 (
            .O(N__36161),
            .I(\current_shift_inst.timer_s1.counter_cry_20 ));
    CascadeMux I__7525 (
            .O(N__36158),
            .I(N__36154));
    CascadeMux I__7524 (
            .O(N__36157),
            .I(N__36151));
    InMux I__7523 (
            .O(N__36154),
            .I(N__36145));
    InMux I__7522 (
            .O(N__36151),
            .I(N__36145));
    InMux I__7521 (
            .O(N__36150),
            .I(N__36142));
    LocalMux I__7520 (
            .O(N__36145),
            .I(N__36139));
    LocalMux I__7519 (
            .O(N__36142),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    Odrv12 I__7518 (
            .O(N__36139),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    InMux I__7517 (
            .O(N__36134),
            .I(\current_shift_inst.timer_s1.counter_cry_21 ));
    InMux I__7516 (
            .O(N__36131),
            .I(N__36124));
    InMux I__7515 (
            .O(N__36130),
            .I(N__36124));
    InMux I__7514 (
            .O(N__36129),
            .I(N__36121));
    LocalMux I__7513 (
            .O(N__36124),
            .I(N__36118));
    LocalMux I__7512 (
            .O(N__36121),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    Odrv12 I__7511 (
            .O(N__36118),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    InMux I__7510 (
            .O(N__36113),
            .I(\current_shift_inst.timer_s1.counter_cry_5 ));
    InMux I__7509 (
            .O(N__36110),
            .I(N__36103));
    InMux I__7508 (
            .O(N__36109),
            .I(N__36103));
    InMux I__7507 (
            .O(N__36108),
            .I(N__36100));
    LocalMux I__7506 (
            .O(N__36103),
            .I(N__36097));
    LocalMux I__7505 (
            .O(N__36100),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    Odrv12 I__7504 (
            .O(N__36097),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    InMux I__7503 (
            .O(N__36092),
            .I(\current_shift_inst.timer_s1.counter_cry_6 ));
    CascadeMux I__7502 (
            .O(N__36089),
            .I(N__36086));
    InMux I__7501 (
            .O(N__36086),
            .I(N__36083));
    LocalMux I__7500 (
            .O(N__36083),
            .I(N__36079));
    InMux I__7499 (
            .O(N__36082),
            .I(N__36075));
    Span4Mux_v I__7498 (
            .O(N__36079),
            .I(N__36072));
    InMux I__7497 (
            .O(N__36078),
            .I(N__36069));
    LocalMux I__7496 (
            .O(N__36075),
            .I(N__36064));
    Span4Mux_h I__7495 (
            .O(N__36072),
            .I(N__36064));
    LocalMux I__7494 (
            .O(N__36069),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    Odrv4 I__7493 (
            .O(N__36064),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    InMux I__7492 (
            .O(N__36059),
            .I(bfn_15_14_0_));
    CascadeMux I__7491 (
            .O(N__36056),
            .I(N__36052));
    InMux I__7490 (
            .O(N__36055),
            .I(N__36049));
    InMux I__7489 (
            .O(N__36052),
            .I(N__36046));
    LocalMux I__7488 (
            .O(N__36049),
            .I(N__36040));
    LocalMux I__7487 (
            .O(N__36046),
            .I(N__36040));
    InMux I__7486 (
            .O(N__36045),
            .I(N__36037));
    Span4Mux_v I__7485 (
            .O(N__36040),
            .I(N__36034));
    LocalMux I__7484 (
            .O(N__36037),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    Odrv4 I__7483 (
            .O(N__36034),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    InMux I__7482 (
            .O(N__36029),
            .I(\current_shift_inst.timer_s1.counter_cry_8 ));
    CascadeMux I__7481 (
            .O(N__36026),
            .I(N__36022));
    CascadeMux I__7480 (
            .O(N__36025),
            .I(N__36019));
    InMux I__7479 (
            .O(N__36022),
            .I(N__36013));
    InMux I__7478 (
            .O(N__36019),
            .I(N__36013));
    InMux I__7477 (
            .O(N__36018),
            .I(N__36010));
    LocalMux I__7476 (
            .O(N__36013),
            .I(N__36007));
    LocalMux I__7475 (
            .O(N__36010),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    Odrv4 I__7474 (
            .O(N__36007),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    InMux I__7473 (
            .O(N__36002),
            .I(\current_shift_inst.timer_s1.counter_cry_9 ));
    CascadeMux I__7472 (
            .O(N__35999),
            .I(N__35995));
    CascadeMux I__7471 (
            .O(N__35998),
            .I(N__35992));
    InMux I__7470 (
            .O(N__35995),
            .I(N__35986));
    InMux I__7469 (
            .O(N__35992),
            .I(N__35986));
    InMux I__7468 (
            .O(N__35991),
            .I(N__35983));
    LocalMux I__7467 (
            .O(N__35986),
            .I(N__35980));
    LocalMux I__7466 (
            .O(N__35983),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    Odrv12 I__7465 (
            .O(N__35980),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    InMux I__7464 (
            .O(N__35975),
            .I(\current_shift_inst.timer_s1.counter_cry_10 ));
    InMux I__7463 (
            .O(N__35972),
            .I(N__35965));
    InMux I__7462 (
            .O(N__35971),
            .I(N__35965));
    InMux I__7461 (
            .O(N__35970),
            .I(N__35962));
    LocalMux I__7460 (
            .O(N__35965),
            .I(N__35959));
    LocalMux I__7459 (
            .O(N__35962),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    Odrv12 I__7458 (
            .O(N__35959),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    InMux I__7457 (
            .O(N__35954),
            .I(\current_shift_inst.timer_s1.counter_cry_11 ));
    InMux I__7456 (
            .O(N__35951),
            .I(N__35944));
    InMux I__7455 (
            .O(N__35950),
            .I(N__35944));
    InMux I__7454 (
            .O(N__35949),
            .I(N__35941));
    LocalMux I__7453 (
            .O(N__35944),
            .I(N__35938));
    LocalMux I__7452 (
            .O(N__35941),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    Odrv4 I__7451 (
            .O(N__35938),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    InMux I__7450 (
            .O(N__35933),
            .I(\current_shift_inst.timer_s1.counter_cry_12 ));
    InMux I__7449 (
            .O(N__35930),
            .I(N__35926));
    InMux I__7448 (
            .O(N__35929),
            .I(N__35923));
    LocalMux I__7447 (
            .O(N__35926),
            .I(N__35920));
    LocalMux I__7446 (
            .O(N__35923),
            .I(N__35917));
    Span4Mux_v I__7445 (
            .O(N__35920),
            .I(N__35911));
    Span4Mux_h I__7444 (
            .O(N__35917),
            .I(N__35911));
    InMux I__7443 (
            .O(N__35916),
            .I(N__35908));
    Odrv4 I__7442 (
            .O(N__35911),
            .I(\delay_measurement_inst.hc_stateZ0Z_0 ));
    LocalMux I__7441 (
            .O(N__35908),
            .I(\delay_measurement_inst.hc_stateZ0Z_0 ));
    InMux I__7440 (
            .O(N__35903),
            .I(N__35900));
    LocalMux I__7439 (
            .O(N__35900),
            .I(N__35896));
    InMux I__7438 (
            .O(N__35899),
            .I(N__35893));
    Span4Mux_v I__7437 (
            .O(N__35896),
            .I(N__35888));
    LocalMux I__7436 (
            .O(N__35893),
            .I(N__35888));
    Span4Mux_v I__7435 (
            .O(N__35888),
            .I(N__35885));
    Odrv4 I__7434 (
            .O(N__35885),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    InMux I__7433 (
            .O(N__35882),
            .I(N__35878));
    InMux I__7432 (
            .O(N__35881),
            .I(N__35875));
    LocalMux I__7431 (
            .O(N__35878),
            .I(N__35872));
    LocalMux I__7430 (
            .O(N__35875),
            .I(N__35869));
    Span4Mux_v I__7429 (
            .O(N__35872),
            .I(N__35863));
    Span4Mux_v I__7428 (
            .O(N__35869),
            .I(N__35863));
    InMux I__7427 (
            .O(N__35868),
            .I(N__35860));
    Odrv4 I__7426 (
            .O(N__35863),
            .I(\delay_measurement_inst.prev_hc_sigZ0 ));
    LocalMux I__7425 (
            .O(N__35860),
            .I(\delay_measurement_inst.prev_hc_sigZ0 ));
    CascadeMux I__7424 (
            .O(N__35855),
            .I(N__35851));
    InMux I__7423 (
            .O(N__35854),
            .I(N__35847));
    InMux I__7422 (
            .O(N__35851),
            .I(N__35844));
    InMux I__7421 (
            .O(N__35850),
            .I(N__35841));
    LocalMux I__7420 (
            .O(N__35847),
            .I(N__35836));
    LocalMux I__7419 (
            .O(N__35844),
            .I(N__35836));
    LocalMux I__7418 (
            .O(N__35841),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    Odrv12 I__7417 (
            .O(N__35836),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    InMux I__7416 (
            .O(N__35831),
            .I(bfn_15_13_0_));
    CascadeMux I__7415 (
            .O(N__35828),
            .I(N__35824));
    InMux I__7414 (
            .O(N__35827),
            .I(N__35821));
    InMux I__7413 (
            .O(N__35824),
            .I(N__35817));
    LocalMux I__7412 (
            .O(N__35821),
            .I(N__35814));
    InMux I__7411 (
            .O(N__35820),
            .I(N__35811));
    LocalMux I__7410 (
            .O(N__35817),
            .I(N__35808));
    Odrv12 I__7409 (
            .O(N__35814),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    LocalMux I__7408 (
            .O(N__35811),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    Odrv4 I__7407 (
            .O(N__35808),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    InMux I__7406 (
            .O(N__35801),
            .I(\current_shift_inst.timer_s1.counter_cry_0 ));
    InMux I__7405 (
            .O(N__35798),
            .I(N__35791));
    InMux I__7404 (
            .O(N__35797),
            .I(N__35791));
    InMux I__7403 (
            .O(N__35796),
            .I(N__35788));
    LocalMux I__7402 (
            .O(N__35791),
            .I(N__35785));
    LocalMux I__7401 (
            .O(N__35788),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    Odrv4 I__7400 (
            .O(N__35785),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    InMux I__7399 (
            .O(N__35780),
            .I(\current_shift_inst.timer_s1.counter_cry_1 ));
    InMux I__7398 (
            .O(N__35777),
            .I(N__35770));
    InMux I__7397 (
            .O(N__35776),
            .I(N__35770));
    InMux I__7396 (
            .O(N__35775),
            .I(N__35767));
    LocalMux I__7395 (
            .O(N__35770),
            .I(N__35764));
    LocalMux I__7394 (
            .O(N__35767),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    Odrv4 I__7393 (
            .O(N__35764),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    InMux I__7392 (
            .O(N__35759),
            .I(\current_shift_inst.timer_s1.counter_cry_2 ));
    CascadeMux I__7391 (
            .O(N__35756),
            .I(N__35752));
    CascadeMux I__7390 (
            .O(N__35755),
            .I(N__35749));
    InMux I__7389 (
            .O(N__35752),
            .I(N__35744));
    InMux I__7388 (
            .O(N__35749),
            .I(N__35744));
    LocalMux I__7387 (
            .O(N__35744),
            .I(N__35740));
    InMux I__7386 (
            .O(N__35743),
            .I(N__35737));
    Span4Mux_h I__7385 (
            .O(N__35740),
            .I(N__35734));
    LocalMux I__7384 (
            .O(N__35737),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    Odrv4 I__7383 (
            .O(N__35734),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    InMux I__7382 (
            .O(N__35729),
            .I(\current_shift_inst.timer_s1.counter_cry_3 ));
    CascadeMux I__7381 (
            .O(N__35726),
            .I(N__35722));
    CascadeMux I__7380 (
            .O(N__35725),
            .I(N__35719));
    InMux I__7379 (
            .O(N__35722),
            .I(N__35713));
    InMux I__7378 (
            .O(N__35719),
            .I(N__35713));
    InMux I__7377 (
            .O(N__35718),
            .I(N__35710));
    LocalMux I__7376 (
            .O(N__35713),
            .I(N__35707));
    LocalMux I__7375 (
            .O(N__35710),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    Odrv12 I__7374 (
            .O(N__35707),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    InMux I__7373 (
            .O(N__35702),
            .I(\current_shift_inst.timer_s1.counter_cry_4 ));
    CEMux I__7372 (
            .O(N__35699),
            .I(N__35684));
    CEMux I__7371 (
            .O(N__35698),
            .I(N__35684));
    CEMux I__7370 (
            .O(N__35697),
            .I(N__35684));
    CEMux I__7369 (
            .O(N__35696),
            .I(N__35684));
    CEMux I__7368 (
            .O(N__35695),
            .I(N__35684));
    GlobalMux I__7367 (
            .O(N__35684),
            .I(N__35681));
    gio2CtrlBuf I__7366 (
            .O(N__35681),
            .I(\delay_measurement_inst.delay_hc_timer.N_321_i_g ));
    InMux I__7365 (
            .O(N__35678),
            .I(N__35674));
    CascadeMux I__7364 (
            .O(N__35677),
            .I(N__35671));
    LocalMux I__7363 (
            .O(N__35674),
            .I(N__35667));
    InMux I__7362 (
            .O(N__35671),
            .I(N__35664));
    InMux I__7361 (
            .O(N__35670),
            .I(N__35661));
    Span4Mux_h I__7360 (
            .O(N__35667),
            .I(N__35658));
    LocalMux I__7359 (
            .O(N__35664),
            .I(N__35651));
    LocalMux I__7358 (
            .O(N__35661),
            .I(N__35651));
    Span4Mux_h I__7357 (
            .O(N__35658),
            .I(N__35648));
    InMux I__7356 (
            .O(N__35657),
            .I(N__35645));
    InMux I__7355 (
            .O(N__35656),
            .I(N__35642));
    Odrv12 I__7354 (
            .O(N__35651),
            .I(measured_delay_hc_10));
    Odrv4 I__7353 (
            .O(N__35648),
            .I(measured_delay_hc_10));
    LocalMux I__7352 (
            .O(N__35645),
            .I(measured_delay_hc_10));
    LocalMux I__7351 (
            .O(N__35642),
            .I(measured_delay_hc_10));
    InMux I__7350 (
            .O(N__35633),
            .I(N__35630));
    LocalMux I__7349 (
            .O(N__35630),
            .I(N__35627));
    Odrv4 I__7348 (
            .O(N__35627),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7 ));
    InMux I__7347 (
            .O(N__35624),
            .I(N__35621));
    LocalMux I__7346 (
            .O(N__35621),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    InMux I__7345 (
            .O(N__35618),
            .I(N__35615));
    LocalMux I__7344 (
            .O(N__35615),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    CascadeMux I__7343 (
            .O(N__35612),
            .I(N__35609));
    InMux I__7342 (
            .O(N__35609),
            .I(N__35606));
    LocalMux I__7341 (
            .O(N__35606),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    InMux I__7340 (
            .O(N__35603),
            .I(N__35600));
    LocalMux I__7339 (
            .O(N__35600),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    InMux I__7338 (
            .O(N__35597),
            .I(N__35594));
    LocalMux I__7337 (
            .O(N__35594),
            .I(N__35589));
    InMux I__7336 (
            .O(N__35593),
            .I(N__35584));
    InMux I__7335 (
            .O(N__35592),
            .I(N__35584));
    Span4Mux_h I__7334 (
            .O(N__35589),
            .I(N__35579));
    LocalMux I__7333 (
            .O(N__35584),
            .I(N__35579));
    Odrv4 I__7332 (
            .O(N__35579),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9 ));
    InMux I__7331 (
            .O(N__35576),
            .I(N__35573));
    LocalMux I__7330 (
            .O(N__35573),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2 ));
    InMux I__7329 (
            .O(N__35570),
            .I(N__35566));
    InMux I__7328 (
            .O(N__35569),
            .I(N__35563));
    LocalMux I__7327 (
            .O(N__35566),
            .I(N__35560));
    LocalMux I__7326 (
            .O(N__35563),
            .I(N__35553));
    Span4Mux_v I__7325 (
            .O(N__35560),
            .I(N__35553));
    InMux I__7324 (
            .O(N__35559),
            .I(N__35548));
    InMux I__7323 (
            .O(N__35558),
            .I(N__35548));
    Odrv4 I__7322 (
            .O(N__35553),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    LocalMux I__7321 (
            .O(N__35548),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    InMux I__7320 (
            .O(N__35543),
            .I(N__35540));
    LocalMux I__7319 (
            .O(N__35540),
            .I(N__35535));
    InMux I__7318 (
            .O(N__35539),
            .I(N__35532));
    InMux I__7317 (
            .O(N__35538),
            .I(N__35529));
    Odrv12 I__7316 (
            .O(N__35535),
            .I(\delay_measurement_inst.elapsed_time_hc_3 ));
    LocalMux I__7315 (
            .O(N__35532),
            .I(\delay_measurement_inst.elapsed_time_hc_3 ));
    LocalMux I__7314 (
            .O(N__35529),
            .I(\delay_measurement_inst.elapsed_time_hc_3 ));
    InMux I__7313 (
            .O(N__35522),
            .I(N__35519));
    LocalMux I__7312 (
            .O(N__35519),
            .I(N__35514));
    CascadeMux I__7311 (
            .O(N__35518),
            .I(N__35510));
    CascadeMux I__7310 (
            .O(N__35517),
            .I(N__35507));
    Span4Mux_v I__7309 (
            .O(N__35514),
            .I(N__35504));
    InMux I__7308 (
            .O(N__35513),
            .I(N__35501));
    InMux I__7307 (
            .O(N__35510),
            .I(N__35497));
    InMux I__7306 (
            .O(N__35507),
            .I(N__35494));
    Span4Mux_h I__7305 (
            .O(N__35504),
            .I(N__35491));
    LocalMux I__7304 (
            .O(N__35501),
            .I(N__35488));
    CascadeMux I__7303 (
            .O(N__35500),
            .I(N__35485));
    LocalMux I__7302 (
            .O(N__35497),
            .I(N__35482));
    LocalMux I__7301 (
            .O(N__35494),
            .I(N__35479));
    Span4Mux_h I__7300 (
            .O(N__35491),
            .I(N__35474));
    Span4Mux_v I__7299 (
            .O(N__35488),
            .I(N__35474));
    InMux I__7298 (
            .O(N__35485),
            .I(N__35471));
    Sp12to4 I__7297 (
            .O(N__35482),
            .I(N__35468));
    Span4Mux_h I__7296 (
            .O(N__35479),
            .I(N__35465));
    Span4Mux_h I__7295 (
            .O(N__35474),
            .I(N__35462));
    LocalMux I__7294 (
            .O(N__35471),
            .I(measured_delay_hc_3));
    Odrv12 I__7293 (
            .O(N__35468),
            .I(measured_delay_hc_3));
    Odrv4 I__7292 (
            .O(N__35465),
            .I(measured_delay_hc_3));
    Odrv4 I__7291 (
            .O(N__35462),
            .I(measured_delay_hc_3));
    InMux I__7290 (
            .O(N__35453),
            .I(N__35450));
    LocalMux I__7289 (
            .O(N__35450),
            .I(N__35445));
    InMux I__7288 (
            .O(N__35449),
            .I(N__35442));
    InMux I__7287 (
            .O(N__35448),
            .I(N__35439));
    Odrv12 I__7286 (
            .O(N__35445),
            .I(\delay_measurement_inst.elapsed_time_hc_4 ));
    LocalMux I__7285 (
            .O(N__35442),
            .I(\delay_measurement_inst.elapsed_time_hc_4 ));
    LocalMux I__7284 (
            .O(N__35439),
            .I(\delay_measurement_inst.elapsed_time_hc_4 ));
    InMux I__7283 (
            .O(N__35432),
            .I(N__35428));
    InMux I__7282 (
            .O(N__35431),
            .I(N__35423));
    LocalMux I__7281 (
            .O(N__35428),
            .I(N__35419));
    InMux I__7280 (
            .O(N__35427),
            .I(N__35416));
    InMux I__7279 (
            .O(N__35426),
            .I(N__35413));
    LocalMux I__7278 (
            .O(N__35423),
            .I(N__35410));
    CascadeMux I__7277 (
            .O(N__35422),
            .I(N__35407));
    Span4Mux_v I__7276 (
            .O(N__35419),
            .I(N__35404));
    LocalMux I__7275 (
            .O(N__35416),
            .I(N__35401));
    LocalMux I__7274 (
            .O(N__35413),
            .I(N__35398));
    Span4Mux_v I__7273 (
            .O(N__35410),
            .I(N__35395));
    InMux I__7272 (
            .O(N__35407),
            .I(N__35392));
    Span4Mux_h I__7271 (
            .O(N__35404),
            .I(N__35389));
    Sp12to4 I__7270 (
            .O(N__35401),
            .I(N__35386));
    Span4Mux_h I__7269 (
            .O(N__35398),
            .I(N__35383));
    Span4Mux_h I__7268 (
            .O(N__35395),
            .I(N__35380));
    LocalMux I__7267 (
            .O(N__35392),
            .I(measured_delay_hc_4));
    Odrv4 I__7266 (
            .O(N__35389),
            .I(measured_delay_hc_4));
    Odrv12 I__7265 (
            .O(N__35386),
            .I(measured_delay_hc_4));
    Odrv4 I__7264 (
            .O(N__35383),
            .I(measured_delay_hc_4));
    Odrv4 I__7263 (
            .O(N__35380),
            .I(measured_delay_hc_4));
    InMux I__7262 (
            .O(N__35369),
            .I(N__35366));
    LocalMux I__7261 (
            .O(N__35366),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    InMux I__7260 (
            .O(N__35363),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ));
    InMux I__7259 (
            .O(N__35360),
            .I(N__35357));
    LocalMux I__7258 (
            .O(N__35357),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    InMux I__7257 (
            .O(N__35354),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ));
    InMux I__7256 (
            .O(N__35351),
            .I(N__35348));
    LocalMux I__7255 (
            .O(N__35348),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    InMux I__7254 (
            .O(N__35345),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__7253 (
            .O(N__35342),
            .I(N__35339));
    InMux I__7252 (
            .O(N__35339),
            .I(N__35336));
    LocalMux I__7251 (
            .O(N__35336),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    InMux I__7250 (
            .O(N__35333),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ));
    InMux I__7249 (
            .O(N__35330),
            .I(bfn_15_10_0_));
    InMux I__7248 (
            .O(N__35327),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__7247 (
            .O(N__35324),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__7246 (
            .O(N__35321),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__7245 (
            .O(N__35318),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ));
    InMux I__7244 (
            .O(N__35315),
            .I(N__35306));
    InMux I__7243 (
            .O(N__35314),
            .I(N__35306));
    InMux I__7242 (
            .O(N__35313),
            .I(N__35306));
    LocalMux I__7241 (
            .O(N__35306),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    InMux I__7240 (
            .O(N__35303),
            .I(N__35299));
    InMux I__7239 (
            .O(N__35302),
            .I(N__35295));
    LocalMux I__7238 (
            .O(N__35299),
            .I(N__35292));
    InMux I__7237 (
            .O(N__35298),
            .I(N__35289));
    LocalMux I__7236 (
            .O(N__35295),
            .I(N__35285));
    Span4Mux_h I__7235 (
            .O(N__35292),
            .I(N__35280));
    LocalMux I__7234 (
            .O(N__35289),
            .I(N__35280));
    InMux I__7233 (
            .O(N__35288),
            .I(N__35277));
    Odrv4 I__7232 (
            .O(N__35285),
            .I(\delay_measurement_inst.delay_hc_reg3lto14 ));
    Odrv4 I__7231 (
            .O(N__35280),
            .I(\delay_measurement_inst.delay_hc_reg3lto14 ));
    LocalMux I__7230 (
            .O(N__35277),
            .I(\delay_measurement_inst.delay_hc_reg3lto14 ));
    InMux I__7229 (
            .O(N__35270),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ));
    CascadeMux I__7228 (
            .O(N__35267),
            .I(N__35264));
    InMux I__7227 (
            .O(N__35264),
            .I(N__35261));
    LocalMux I__7226 (
            .O(N__35261),
            .I(N__35253));
    InMux I__7225 (
            .O(N__35260),
            .I(N__35250));
    InMux I__7224 (
            .O(N__35259),
            .I(N__35246));
    InMux I__7223 (
            .O(N__35258),
            .I(N__35243));
    InMux I__7222 (
            .O(N__35257),
            .I(N__35240));
    InMux I__7221 (
            .O(N__35256),
            .I(N__35237));
    Span4Mux_h I__7220 (
            .O(N__35253),
            .I(N__35232));
    LocalMux I__7219 (
            .O(N__35250),
            .I(N__35232));
    InMux I__7218 (
            .O(N__35249),
            .I(N__35229));
    LocalMux I__7217 (
            .O(N__35246),
            .I(N__35224));
    LocalMux I__7216 (
            .O(N__35243),
            .I(N__35224));
    LocalMux I__7215 (
            .O(N__35240),
            .I(\delay_measurement_inst.delay_hc_reg3lto15 ));
    LocalMux I__7214 (
            .O(N__35237),
            .I(\delay_measurement_inst.delay_hc_reg3lto15 ));
    Odrv4 I__7213 (
            .O(N__35232),
            .I(\delay_measurement_inst.delay_hc_reg3lto15 ));
    LocalMux I__7212 (
            .O(N__35229),
            .I(\delay_measurement_inst.delay_hc_reg3lto15 ));
    Odrv4 I__7211 (
            .O(N__35224),
            .I(\delay_measurement_inst.delay_hc_reg3lto15 ));
    InMux I__7210 (
            .O(N__35213),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ));
    CascadeMux I__7209 (
            .O(N__35210),
            .I(N__35207));
    InMux I__7208 (
            .O(N__35207),
            .I(N__35203));
    InMux I__7207 (
            .O(N__35206),
            .I(N__35200));
    LocalMux I__7206 (
            .O(N__35203),
            .I(N__35195));
    LocalMux I__7205 (
            .O(N__35200),
            .I(N__35195));
    Span4Mux_v I__7204 (
            .O(N__35195),
            .I(N__35191));
    InMux I__7203 (
            .O(N__35194),
            .I(N__35188));
    Odrv4 I__7202 (
            .O(N__35191),
            .I(\delay_measurement_inst.elapsed_time_hc_16 ));
    LocalMux I__7201 (
            .O(N__35188),
            .I(\delay_measurement_inst.elapsed_time_hc_16 ));
    InMux I__7200 (
            .O(N__35183),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ));
    InMux I__7199 (
            .O(N__35180),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ));
    InMux I__7198 (
            .O(N__35177),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ));
    InMux I__7197 (
            .O(N__35174),
            .I(bfn_15_9_0_));
    CascadeMux I__7196 (
            .O(N__35171),
            .I(N__35167));
    InMux I__7195 (
            .O(N__35170),
            .I(N__35162));
    InMux I__7194 (
            .O(N__35167),
            .I(N__35162));
    LocalMux I__7193 (
            .O(N__35162),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    InMux I__7192 (
            .O(N__35159),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ));
    InMux I__7191 (
            .O(N__35156),
            .I(N__35150));
    InMux I__7190 (
            .O(N__35155),
            .I(N__35150));
    LocalMux I__7189 (
            .O(N__35150),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    InMux I__7188 (
            .O(N__35147),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__7187 (
            .O(N__35144),
            .I(N__35140));
    InMux I__7186 (
            .O(N__35143),
            .I(N__35137));
    LocalMux I__7185 (
            .O(N__35140),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    LocalMux I__7184 (
            .O(N__35137),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    InMux I__7183 (
            .O(N__35132),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ));
    InMux I__7182 (
            .O(N__35129),
            .I(N__35125));
    InMux I__7181 (
            .O(N__35128),
            .I(N__35121));
    LocalMux I__7180 (
            .O(N__35125),
            .I(N__35118));
    CascadeMux I__7179 (
            .O(N__35124),
            .I(N__35114));
    LocalMux I__7178 (
            .O(N__35121),
            .I(N__35111));
    Span4Mux_v I__7177 (
            .O(N__35118),
            .I(N__35108));
    InMux I__7176 (
            .O(N__35117),
            .I(N__35105));
    InMux I__7175 (
            .O(N__35114),
            .I(N__35102));
    Span4Mux_v I__7174 (
            .O(N__35111),
            .I(N__35099));
    Odrv4 I__7173 (
            .O(N__35108),
            .I(\delay_measurement_inst.delay_hc_reg3lto6 ));
    LocalMux I__7172 (
            .O(N__35105),
            .I(\delay_measurement_inst.delay_hc_reg3lto6 ));
    LocalMux I__7171 (
            .O(N__35102),
            .I(\delay_measurement_inst.delay_hc_reg3lto6 ));
    Odrv4 I__7170 (
            .O(N__35099),
            .I(\delay_measurement_inst.delay_hc_reg3lto6 ));
    InMux I__7169 (
            .O(N__35090),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ));
    InMux I__7168 (
            .O(N__35087),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ));
    InMux I__7167 (
            .O(N__35084),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ));
    InMux I__7166 (
            .O(N__35081),
            .I(N__35077));
    InMux I__7165 (
            .O(N__35080),
            .I(N__35072));
    LocalMux I__7164 (
            .O(N__35077),
            .I(N__35069));
    CascadeMux I__7163 (
            .O(N__35076),
            .I(N__35066));
    InMux I__7162 (
            .O(N__35075),
            .I(N__35063));
    LocalMux I__7161 (
            .O(N__35072),
            .I(N__35060));
    Span4Mux_h I__7160 (
            .O(N__35069),
            .I(N__35057));
    InMux I__7159 (
            .O(N__35066),
            .I(N__35054));
    LocalMux I__7158 (
            .O(N__35063),
            .I(N__35049));
    Span4Mux_h I__7157 (
            .O(N__35060),
            .I(N__35049));
    Odrv4 I__7156 (
            .O(N__35057),
            .I(\delay_measurement_inst.delay_hc_reg3lto9 ));
    LocalMux I__7155 (
            .O(N__35054),
            .I(\delay_measurement_inst.delay_hc_reg3lto9 ));
    Odrv4 I__7154 (
            .O(N__35049),
            .I(\delay_measurement_inst.delay_hc_reg3lto9 ));
    InMux I__7153 (
            .O(N__35042),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ));
    InMux I__7152 (
            .O(N__35039),
            .I(N__35035));
    CascadeMux I__7151 (
            .O(N__35038),
            .I(N__35032));
    LocalMux I__7150 (
            .O(N__35035),
            .I(N__35028));
    InMux I__7149 (
            .O(N__35032),
            .I(N__35025));
    InMux I__7148 (
            .O(N__35031),
            .I(N__35022));
    Odrv4 I__7147 (
            .O(N__35028),
            .I(\delay_measurement_inst.elapsed_time_hc_10 ));
    LocalMux I__7146 (
            .O(N__35025),
            .I(\delay_measurement_inst.elapsed_time_hc_10 ));
    LocalMux I__7145 (
            .O(N__35022),
            .I(\delay_measurement_inst.elapsed_time_hc_10 ));
    InMux I__7144 (
            .O(N__35015),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__7143 (
            .O(N__35012),
            .I(N__35008));
    InMux I__7142 (
            .O(N__35011),
            .I(N__35003));
    InMux I__7141 (
            .O(N__35008),
            .I(N__35003));
    LocalMux I__7140 (
            .O(N__35003),
            .I(N__34999));
    InMux I__7139 (
            .O(N__35002),
            .I(N__34996));
    Span4Mux_v I__7138 (
            .O(N__34999),
            .I(N__34991));
    LocalMux I__7137 (
            .O(N__34996),
            .I(N__34991));
    Odrv4 I__7136 (
            .O(N__34991),
            .I(\delay_measurement_inst.elapsed_time_hc_11 ));
    InMux I__7135 (
            .O(N__34988),
            .I(bfn_15_8_0_));
    InMux I__7134 (
            .O(N__34985),
            .I(N__34978));
    InMux I__7133 (
            .O(N__34984),
            .I(N__34978));
    CascadeMux I__7132 (
            .O(N__34983),
            .I(N__34975));
    LocalMux I__7131 (
            .O(N__34978),
            .I(N__34972));
    InMux I__7130 (
            .O(N__34975),
            .I(N__34969));
    Odrv4 I__7129 (
            .O(N__34972),
            .I(\delay_measurement_inst.elapsed_time_hc_12 ));
    LocalMux I__7128 (
            .O(N__34969),
            .I(\delay_measurement_inst.elapsed_time_hc_12 ));
    InMux I__7127 (
            .O(N__34964),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__7126 (
            .O(N__34961),
            .I(N__34957));
    InMux I__7125 (
            .O(N__34960),
            .I(N__34954));
    InMux I__7124 (
            .O(N__34957),
            .I(N__34951));
    LocalMux I__7123 (
            .O(N__34954),
            .I(N__34948));
    LocalMux I__7122 (
            .O(N__34951),
            .I(N__34944));
    Span4Mux_v I__7121 (
            .O(N__34948),
            .I(N__34941));
    InMux I__7120 (
            .O(N__34947),
            .I(N__34938));
    Span4Mux_h I__7119 (
            .O(N__34944),
            .I(N__34935));
    Odrv4 I__7118 (
            .O(N__34941),
            .I(\delay_measurement_inst.elapsed_time_hc_13 ));
    LocalMux I__7117 (
            .O(N__34938),
            .I(\delay_measurement_inst.elapsed_time_hc_13 ));
    Odrv4 I__7116 (
            .O(N__34935),
            .I(\delay_measurement_inst.elapsed_time_hc_13 ));
    InMux I__7115 (
            .O(N__34928),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ));
    InMux I__7114 (
            .O(N__34925),
            .I(N__34922));
    LocalMux I__7113 (
            .O(N__34922),
            .I(N__34919));
    Odrv12 I__7112 (
            .O(N__34919),
            .I(delay_tr_input_c));
    InMux I__7111 (
            .O(N__34916),
            .I(N__34913));
    LocalMux I__7110 (
            .O(N__34913),
            .I(delay_tr_d1));
    InMux I__7109 (
            .O(N__34910),
            .I(N__34907));
    LocalMux I__7108 (
            .O(N__34907),
            .I(N__34901));
    InMux I__7107 (
            .O(N__34906),
            .I(N__34894));
    InMux I__7106 (
            .O(N__34905),
            .I(N__34894));
    InMux I__7105 (
            .O(N__34904),
            .I(N__34894));
    Span4Mux_v I__7104 (
            .O(N__34901),
            .I(N__34891));
    LocalMux I__7103 (
            .O(N__34894),
            .I(N__34888));
    Span4Mux_h I__7102 (
            .O(N__34891),
            .I(N__34885));
    Span4Mux_v I__7101 (
            .O(N__34888),
            .I(N__34882));
    Span4Mux_v I__7100 (
            .O(N__34885),
            .I(N__34879));
    Span4Mux_v I__7099 (
            .O(N__34882),
            .I(N__34876));
    Odrv4 I__7098 (
            .O(N__34879),
            .I(delay_tr_d2));
    Odrv4 I__7097 (
            .O(N__34876),
            .I(delay_tr_d2));
    InMux I__7096 (
            .O(N__34871),
            .I(N__34868));
    LocalMux I__7095 (
            .O(N__34868),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_4 ));
    InMux I__7094 (
            .O(N__34865),
            .I(N__34862));
    LocalMux I__7093 (
            .O(N__34862),
            .I(N__34859));
    Span4Mux_v I__7092 (
            .O(N__34859),
            .I(N__34855));
    InMux I__7091 (
            .O(N__34858),
            .I(N__34852));
    Odrv4 I__7090 (
            .O(N__34855),
            .I(\delay_measurement_inst.elapsed_time_hc_1 ));
    LocalMux I__7089 (
            .O(N__34852),
            .I(\delay_measurement_inst.elapsed_time_hc_1 ));
    InMux I__7088 (
            .O(N__34847),
            .I(N__34844));
    LocalMux I__7087 (
            .O(N__34844),
            .I(N__34841));
    Span4Mux_h I__7086 (
            .O(N__34841),
            .I(N__34836));
    InMux I__7085 (
            .O(N__34840),
            .I(N__34833));
    InMux I__7084 (
            .O(N__34839),
            .I(N__34830));
    Odrv4 I__7083 (
            .O(N__34836),
            .I(\delay_measurement_inst.elapsed_time_hc_2 ));
    LocalMux I__7082 (
            .O(N__34833),
            .I(\delay_measurement_inst.elapsed_time_hc_2 ));
    LocalMux I__7081 (
            .O(N__34830),
            .I(\delay_measurement_inst.elapsed_time_hc_2 ));
    InMux I__7080 (
            .O(N__34823),
            .I(N__34820));
    LocalMux I__7079 (
            .O(N__34820),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6 ));
    InMux I__7078 (
            .O(N__34817),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ));
    InMux I__7077 (
            .O(N__34814),
            .I(N__34810));
    CascadeMux I__7076 (
            .O(N__34813),
            .I(N__34807));
    LocalMux I__7075 (
            .O(N__34810),
            .I(N__34804));
    InMux I__7074 (
            .O(N__34807),
            .I(N__34800));
    Span4Mux_v I__7073 (
            .O(N__34804),
            .I(N__34797));
    InMux I__7072 (
            .O(N__34803),
            .I(N__34794));
    LocalMux I__7071 (
            .O(N__34800),
            .I(N__34791));
    Odrv4 I__7070 (
            .O(N__34797),
            .I(\delay_measurement_inst.elapsed_time_hc_5 ));
    LocalMux I__7069 (
            .O(N__34794),
            .I(\delay_measurement_inst.elapsed_time_hc_5 ));
    Odrv4 I__7068 (
            .O(N__34791),
            .I(\delay_measurement_inst.elapsed_time_hc_5 ));
    InMux I__7067 (
            .O(N__34784),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ));
    InMux I__7066 (
            .O(N__34781),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12 ));
    InMux I__7065 (
            .O(N__34778),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13 ));
    InMux I__7064 (
            .O(N__34775),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14 ));
    InMux I__7063 (
            .O(N__34772),
            .I(bfn_14_24_0_));
    InMux I__7062 (
            .O(N__34769),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16 ));
    InMux I__7061 (
            .O(N__34766),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17 ));
    InMux I__7060 (
            .O(N__34763),
            .I(N__34760));
    LocalMux I__7059 (
            .O(N__34760),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13 ));
    InMux I__7058 (
            .O(N__34757),
            .I(N__34754));
    LocalMux I__7057 (
            .O(N__34754),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17 ));
    InMux I__7056 (
            .O(N__34751),
            .I(N__34748));
    LocalMux I__7055 (
            .O(N__34748),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18 ));
    InMux I__7054 (
            .O(N__34745),
            .I(N__34742));
    LocalMux I__7053 (
            .O(N__34742),
            .I(N__34739));
    Span4Mux_v I__7052 (
            .O(N__34739),
            .I(N__34736));
    Odrv4 I__7051 (
            .O(N__34736),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5 ));
    InMux I__7050 (
            .O(N__34733),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3 ));
    InMux I__7049 (
            .O(N__34730),
            .I(N__34727));
    LocalMux I__7048 (
            .O(N__34727),
            .I(N__34723));
    InMux I__7047 (
            .O(N__34726),
            .I(N__34720));
    Odrv4 I__7046 (
            .O(N__34723),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6 ));
    LocalMux I__7045 (
            .O(N__34720),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__7044 (
            .O(N__34715),
            .I(N__34712));
    LocalMux I__7043 (
            .O(N__34712),
            .I(N__34709));
    Odrv4 I__7042 (
            .O(N__34709),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6 ));
    InMux I__7041 (
            .O(N__34706),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4 ));
    InMux I__7040 (
            .O(N__34703),
            .I(N__34700));
    LocalMux I__7039 (
            .O(N__34700),
            .I(N__34696));
    InMux I__7038 (
            .O(N__34699),
            .I(N__34693));
    Odrv4 I__7037 (
            .O(N__34696),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7 ));
    LocalMux I__7036 (
            .O(N__34693),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__7035 (
            .O(N__34688),
            .I(N__34685));
    LocalMux I__7034 (
            .O(N__34685),
            .I(N__34682));
    Span4Mux_v I__7033 (
            .O(N__34682),
            .I(N__34679));
    Span4Mux_h I__7032 (
            .O(N__34679),
            .I(N__34676));
    Odrv4 I__7031 (
            .O(N__34676),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7 ));
    InMux I__7030 (
            .O(N__34673),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5 ));
    InMux I__7029 (
            .O(N__34670),
            .I(N__34667));
    LocalMux I__7028 (
            .O(N__34667),
            .I(N__34663));
    InMux I__7027 (
            .O(N__34666),
            .I(N__34660));
    Odrv4 I__7026 (
            .O(N__34663),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8 ));
    LocalMux I__7025 (
            .O(N__34660),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8 ));
    CascadeMux I__7024 (
            .O(N__34655),
            .I(N__34652));
    InMux I__7023 (
            .O(N__34652),
            .I(N__34649));
    LocalMux I__7022 (
            .O(N__34649),
            .I(N__34646));
    Odrv12 I__7021 (
            .O(N__34646),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8 ));
    InMux I__7020 (
            .O(N__34643),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6 ));
    InMux I__7019 (
            .O(N__34640),
            .I(bfn_14_23_0_));
    InMux I__7018 (
            .O(N__34637),
            .I(N__34633));
    InMux I__7017 (
            .O(N__34636),
            .I(N__34630));
    LocalMux I__7016 (
            .O(N__34633),
            .I(N__34627));
    LocalMux I__7015 (
            .O(N__34630),
            .I(N__34624));
    Odrv12 I__7014 (
            .O(N__34627),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10 ));
    Odrv4 I__7013 (
            .O(N__34624),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__7012 (
            .O(N__34619),
            .I(N__34616));
    LocalMux I__7011 (
            .O(N__34616),
            .I(N__34613));
    Odrv12 I__7010 (
            .O(N__34613),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10 ));
    InMux I__7009 (
            .O(N__34610),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8 ));
    InMux I__7008 (
            .O(N__34607),
            .I(N__34603));
    InMux I__7007 (
            .O(N__34606),
            .I(N__34600));
    LocalMux I__7006 (
            .O(N__34603),
            .I(N__34597));
    LocalMux I__7005 (
            .O(N__34600),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11 ));
    Odrv4 I__7004 (
            .O(N__34597),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__7003 (
            .O(N__34592),
            .I(N__34589));
    LocalMux I__7002 (
            .O(N__34589),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11 ));
    InMux I__7001 (
            .O(N__34586),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9 ));
    InMux I__7000 (
            .O(N__34583),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10 ));
    InMux I__6999 (
            .O(N__34580),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11 ));
    InMux I__6998 (
            .O(N__34577),
            .I(N__34574));
    LocalMux I__6997 (
            .O(N__34574),
            .I(N__34571));
    Odrv4 I__6996 (
            .O(N__34571),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0 ));
    InMux I__6995 (
            .O(N__34568),
            .I(N__34565));
    LocalMux I__6994 (
            .O(N__34565),
            .I(N__34561));
    InMux I__6993 (
            .O(N__34564),
            .I(N__34558));
    Span4Mux_s1_v I__6992 (
            .O(N__34561),
            .I(N__34552));
    LocalMux I__6991 (
            .O(N__34558),
            .I(N__34552));
    InMux I__6990 (
            .O(N__34557),
            .I(N__34549));
    Span4Mux_v I__6989 (
            .O(N__34552),
            .I(N__34546));
    LocalMux I__6988 (
            .O(N__34549),
            .I(N__34541));
    Span4Mux_h I__6987 (
            .O(N__34546),
            .I(N__34538));
    InMux I__6986 (
            .O(N__34545),
            .I(N__34531));
    InMux I__6985 (
            .O(N__34544),
            .I(N__34531));
    Span4Mux_v I__6984 (
            .O(N__34541),
            .I(N__34528));
    Sp12to4 I__6983 (
            .O(N__34538),
            .I(N__34525));
    InMux I__6982 (
            .O(N__34537),
            .I(N__34522));
    CascadeMux I__6981 (
            .O(N__34536),
            .I(N__34519));
    LocalMux I__6980 (
            .O(N__34531),
            .I(N__34516));
    Span4Mux_h I__6979 (
            .O(N__34528),
            .I(N__34513));
    Span12Mux_s11_v I__6978 (
            .O(N__34525),
            .I(N__34510));
    LocalMux I__6977 (
            .O(N__34522),
            .I(N__34507));
    InMux I__6976 (
            .O(N__34519),
            .I(N__34504));
    Span4Mux_v I__6975 (
            .O(N__34516),
            .I(N__34501));
    Sp12to4 I__6974 (
            .O(N__34513),
            .I(N__34498));
    Span12Mux_v I__6973 (
            .O(N__34510),
            .I(N__34491));
    Sp12to4 I__6972 (
            .O(N__34507),
            .I(N__34491));
    LocalMux I__6971 (
            .O(N__34504),
            .I(N__34491));
    Span4Mux_h I__6970 (
            .O(N__34501),
            .I(N__34488));
    Span12Mux_v I__6969 (
            .O(N__34498),
            .I(N__34483));
    Span12Mux_h I__6968 (
            .O(N__34491),
            .I(N__34483));
    Span4Mux_v I__6967 (
            .O(N__34488),
            .I(N__34480));
    Odrv12 I__6966 (
            .O(N__34483),
            .I(start_stop_c));
    Odrv4 I__6965 (
            .O(N__34480),
            .I(start_stop_c));
    InMux I__6964 (
            .O(N__34475),
            .I(N__34471));
    CascadeMux I__6963 (
            .O(N__34474),
            .I(N__34468));
    LocalMux I__6962 (
            .O(N__34471),
            .I(N__34465));
    InMux I__6961 (
            .O(N__34468),
            .I(N__34462));
    Span12Mux_s10_v I__6960 (
            .O(N__34465),
            .I(N__34459));
    LocalMux I__6959 (
            .O(N__34462),
            .I(shift_flag_start));
    Odrv12 I__6958 (
            .O(N__34459),
            .I(shift_flag_start));
    InMux I__6957 (
            .O(N__34454),
            .I(N__34448));
    InMux I__6956 (
            .O(N__34453),
            .I(N__34448));
    LocalMux I__6955 (
            .O(N__34448),
            .I(N__34445));
    Span4Mux_v I__6954 (
            .O(N__34445),
            .I(N__34442));
    Odrv4 I__6953 (
            .O(N__34442),
            .I(\phase_controller_slave.un1_startZ0 ));
    InMux I__6952 (
            .O(N__34439),
            .I(N__34436));
    LocalMux I__6951 (
            .O(N__34436),
            .I(N__34433));
    Span4Mux_h I__6950 (
            .O(N__34433),
            .I(N__34428));
    InMux I__6949 (
            .O(N__34432),
            .I(N__34423));
    InMux I__6948 (
            .O(N__34431),
            .I(N__34423));
    Odrv4 I__6947 (
            .O(N__34428),
            .I(\phase_controller_slave.stoper_tr.time_passed11 ));
    LocalMux I__6946 (
            .O(N__34423),
            .I(\phase_controller_slave.stoper_tr.time_passed11 ));
    InMux I__6945 (
            .O(N__34418),
            .I(N__34412));
    InMux I__6944 (
            .O(N__34417),
            .I(N__34412));
    LocalMux I__6943 (
            .O(N__34412),
            .I(N__34407));
    InMux I__6942 (
            .O(N__34411),
            .I(N__34404));
    InMux I__6941 (
            .O(N__34410),
            .I(N__34399));
    Span4Mux_v I__6940 (
            .O(N__34407),
            .I(N__34396));
    LocalMux I__6939 (
            .O(N__34404),
            .I(N__34393));
    InMux I__6938 (
            .O(N__34403),
            .I(N__34388));
    InMux I__6937 (
            .O(N__34402),
            .I(N__34388));
    LocalMux I__6936 (
            .O(N__34399),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__6935 (
            .O(N__34396),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__6934 (
            .O(N__34393),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__6933 (
            .O(N__34388),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    InMux I__6932 (
            .O(N__34379),
            .I(N__34376));
    LocalMux I__6931 (
            .O(N__34376),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2 ));
    CascadeMux I__6930 (
            .O(N__34373),
            .I(N__34370));
    InMux I__6929 (
            .O(N__34370),
            .I(N__34366));
    InMux I__6928 (
            .O(N__34369),
            .I(N__34362));
    LocalMux I__6927 (
            .O(N__34366),
            .I(N__34359));
    InMux I__6926 (
            .O(N__34365),
            .I(N__34356));
    LocalMux I__6925 (
            .O(N__34362),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv12 I__6924 (
            .O(N__34359),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__6923 (
            .O(N__34356),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ));
    InMux I__6922 (
            .O(N__34349),
            .I(N__34346));
    LocalMux I__6921 (
            .O(N__34346),
            .I(N__34342));
    InMux I__6920 (
            .O(N__34345),
            .I(N__34339));
    Odrv12 I__6919 (
            .O(N__34342),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2 ));
    LocalMux I__6918 (
            .O(N__34339),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__6917 (
            .O(N__34334),
            .I(N__34331));
    LocalMux I__6916 (
            .O(N__34331),
            .I(N__34328));
    Odrv4 I__6915 (
            .O(N__34328),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2 ));
    InMux I__6914 (
            .O(N__34325),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0 ));
    InMux I__6913 (
            .O(N__34322),
            .I(N__34319));
    LocalMux I__6912 (
            .O(N__34319),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6 ));
    CascadeMux I__6911 (
            .O(N__34316),
            .I(N__34313));
    InMux I__6910 (
            .O(N__34313),
            .I(N__34310));
    LocalMux I__6909 (
            .O(N__34310),
            .I(N__34306));
    InMux I__6908 (
            .O(N__34309),
            .I(N__34303));
    Odrv12 I__6907 (
            .O(N__34306),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3 ));
    LocalMux I__6906 (
            .O(N__34303),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__6905 (
            .O(N__34298),
            .I(N__34295));
    LocalMux I__6904 (
            .O(N__34295),
            .I(N__34292));
    Span4Mux_v I__6903 (
            .O(N__34292),
            .I(N__34289));
    Odrv4 I__6902 (
            .O(N__34289),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3 ));
    InMux I__6901 (
            .O(N__34286),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1 ));
    InMux I__6900 (
            .O(N__34283),
            .I(N__34280));
    LocalMux I__6899 (
            .O(N__34280),
            .I(N__34276));
    InMux I__6898 (
            .O(N__34279),
            .I(N__34273));
    Odrv4 I__6897 (
            .O(N__34276),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4 ));
    LocalMux I__6896 (
            .O(N__34273),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4 ));
    CascadeMux I__6895 (
            .O(N__34268),
            .I(N__34265));
    InMux I__6894 (
            .O(N__34265),
            .I(N__34262));
    LocalMux I__6893 (
            .O(N__34262),
            .I(N__34259));
    Odrv4 I__6892 (
            .O(N__34259),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4 ));
    InMux I__6891 (
            .O(N__34256),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2 ));
    InMux I__6890 (
            .O(N__34253),
            .I(N__34250));
    LocalMux I__6889 (
            .O(N__34250),
            .I(N__34246));
    InMux I__6888 (
            .O(N__34249),
            .I(N__34243));
    Odrv4 I__6887 (
            .O(N__34246),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5 ));
    LocalMux I__6886 (
            .O(N__34243),
            .I(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__6885 (
            .O(N__34238),
            .I(N__34235));
    LocalMux I__6884 (
            .O(N__34235),
            .I(N__34232));
    Span4Mux_h I__6883 (
            .O(N__34232),
            .I(N__34229));
    Odrv4 I__6882 (
            .O(N__34229),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3 ));
    CascadeMux I__6881 (
            .O(N__34226),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3Z0Z_3_cascade_ ));
    InMux I__6880 (
            .O(N__34223),
            .I(N__34220));
    LocalMux I__6879 (
            .O(N__34220),
            .I(N__34217));
    Span4Mux_h I__6878 (
            .O(N__34217),
            .I(N__34214));
    Odrv4 I__6877 (
            .O(N__34214),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_5Z0Z_3 ));
    CascadeMux I__6876 (
            .O(N__34211),
            .I(\phase_controller_slave.stoper_hc.time_passed11_cascade_ ));
    InMux I__6875 (
            .O(N__34208),
            .I(N__34205));
    LocalMux I__6874 (
            .O(N__34205),
            .I(N__34202));
    Odrv4 I__6873 (
            .O(N__34202),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1 ));
    InMux I__6872 (
            .O(N__34199),
            .I(N__34196));
    LocalMux I__6871 (
            .O(N__34196),
            .I(N__34193));
    Span4Mux_v I__6870 (
            .O(N__34193),
            .I(N__34190));
    Odrv4 I__6869 (
            .O(N__34190),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8 ));
    CascadeMux I__6868 (
            .O(N__34187),
            .I(N__34184));
    InMux I__6867 (
            .O(N__34184),
            .I(N__34181));
    LocalMux I__6866 (
            .O(N__34181),
            .I(N__34178));
    Span4Mux_h I__6865 (
            .O(N__34178),
            .I(N__34175));
    Odrv4 I__6864 (
            .O(N__34175),
            .I(\phase_controller_slave.stoper_hc.time_passed_1_sqmuxa ));
    CascadeMux I__6863 (
            .O(N__34172),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ));
    InMux I__6862 (
            .O(N__34169),
            .I(N__34166));
    LocalMux I__6861 (
            .O(N__34166),
            .I(N__34162));
    InMux I__6860 (
            .O(N__34165),
            .I(N__34159));
    Span4Mux_v I__6859 (
            .O(N__34162),
            .I(N__34155));
    LocalMux I__6858 (
            .O(N__34159),
            .I(N__34152));
    CascadeMux I__6857 (
            .O(N__34158),
            .I(N__34147));
    Span4Mux_h I__6856 (
            .O(N__34155),
            .I(N__34144));
    Span4Mux_v I__6855 (
            .O(N__34152),
            .I(N__34141));
    InMux I__6854 (
            .O(N__34151),
            .I(N__34138));
    InMux I__6853 (
            .O(N__34150),
            .I(N__34135));
    InMux I__6852 (
            .O(N__34147),
            .I(N__34132));
    Span4Mux_h I__6851 (
            .O(N__34144),
            .I(N__34125));
    Span4Mux_v I__6850 (
            .O(N__34141),
            .I(N__34125));
    LocalMux I__6849 (
            .O(N__34138),
            .I(N__34125));
    LocalMux I__6848 (
            .O(N__34135),
            .I(N__34122));
    LocalMux I__6847 (
            .O(N__34132),
            .I(measured_delay_hc_6));
    Odrv4 I__6846 (
            .O(N__34125),
            .I(measured_delay_hc_6));
    Odrv4 I__6845 (
            .O(N__34122),
            .I(measured_delay_hc_6));
    InMux I__6844 (
            .O(N__34115),
            .I(N__34111));
    CascadeMux I__6843 (
            .O(N__34114),
            .I(N__34108));
    LocalMux I__6842 (
            .O(N__34111),
            .I(N__34103));
    InMux I__6841 (
            .O(N__34108),
            .I(N__34100));
    InMux I__6840 (
            .O(N__34107),
            .I(N__34096));
    CascadeMux I__6839 (
            .O(N__34106),
            .I(N__34093));
    Span4Mux_v I__6838 (
            .O(N__34103),
            .I(N__34090));
    LocalMux I__6837 (
            .O(N__34100),
            .I(N__34087));
    InMux I__6836 (
            .O(N__34099),
            .I(N__34084));
    LocalMux I__6835 (
            .O(N__34096),
            .I(N__34081));
    InMux I__6834 (
            .O(N__34093),
            .I(N__34078));
    Span4Mux_v I__6833 (
            .O(N__34090),
            .I(N__34075));
    Span12Mux_h I__6832 (
            .O(N__34087),
            .I(N__34072));
    LocalMux I__6831 (
            .O(N__34084),
            .I(N__34069));
    Span4Mux_v I__6830 (
            .O(N__34081),
            .I(N__34066));
    LocalMux I__6829 (
            .O(N__34078),
            .I(measured_delay_hc_2));
    Odrv4 I__6828 (
            .O(N__34075),
            .I(measured_delay_hc_2));
    Odrv12 I__6827 (
            .O(N__34072),
            .I(measured_delay_hc_2));
    Odrv4 I__6826 (
            .O(N__34069),
            .I(measured_delay_hc_2));
    Odrv4 I__6825 (
            .O(N__34066),
            .I(measured_delay_hc_2));
    CascadeMux I__6824 (
            .O(N__34055),
            .I(N__34052));
    InMux I__6823 (
            .O(N__34052),
            .I(N__34049));
    LocalMux I__6822 (
            .O(N__34049),
            .I(N__34043));
    InMux I__6821 (
            .O(N__34048),
            .I(N__34040));
    InMux I__6820 (
            .O(N__34047),
            .I(N__34037));
    CascadeMux I__6819 (
            .O(N__34046),
            .I(N__34034));
    Span4Mux_h I__6818 (
            .O(N__34043),
            .I(N__34031));
    LocalMux I__6817 (
            .O(N__34040),
            .I(N__34024));
    LocalMux I__6816 (
            .O(N__34037),
            .I(N__34024));
    InMux I__6815 (
            .O(N__34034),
            .I(N__34021));
    Span4Mux_v I__6814 (
            .O(N__34031),
            .I(N__34018));
    InMux I__6813 (
            .O(N__34030),
            .I(N__34015));
    InMux I__6812 (
            .O(N__34029),
            .I(N__34012));
    Span4Mux_v I__6811 (
            .O(N__34024),
            .I(N__34009));
    LocalMux I__6810 (
            .O(N__34021),
            .I(measured_delay_hc_9));
    Odrv4 I__6809 (
            .O(N__34018),
            .I(measured_delay_hc_9));
    LocalMux I__6808 (
            .O(N__34015),
            .I(measured_delay_hc_9));
    LocalMux I__6807 (
            .O(N__34012),
            .I(measured_delay_hc_9));
    Odrv4 I__6806 (
            .O(N__34009),
            .I(measured_delay_hc_9));
    InMux I__6805 (
            .O(N__33998),
            .I(N__33995));
    LocalMux I__6804 (
            .O(N__33995),
            .I(N__33992));
    Span4Mux_v I__6803 (
            .O(N__33992),
            .I(N__33989));
    Odrv4 I__6802 (
            .O(N__33989),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7 ));
    InMux I__6801 (
            .O(N__33986),
            .I(N__33983));
    LocalMux I__6800 (
            .O(N__33983),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_9 ));
    InMux I__6799 (
            .O(N__33980),
            .I(N__33977));
    LocalMux I__6798 (
            .O(N__33977),
            .I(N__33974));
    Span4Mux_v I__6797 (
            .O(N__33974),
            .I(N__33971));
    Odrv4 I__6796 (
            .O(N__33971),
            .I(\current_shift_inst.un4_control_input_axb_9 ));
    InMux I__6795 (
            .O(N__33968),
            .I(N__33965));
    LocalMux I__6794 (
            .O(N__33965),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_16 ));
    InMux I__6793 (
            .O(N__33962),
            .I(N__33959));
    LocalMux I__6792 (
            .O(N__33959),
            .I(N__33956));
    Span4Mux_h I__6791 (
            .O(N__33956),
            .I(N__33953));
    Odrv4 I__6790 (
            .O(N__33953),
            .I(\current_shift_inst.un4_control_input_axb_16 ));
    InMux I__6789 (
            .O(N__33950),
            .I(N__33947));
    LocalMux I__6788 (
            .O(N__33947),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_17 ));
    InMux I__6787 (
            .O(N__33944),
            .I(N__33941));
    LocalMux I__6786 (
            .O(N__33941),
            .I(N__33938));
    Span4Mux_h I__6785 (
            .O(N__33938),
            .I(N__33935));
    Odrv4 I__6784 (
            .O(N__33935),
            .I(\current_shift_inst.un4_control_input_axb_17 ));
    InMux I__6783 (
            .O(N__33932),
            .I(N__33929));
    LocalMux I__6782 (
            .O(N__33929),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_13 ));
    InMux I__6781 (
            .O(N__33926),
            .I(N__33923));
    LocalMux I__6780 (
            .O(N__33923),
            .I(N__33920));
    Odrv4 I__6779 (
            .O(N__33920),
            .I(\current_shift_inst.un4_control_input_axb_13 ));
    InMux I__6778 (
            .O(N__33917),
            .I(N__33913));
    InMux I__6777 (
            .O(N__33916),
            .I(N__33910));
    LocalMux I__6776 (
            .O(N__33913),
            .I(N__33907));
    LocalMux I__6775 (
            .O(N__33910),
            .I(N__33904));
    Span4Mux_v I__6774 (
            .O(N__33907),
            .I(N__33898));
    Span4Mux_h I__6773 (
            .O(N__33904),
            .I(N__33895));
    InMux I__6772 (
            .O(N__33903),
            .I(N__33892));
    InMux I__6771 (
            .O(N__33902),
            .I(N__33887));
    InMux I__6770 (
            .O(N__33901),
            .I(N__33887));
    Odrv4 I__6769 (
            .O(N__33898),
            .I(measured_delay_hc_15));
    Odrv4 I__6768 (
            .O(N__33895),
            .I(measured_delay_hc_15));
    LocalMux I__6767 (
            .O(N__33892),
            .I(measured_delay_hc_15));
    LocalMux I__6766 (
            .O(N__33887),
            .I(measured_delay_hc_15));
    InMux I__6765 (
            .O(N__33878),
            .I(N__33873));
    InMux I__6764 (
            .O(N__33877),
            .I(N__33870));
    CascadeMux I__6763 (
            .O(N__33876),
            .I(N__33867));
    LocalMux I__6762 (
            .O(N__33873),
            .I(N__33863));
    LocalMux I__6761 (
            .O(N__33870),
            .I(N__33860));
    InMux I__6760 (
            .O(N__33867),
            .I(N__33857));
    CascadeMux I__6759 (
            .O(N__33866),
            .I(N__33854));
    Span4Mux_v I__6758 (
            .O(N__33863),
            .I(N__33850));
    Span4Mux_v I__6757 (
            .O(N__33860),
            .I(N__33845));
    LocalMux I__6756 (
            .O(N__33857),
            .I(N__33845));
    InMux I__6755 (
            .O(N__33854),
            .I(N__33840));
    InMux I__6754 (
            .O(N__33853),
            .I(N__33840));
    Odrv4 I__6753 (
            .O(N__33850),
            .I(measured_delay_hc_14));
    Odrv4 I__6752 (
            .O(N__33845),
            .I(measured_delay_hc_14));
    LocalMux I__6751 (
            .O(N__33840),
            .I(measured_delay_hc_14));
    InMux I__6750 (
            .O(N__33833),
            .I(N__33827));
    InMux I__6749 (
            .O(N__33832),
            .I(N__33827));
    LocalMux I__6748 (
            .O(N__33827),
            .I(N__33823));
    InMux I__6747 (
            .O(N__33826),
            .I(N__33820));
    Span4Mux_h I__6746 (
            .O(N__33823),
            .I(N__33817));
    LocalMux I__6745 (
            .O(N__33820),
            .I(\delay_measurement_inst.tr_stateZ0Z_0 ));
    Odrv4 I__6744 (
            .O(N__33817),
            .I(\delay_measurement_inst.tr_stateZ0Z_0 ));
    InMux I__6743 (
            .O(N__33812),
            .I(N__33809));
    LocalMux I__6742 (
            .O(N__33809),
            .I(N__33806));
    Span4Mux_v I__6741 (
            .O(N__33806),
            .I(N__33801));
    InMux I__6740 (
            .O(N__33805),
            .I(N__33796));
    InMux I__6739 (
            .O(N__33804),
            .I(N__33796));
    Odrv4 I__6738 (
            .O(N__33801),
            .I(\delay_measurement_inst.prev_tr_sigZ0 ));
    LocalMux I__6737 (
            .O(N__33796),
            .I(\delay_measurement_inst.prev_tr_sigZ0 ));
    CascadeMux I__6736 (
            .O(N__33791),
            .I(\delay_measurement_inst.tr_state_RNIMR6LZ0Z_0_cascade_ ));
    InMux I__6735 (
            .O(N__33788),
            .I(N__33784));
    CascadeMux I__6734 (
            .O(N__33787),
            .I(N__33780));
    LocalMux I__6733 (
            .O(N__33784),
            .I(N__33777));
    CascadeMux I__6732 (
            .O(N__33783),
            .I(N__33774));
    InMux I__6731 (
            .O(N__33780),
            .I(N__33770));
    Span4Mux_v I__6730 (
            .O(N__33777),
            .I(N__33767));
    InMux I__6729 (
            .O(N__33774),
            .I(N__33762));
    InMux I__6728 (
            .O(N__33773),
            .I(N__33762));
    LocalMux I__6727 (
            .O(N__33770),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    Odrv4 I__6726 (
            .O(N__33767),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    LocalMux I__6725 (
            .O(N__33762),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    InMux I__6724 (
            .O(N__33755),
            .I(N__33752));
    LocalMux I__6723 (
            .O(N__33752),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_8 ));
    InMux I__6722 (
            .O(N__33749),
            .I(N__33746));
    LocalMux I__6721 (
            .O(N__33746),
            .I(N__33743));
    Odrv4 I__6720 (
            .O(N__33743),
            .I(\current_shift_inst.un4_control_input_axb_8 ));
    InMux I__6719 (
            .O(N__33740),
            .I(N__33737));
    LocalMux I__6718 (
            .O(N__33737),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_23 ));
    InMux I__6717 (
            .O(N__33734),
            .I(N__33731));
    LocalMux I__6716 (
            .O(N__33731),
            .I(N__33728));
    Span4Mux_h I__6715 (
            .O(N__33728),
            .I(N__33725));
    Odrv4 I__6714 (
            .O(N__33725),
            .I(\current_shift_inst.un4_control_input_axb_23 ));
    CascadeMux I__6713 (
            .O(N__33722),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto13_3Z0Z_1_cascade_ ));
    InMux I__6712 (
            .O(N__33719),
            .I(N__33716));
    LocalMux I__6711 (
            .O(N__33716),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto13 ));
    InMux I__6710 (
            .O(N__33713),
            .I(N__33704));
    InMux I__6709 (
            .O(N__33712),
            .I(N__33704));
    InMux I__6708 (
            .O(N__33711),
            .I(N__33704));
    LocalMux I__6707 (
            .O(N__33704),
            .I(measured_delay_hc_20));
    CascadeMux I__6706 (
            .O(N__33701),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto30_2_cascade_ ));
    InMux I__6705 (
            .O(N__33698),
            .I(N__33695));
    LocalMux I__6704 (
            .O(N__33695),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt15 ));
    InMux I__6703 (
            .O(N__33692),
            .I(N__33688));
    InMux I__6702 (
            .O(N__33691),
            .I(N__33685));
    LocalMux I__6701 (
            .O(N__33688),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1 ));
    LocalMux I__6700 (
            .O(N__33685),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1 ));
    InMux I__6699 (
            .O(N__33680),
            .I(N__33677));
    LocalMux I__6698 (
            .O(N__33677),
            .I(N__33674));
    Odrv4 I__6697 (
            .O(N__33674),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_2_tz ));
    CascadeMux I__6696 (
            .O(N__33671),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a1_1_cascade_ ));
    InMux I__6695 (
            .O(N__33668),
            .I(N__33665));
    LocalMux I__6694 (
            .O(N__33665),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_0 ));
    CascadeMux I__6693 (
            .O(N__33662),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_1_cascade_ ));
    CascadeMux I__6692 (
            .O(N__33659),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2_cascade_ ));
    InMux I__6691 (
            .O(N__33656),
            .I(N__33653));
    LocalMux I__6690 (
            .O(N__33653),
            .I(N__33650));
    Odrv4 I__6689 (
            .O(N__33650),
            .I(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2 ));
    InMux I__6688 (
            .O(N__33647),
            .I(N__33641));
    InMux I__6687 (
            .O(N__33646),
            .I(N__33641));
    LocalMux I__6686 (
            .O(N__33641),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8 ));
    CascadeMux I__6685 (
            .O(N__33638),
            .I(N__33635));
    InMux I__6684 (
            .O(N__33635),
            .I(N__33632));
    LocalMux I__6683 (
            .O(N__33632),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_1 ));
    InMux I__6682 (
            .O(N__33629),
            .I(N__33623));
    InMux I__6681 (
            .O(N__33628),
            .I(N__33623));
    LocalMux I__6680 (
            .O(N__33623),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt30 ));
    InMux I__6679 (
            .O(N__33620),
            .I(N__33617));
    LocalMux I__6678 (
            .O(N__33617),
            .I(N__33614));
    Odrv4 I__6677 (
            .O(N__33614),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9 ));
    InMux I__6676 (
            .O(N__33611),
            .I(N__33608));
    LocalMux I__6675 (
            .O(N__33608),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0 ));
    CascadeMux I__6674 (
            .O(N__33605),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0_cascade_ ));
    CascadeMux I__6673 (
            .O(N__33602),
            .I(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1_cascade_ ));
    InMux I__6672 (
            .O(N__33599),
            .I(N__33596));
    LocalMux I__6671 (
            .O(N__33596),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt30_0 ));
    InMux I__6670 (
            .O(N__33593),
            .I(N__33586));
    InMux I__6669 (
            .O(N__33592),
            .I(N__33586));
    InMux I__6668 (
            .O(N__33591),
            .I(N__33582));
    LocalMux I__6667 (
            .O(N__33586),
            .I(N__33579));
    InMux I__6666 (
            .O(N__33585),
            .I(N__33576));
    LocalMux I__6665 (
            .O(N__33582),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    Odrv12 I__6664 (
            .O(N__33579),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    LocalMux I__6663 (
            .O(N__33576),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    InMux I__6662 (
            .O(N__33569),
            .I(N__33566));
    LocalMux I__6661 (
            .O(N__33566),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8 ));
    CascadeMux I__6660 (
            .O(N__33563),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_2_cascade_ ));
    InMux I__6659 (
            .O(N__33560),
            .I(N__33557));
    LocalMux I__6658 (
            .O(N__33557),
            .I(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_11 ));
    InMux I__6657 (
            .O(N__33554),
            .I(N__33550));
    InMux I__6656 (
            .O(N__33553),
            .I(N__33547));
    LocalMux I__6655 (
            .O(N__33550),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_1 ));
    LocalMux I__6654 (
            .O(N__33547),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_1 ));
    InMux I__6653 (
            .O(N__33542),
            .I(N__33538));
    InMux I__6652 (
            .O(N__33541),
            .I(N__33535));
    LocalMux I__6651 (
            .O(N__33538),
            .I(N__33530));
    LocalMux I__6650 (
            .O(N__33535),
            .I(N__33530));
    Sp12to4 I__6649 (
            .O(N__33530),
            .I(N__33526));
    InMux I__6648 (
            .O(N__33529),
            .I(N__33523));
    Span12Mux_v I__6647 (
            .O(N__33526),
            .I(N__33520));
    LocalMux I__6646 (
            .O(N__33523),
            .I(\current_shift_inst.start_timer_phaseZ0 ));
    Odrv12 I__6645 (
            .O(N__33520),
            .I(\current_shift_inst.start_timer_phaseZ0 ));
    InMux I__6644 (
            .O(N__33515),
            .I(N__33509));
    InMux I__6643 (
            .O(N__33514),
            .I(N__33506));
    InMux I__6642 (
            .O(N__33513),
            .I(N__33503));
    InMux I__6641 (
            .O(N__33512),
            .I(N__33500));
    LocalMux I__6640 (
            .O(N__33509),
            .I(\current_shift_inst.timer_phase.runningZ0 ));
    LocalMux I__6639 (
            .O(N__33506),
            .I(\current_shift_inst.timer_phase.runningZ0 ));
    LocalMux I__6638 (
            .O(N__33503),
            .I(\current_shift_inst.timer_phase.runningZ0 ));
    LocalMux I__6637 (
            .O(N__33500),
            .I(\current_shift_inst.timer_phase.runningZ0 ));
    InMux I__6636 (
            .O(N__33491),
            .I(N__33486));
    InMux I__6635 (
            .O(N__33490),
            .I(N__33483));
    InMux I__6634 (
            .O(N__33489),
            .I(N__33479));
    LocalMux I__6633 (
            .O(N__33486),
            .I(N__33476));
    LocalMux I__6632 (
            .O(N__33483),
            .I(N__33473));
    CascadeMux I__6631 (
            .O(N__33482),
            .I(N__33470));
    LocalMux I__6630 (
            .O(N__33479),
            .I(N__33463));
    Sp12to4 I__6629 (
            .O(N__33476),
            .I(N__33463));
    Span12Mux_s4_v I__6628 (
            .O(N__33473),
            .I(N__33463));
    InMux I__6627 (
            .O(N__33470),
            .I(N__33460));
    Span12Mux_v I__6626 (
            .O(N__33463),
            .I(N__33457));
    LocalMux I__6625 (
            .O(N__33460),
            .I(\current_shift_inst.stop_timer_phaseZ0 ));
    Odrv12 I__6624 (
            .O(N__33457),
            .I(\current_shift_inst.stop_timer_phaseZ0 ));
    IoInMux I__6623 (
            .O(N__33452),
            .I(N__33449));
    LocalMux I__6622 (
            .O(N__33449),
            .I(N__33446));
    Odrv12 I__6621 (
            .O(N__33446),
            .I(\current_shift_inst.timer_phase.N_188_i ));
    IoInMux I__6620 (
            .O(N__33443),
            .I(N__33440));
    LocalMux I__6619 (
            .O(N__33440),
            .I(N__33437));
    Odrv4 I__6618 (
            .O(N__33437),
            .I(s2_phy_c));
    CascadeMux I__6617 (
            .O(N__33434),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_3_cascade_ ));
    InMux I__6616 (
            .O(N__33431),
            .I(N__33428));
    LocalMux I__6615 (
            .O(N__33428),
            .I(N__33423));
    InMux I__6614 (
            .O(N__33427),
            .I(N__33420));
    InMux I__6613 (
            .O(N__33426),
            .I(N__33417));
    Span4Mux_v I__6612 (
            .O(N__33423),
            .I(N__33412));
    LocalMux I__6611 (
            .O(N__33420),
            .I(N__33412));
    LocalMux I__6610 (
            .O(N__33417),
            .I(N__33409));
    Odrv4 I__6609 (
            .O(N__33412),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    Odrv12 I__6608 (
            .O(N__33409),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    CascadeMux I__6607 (
            .O(N__33404),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt14_cascade_ ));
    InMux I__6606 (
            .O(N__33401),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9 ));
    InMux I__6605 (
            .O(N__33398),
            .I(N__33395));
    LocalMux I__6604 (
            .O(N__33395),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12 ));
    InMux I__6603 (
            .O(N__33392),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10 ));
    InMux I__6602 (
            .O(N__33389),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11 ));
    InMux I__6601 (
            .O(N__33386),
            .I(N__33383));
    LocalMux I__6600 (
            .O(N__33383),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14 ));
    InMux I__6599 (
            .O(N__33380),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12 ));
    InMux I__6598 (
            .O(N__33377),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13 ));
    InMux I__6597 (
            .O(N__33374),
            .I(N__33371));
    LocalMux I__6596 (
            .O(N__33371),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16 ));
    InMux I__6595 (
            .O(N__33368),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14 ));
    InMux I__6594 (
            .O(N__33365),
            .I(bfn_13_25_0_));
    InMux I__6593 (
            .O(N__33362),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16 ));
    InMux I__6592 (
            .O(N__33359),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17 ));
    InMux I__6591 (
            .O(N__33356),
            .I(N__33353));
    LocalMux I__6590 (
            .O(N__33353),
            .I(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19 ));
    InMux I__6589 (
            .O(N__33350),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0 ));
    InMux I__6588 (
            .O(N__33347),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1 ));
    InMux I__6587 (
            .O(N__33344),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2 ));
    InMux I__6586 (
            .O(N__33341),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3 ));
    InMux I__6585 (
            .O(N__33338),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4 ));
    InMux I__6584 (
            .O(N__33335),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5 ));
    InMux I__6583 (
            .O(N__33332),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6 ));
    InMux I__6582 (
            .O(N__33329),
            .I(bfn_13_24_0_));
    InMux I__6581 (
            .O(N__33326),
            .I(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8 ));
    CascadeMux I__6580 (
            .O(N__33323),
            .I(N__33320));
    InMux I__6579 (
            .O(N__33320),
            .I(N__33317));
    LocalMux I__6578 (
            .O(N__33317),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_18 ));
    CascadeMux I__6577 (
            .O(N__33314),
            .I(N__33311));
    InMux I__6576 (
            .O(N__33311),
            .I(N__33308));
    LocalMux I__6575 (
            .O(N__33308),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_19 ));
    InMux I__6574 (
            .O(N__33305),
            .I(N__33298));
    InMux I__6573 (
            .O(N__33304),
            .I(N__33298));
    InMux I__6572 (
            .O(N__33303),
            .I(N__33295));
    LocalMux I__6571 (
            .O(N__33298),
            .I(\phase_controller_slave.stateZ0Z_0 ));
    LocalMux I__6570 (
            .O(N__33295),
            .I(\phase_controller_slave.stateZ0Z_0 ));
    CascadeMux I__6569 (
            .O(N__33290),
            .I(N__33284));
    InMux I__6568 (
            .O(N__33289),
            .I(N__33281));
    InMux I__6567 (
            .O(N__33288),
            .I(N__33278));
    InMux I__6566 (
            .O(N__33287),
            .I(N__33273));
    InMux I__6565 (
            .O(N__33284),
            .I(N__33273));
    LocalMux I__6564 (
            .O(N__33281),
            .I(\phase_controller_slave.stateZ0Z_4 ));
    LocalMux I__6563 (
            .O(N__33278),
            .I(\phase_controller_slave.stateZ0Z_4 ));
    LocalMux I__6562 (
            .O(N__33273),
            .I(\phase_controller_slave.stateZ0Z_4 ));
    InMux I__6561 (
            .O(N__33266),
            .I(N__33263));
    LocalMux I__6560 (
            .O(N__33263),
            .I(N__33260));
    Span4Mux_v I__6559 (
            .O(N__33260),
            .I(N__33257));
    Odrv4 I__6558 (
            .O(N__33257),
            .I(\phase_controller_slave.start_timer_tr_0_sqmuxa ));
    CascadeMux I__6557 (
            .O(N__33254),
            .I(\phase_controller_slave.N_210_cascade_ ));
    CascadeMux I__6556 (
            .O(N__33251),
            .I(\phase_controller_slave.stoper_tr.time_passed11_cascade_ ));
    CascadeMux I__6555 (
            .O(N__33248),
            .I(N__33244));
    InMux I__6554 (
            .O(N__33247),
            .I(N__33239));
    InMux I__6553 (
            .O(N__33244),
            .I(N__33236));
    InMux I__6552 (
            .O(N__33243),
            .I(N__33231));
    InMux I__6551 (
            .O(N__33242),
            .I(N__33231));
    LocalMux I__6550 (
            .O(N__33239),
            .I(\phase_controller_slave.tr_time_passed ));
    LocalMux I__6549 (
            .O(N__33236),
            .I(\phase_controller_slave.tr_time_passed ));
    LocalMux I__6548 (
            .O(N__33231),
            .I(\phase_controller_slave.tr_time_passed ));
    InMux I__6547 (
            .O(N__33224),
            .I(N__33221));
    LocalMux I__6546 (
            .O(N__33221),
            .I(\phase_controller_slave.stoper_tr.time_passed_1_sqmuxa ));
    CascadeMux I__6545 (
            .O(N__33218),
            .I(N__33215));
    InMux I__6544 (
            .O(N__33215),
            .I(N__33212));
    LocalMux I__6543 (
            .O(N__33212),
            .I(N__33209));
    Span4Mux_h I__6542 (
            .O(N__33209),
            .I(N__33206));
    Odrv4 I__6541 (
            .O(N__33206),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_14 ));
    InMux I__6540 (
            .O(N__33203),
            .I(N__33200));
    LocalMux I__6539 (
            .O(N__33200),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_14 ));
    CascadeMux I__6538 (
            .O(N__33197),
            .I(N__33194));
    InMux I__6537 (
            .O(N__33194),
            .I(N__33191));
    LocalMux I__6536 (
            .O(N__33191),
            .I(N__33188));
    Span4Mux_v I__6535 (
            .O(N__33188),
            .I(N__33185));
    Span4Mux_v I__6534 (
            .O(N__33185),
            .I(N__33182));
    Odrv4 I__6533 (
            .O(N__33182),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_15 ));
    InMux I__6532 (
            .O(N__33179),
            .I(N__33176));
    LocalMux I__6531 (
            .O(N__33176),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_15 ));
    InMux I__6530 (
            .O(N__33173),
            .I(N__33170));
    LocalMux I__6529 (
            .O(N__33170),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_16 ));
    InMux I__6528 (
            .O(N__33167),
            .I(N__33164));
    LocalMux I__6527 (
            .O(N__33164),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_17 ));
    InMux I__6526 (
            .O(N__33161),
            .I(N__33158));
    LocalMux I__6525 (
            .O(N__33158),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_18 ));
    InMux I__6524 (
            .O(N__33155),
            .I(N__33152));
    LocalMux I__6523 (
            .O(N__33152),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_19 ));
    InMux I__6522 (
            .O(N__33149),
            .I(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19 ));
    CascadeMux I__6521 (
            .O(N__33146),
            .I(N__33143));
    InMux I__6520 (
            .O(N__33143),
            .I(N__33140));
    LocalMux I__6519 (
            .O(N__33140),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_17 ));
    CascadeMux I__6518 (
            .O(N__33137),
            .I(N__33134));
    InMux I__6517 (
            .O(N__33134),
            .I(N__33131));
    LocalMux I__6516 (
            .O(N__33131),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_6 ));
    InMux I__6515 (
            .O(N__33128),
            .I(N__33125));
    LocalMux I__6514 (
            .O(N__33125),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_6 ));
    CascadeMux I__6513 (
            .O(N__33122),
            .I(N__33119));
    InMux I__6512 (
            .O(N__33119),
            .I(N__33116));
    LocalMux I__6511 (
            .O(N__33116),
            .I(N__33113));
    Odrv4 I__6510 (
            .O(N__33113),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_7 ));
    InMux I__6509 (
            .O(N__33110),
            .I(N__33107));
    LocalMux I__6508 (
            .O(N__33107),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_7 ));
    CascadeMux I__6507 (
            .O(N__33104),
            .I(N__33101));
    InMux I__6506 (
            .O(N__33101),
            .I(N__33098));
    LocalMux I__6505 (
            .O(N__33098),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_8 ));
    InMux I__6504 (
            .O(N__33095),
            .I(N__33092));
    LocalMux I__6503 (
            .O(N__33092),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_8 ));
    CascadeMux I__6502 (
            .O(N__33089),
            .I(N__33086));
    InMux I__6501 (
            .O(N__33086),
            .I(N__33083));
    LocalMux I__6500 (
            .O(N__33083),
            .I(N__33080));
    Odrv4 I__6499 (
            .O(N__33080),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_9 ));
    InMux I__6498 (
            .O(N__33077),
            .I(N__33074));
    LocalMux I__6497 (
            .O(N__33074),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_9 ));
    CascadeMux I__6496 (
            .O(N__33071),
            .I(N__33068));
    InMux I__6495 (
            .O(N__33068),
            .I(N__33065));
    LocalMux I__6494 (
            .O(N__33065),
            .I(N__33062));
    Span12Mux_h I__6493 (
            .O(N__33062),
            .I(N__33059));
    Odrv12 I__6492 (
            .O(N__33059),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_10 ));
    InMux I__6491 (
            .O(N__33056),
            .I(N__33053));
    LocalMux I__6490 (
            .O(N__33053),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_10 ));
    CascadeMux I__6489 (
            .O(N__33050),
            .I(N__33047));
    InMux I__6488 (
            .O(N__33047),
            .I(N__33044));
    LocalMux I__6487 (
            .O(N__33044),
            .I(N__33041));
    Span4Mux_v I__6486 (
            .O(N__33041),
            .I(N__33038));
    Span4Mux_v I__6485 (
            .O(N__33038),
            .I(N__33035));
    Odrv4 I__6484 (
            .O(N__33035),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_11 ));
    InMux I__6483 (
            .O(N__33032),
            .I(N__33029));
    LocalMux I__6482 (
            .O(N__33029),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_11 ));
    CascadeMux I__6481 (
            .O(N__33026),
            .I(N__33023));
    InMux I__6480 (
            .O(N__33023),
            .I(N__33020));
    LocalMux I__6479 (
            .O(N__33020),
            .I(N__33017));
    Span4Mux_v I__6478 (
            .O(N__33017),
            .I(N__33014));
    Span4Mux_v I__6477 (
            .O(N__33014),
            .I(N__33011));
    Odrv4 I__6476 (
            .O(N__33011),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_12 ));
    InMux I__6475 (
            .O(N__33008),
            .I(N__33005));
    LocalMux I__6474 (
            .O(N__33005),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_12 ));
    CascadeMux I__6473 (
            .O(N__33002),
            .I(N__32999));
    InMux I__6472 (
            .O(N__32999),
            .I(N__32996));
    LocalMux I__6471 (
            .O(N__32996),
            .I(N__32993));
    Span4Mux_v I__6470 (
            .O(N__32993),
            .I(N__32990));
    Span4Mux_v I__6469 (
            .O(N__32990),
            .I(N__32987));
    Odrv4 I__6468 (
            .O(N__32987),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_13 ));
    InMux I__6467 (
            .O(N__32984),
            .I(N__32981));
    LocalMux I__6466 (
            .O(N__32981),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_13 ));
    CascadeMux I__6465 (
            .O(N__32978),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6_cascade_ ));
    CascadeMux I__6464 (
            .O(N__32975),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13_cascade_ ));
    CascadeMux I__6463 (
            .O(N__32972),
            .I(N__32969));
    InMux I__6462 (
            .O(N__32969),
            .I(N__32966));
    LocalMux I__6461 (
            .O(N__32966),
            .I(N__32963));
    Odrv4 I__6460 (
            .O(N__32963),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_1 ));
    InMux I__6459 (
            .O(N__32960),
            .I(N__32957));
    LocalMux I__6458 (
            .O(N__32957),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_1 ));
    CascadeMux I__6457 (
            .O(N__32954),
            .I(N__32951));
    InMux I__6456 (
            .O(N__32951),
            .I(N__32948));
    LocalMux I__6455 (
            .O(N__32948),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_2 ));
    InMux I__6454 (
            .O(N__32945),
            .I(N__32942));
    LocalMux I__6453 (
            .O(N__32942),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_2 ));
    CascadeMux I__6452 (
            .O(N__32939),
            .I(N__32936));
    InMux I__6451 (
            .O(N__32936),
            .I(N__32933));
    LocalMux I__6450 (
            .O(N__32933),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_3 ));
    InMux I__6449 (
            .O(N__32930),
            .I(N__32927));
    LocalMux I__6448 (
            .O(N__32927),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_3 ));
    CascadeMux I__6447 (
            .O(N__32924),
            .I(N__32921));
    InMux I__6446 (
            .O(N__32921),
            .I(N__32918));
    LocalMux I__6445 (
            .O(N__32918),
            .I(N__32915));
    Odrv4 I__6444 (
            .O(N__32915),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_4 ));
    InMux I__6443 (
            .O(N__32912),
            .I(N__32909));
    LocalMux I__6442 (
            .O(N__32909),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_4 ));
    CascadeMux I__6441 (
            .O(N__32906),
            .I(N__32903));
    InMux I__6440 (
            .O(N__32903),
            .I(N__32900));
    LocalMux I__6439 (
            .O(N__32900),
            .I(N__32897));
    Odrv12 I__6438 (
            .O(N__32897),
            .I(\phase_controller_slave.stoper_tr.target_timeZ0Z_5 ));
    InMux I__6437 (
            .O(N__32894),
            .I(N__32891));
    LocalMux I__6436 (
            .O(N__32891),
            .I(\phase_controller_slave.stoper_tr.accumulated_time_i_5 ));
    IoInMux I__6435 (
            .O(N__32888),
            .I(N__32885));
    LocalMux I__6434 (
            .O(N__32885),
            .I(N__32882));
    IoSpan4Mux I__6433 (
            .O(N__32882),
            .I(N__32879));
    Span4Mux_s3_v I__6432 (
            .O(N__32879),
            .I(N__32876));
    Span4Mux_v I__6431 (
            .O(N__32876),
            .I(N__32872));
    InMux I__6430 (
            .O(N__32875),
            .I(N__32869));
    Span4Mux_v I__6429 (
            .O(N__32872),
            .I(N__32866));
    LocalMux I__6428 (
            .O(N__32869),
            .I(N__32863));
    Span4Mux_v I__6427 (
            .O(N__32866),
            .I(N__32858));
    Span4Mux_v I__6426 (
            .O(N__32863),
            .I(N__32858));
    Odrv4 I__6425 (
            .O(N__32858),
            .I(s1_phy_c));
    InMux I__6424 (
            .O(N__32855),
            .I(N__32852));
    LocalMux I__6423 (
            .O(N__32852),
            .I(\current_shift_inst.S1_syncZ0Z0 ));
    InMux I__6422 (
            .O(N__32849),
            .I(N__32846));
    LocalMux I__6421 (
            .O(N__32846),
            .I(\current_shift_inst.S3_sync_prevZ0 ));
    InMux I__6420 (
            .O(N__32843),
            .I(N__32839));
    CascadeMux I__6419 (
            .O(N__32842),
            .I(N__32835));
    LocalMux I__6418 (
            .O(N__32839),
            .I(N__32832));
    InMux I__6417 (
            .O(N__32838),
            .I(N__32827));
    InMux I__6416 (
            .O(N__32835),
            .I(N__32827));
    Span4Mux_h I__6415 (
            .O(N__32832),
            .I(N__32822));
    LocalMux I__6414 (
            .O(N__32827),
            .I(N__32822));
    Sp12to4 I__6413 (
            .O(N__32822),
            .I(N__32819));
    Odrv12 I__6412 (
            .O(N__32819),
            .I(\current_shift_inst.S3_riseZ0 ));
    InMux I__6411 (
            .O(N__32816),
            .I(N__32810));
    InMux I__6410 (
            .O(N__32815),
            .I(N__32810));
    LocalMux I__6409 (
            .O(N__32810),
            .I(\current_shift_inst.S1_syncZ0Z1 ));
    InMux I__6408 (
            .O(N__32807),
            .I(N__32804));
    LocalMux I__6407 (
            .O(N__32804),
            .I(\current_shift_inst.S1_sync_prevZ0 ));
    InMux I__6406 (
            .O(N__32801),
            .I(N__32798));
    LocalMux I__6405 (
            .O(N__32798),
            .I(\current_shift_inst.S3_syncZ0Z0 ));
    InMux I__6404 (
            .O(N__32795),
            .I(N__32789));
    InMux I__6403 (
            .O(N__32794),
            .I(N__32789));
    LocalMux I__6402 (
            .O(N__32789),
            .I(\current_shift_inst.S3_syncZ0Z1 ));
    InMux I__6401 (
            .O(N__32786),
            .I(N__32783));
    LocalMux I__6400 (
            .O(N__32783),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_26 ));
    InMux I__6399 (
            .O(N__32780),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ));
    InMux I__6398 (
            .O(N__32777),
            .I(N__32774));
    LocalMux I__6397 (
            .O(N__32774),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_27 ));
    InMux I__6396 (
            .O(N__32771),
            .I(bfn_13_16_0_));
    InMux I__6395 (
            .O(N__32768),
            .I(N__32765));
    LocalMux I__6394 (
            .O(N__32765),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_28 ));
    InMux I__6393 (
            .O(N__32762),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ));
    InMux I__6392 (
            .O(N__32759),
            .I(N__32756));
    LocalMux I__6391 (
            .O(N__32756),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_29 ));
    InMux I__6390 (
            .O(N__32753),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ));
    InMux I__6389 (
            .O(N__32750),
            .I(N__32747));
    LocalMux I__6388 (
            .O(N__32747),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_30 ));
    InMux I__6387 (
            .O(N__32744),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ));
    CEMux I__6386 (
            .O(N__32741),
            .I(N__32726));
    CEMux I__6385 (
            .O(N__32740),
            .I(N__32726));
    CEMux I__6384 (
            .O(N__32739),
            .I(N__32726));
    CEMux I__6383 (
            .O(N__32738),
            .I(N__32726));
    CEMux I__6382 (
            .O(N__32737),
            .I(N__32726));
    GlobalMux I__6381 (
            .O(N__32726),
            .I(N__32723));
    gio2CtrlBuf I__6380 (
            .O(N__32723),
            .I(\current_shift_inst.timer_s1.N_187_i_g ));
    InMux I__6379 (
            .O(N__32720),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ));
    InMux I__6378 (
            .O(N__32717),
            .I(N__32711));
    InMux I__6377 (
            .O(N__32716),
            .I(N__32711));
    LocalMux I__6376 (
            .O(N__32711),
            .I(N__32708));
    Span4Mux_v I__6375 (
            .O(N__32708),
            .I(N__32705));
    Odrv4 I__6374 (
            .O(N__32705),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    InMux I__6373 (
            .O(N__32702),
            .I(N__32691));
    InMux I__6372 (
            .O(N__32701),
            .I(N__32691));
    InMux I__6371 (
            .O(N__32700),
            .I(N__32680));
    InMux I__6370 (
            .O(N__32699),
            .I(N__32680));
    InMux I__6369 (
            .O(N__32698),
            .I(N__32680));
    InMux I__6368 (
            .O(N__32697),
            .I(N__32680));
    InMux I__6367 (
            .O(N__32696),
            .I(N__32680));
    LocalMux I__6366 (
            .O(N__32691),
            .I(N__32675));
    LocalMux I__6365 (
            .O(N__32680),
            .I(N__32675));
    Odrv12 I__6364 (
            .O(N__32675),
            .I(\current_shift_inst.S1_riseZ0 ));
    InMux I__6363 (
            .O(N__32672),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ));
    InMux I__6362 (
            .O(N__32669),
            .I(N__32666));
    LocalMux I__6361 (
            .O(N__32666),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_18 ));
    InMux I__6360 (
            .O(N__32663),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ));
    InMux I__6359 (
            .O(N__32660),
            .I(N__32657));
    LocalMux I__6358 (
            .O(N__32657),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_19 ));
    InMux I__6357 (
            .O(N__32654),
            .I(bfn_13_15_0_));
    InMux I__6356 (
            .O(N__32651),
            .I(N__32648));
    LocalMux I__6355 (
            .O(N__32648),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_20 ));
    InMux I__6354 (
            .O(N__32645),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ));
    InMux I__6353 (
            .O(N__32642),
            .I(N__32639));
    LocalMux I__6352 (
            .O(N__32639),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_21 ));
    InMux I__6351 (
            .O(N__32636),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ));
    InMux I__6350 (
            .O(N__32633),
            .I(N__32630));
    LocalMux I__6349 (
            .O(N__32630),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_22 ));
    InMux I__6348 (
            .O(N__32627),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ));
    InMux I__6347 (
            .O(N__32624),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ));
    InMux I__6346 (
            .O(N__32621),
            .I(N__32618));
    LocalMux I__6345 (
            .O(N__32618),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_24 ));
    InMux I__6344 (
            .O(N__32615),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ));
    InMux I__6343 (
            .O(N__32612),
            .I(N__32609));
    LocalMux I__6342 (
            .O(N__32609),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_25 ));
    InMux I__6341 (
            .O(N__32606),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ));
    InMux I__6340 (
            .O(N__32603),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ));
    InMux I__6339 (
            .O(N__32600),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ));
    InMux I__6338 (
            .O(N__32597),
            .I(N__32594));
    LocalMux I__6337 (
            .O(N__32594),
            .I(N__32591));
    Odrv4 I__6336 (
            .O(N__32591),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_10 ));
    InMux I__6335 (
            .O(N__32588),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ));
    InMux I__6334 (
            .O(N__32585),
            .I(N__32582));
    LocalMux I__6333 (
            .O(N__32582),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_11 ));
    InMux I__6332 (
            .O(N__32579),
            .I(bfn_13_14_0_));
    InMux I__6331 (
            .O(N__32576),
            .I(N__32573));
    LocalMux I__6330 (
            .O(N__32573),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_12 ));
    InMux I__6329 (
            .O(N__32570),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ));
    InMux I__6328 (
            .O(N__32567),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ));
    InMux I__6327 (
            .O(N__32564),
            .I(N__32561));
    LocalMux I__6326 (
            .O(N__32561),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_14 ));
    InMux I__6325 (
            .O(N__32558),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ));
    InMux I__6324 (
            .O(N__32555),
            .I(N__32552));
    LocalMux I__6323 (
            .O(N__32552),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_15 ));
    InMux I__6322 (
            .O(N__32549),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ));
    InMux I__6321 (
            .O(N__32546),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ));
    InMux I__6320 (
            .O(N__32543),
            .I(N__32540));
    LocalMux I__6319 (
            .O(N__32540),
            .I(N__32535));
    InMux I__6318 (
            .O(N__32539),
            .I(N__32532));
    InMux I__6317 (
            .O(N__32538),
            .I(N__32529));
    Span4Mux_v I__6316 (
            .O(N__32535),
            .I(N__32526));
    LocalMux I__6315 (
            .O(N__32532),
            .I(N__32521));
    LocalMux I__6314 (
            .O(N__32529),
            .I(N__32521));
    Span4Mux_h I__6313 (
            .O(N__32526),
            .I(N__32518));
    Span4Mux_v I__6312 (
            .O(N__32521),
            .I(N__32515));
    Odrv4 I__6311 (
            .O(N__32518),
            .I(il_max_comp1_D2));
    Odrv4 I__6310 (
            .O(N__32515),
            .I(il_max_comp1_D2));
    CascadeMux I__6309 (
            .O(N__32510),
            .I(\phase_controller_inst1.N_86_cascade_ ));
    InMux I__6308 (
            .O(N__32507),
            .I(N__32499));
    InMux I__6307 (
            .O(N__32506),
            .I(N__32499));
    InMux I__6306 (
            .O(N__32505),
            .I(N__32496));
    InMux I__6305 (
            .O(N__32504),
            .I(N__32493));
    LocalMux I__6304 (
            .O(N__32499),
            .I(\phase_controller_inst1.stateZ0Z_3 ));
    LocalMux I__6303 (
            .O(N__32496),
            .I(\phase_controller_inst1.stateZ0Z_3 ));
    LocalMux I__6302 (
            .O(N__32493),
            .I(\phase_controller_inst1.stateZ0Z_3 ));
    InMux I__6301 (
            .O(N__32486),
            .I(N__32483));
    LocalMux I__6300 (
            .O(N__32483),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_3 ));
    InMux I__6299 (
            .O(N__32480),
            .I(N__32477));
    LocalMux I__6298 (
            .O(N__32477),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_4 ));
    InMux I__6297 (
            .O(N__32474),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ));
    InMux I__6296 (
            .O(N__32471),
            .I(N__32468));
    LocalMux I__6295 (
            .O(N__32468),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_5 ));
    InMux I__6294 (
            .O(N__32465),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ));
    InMux I__6293 (
            .O(N__32462),
            .I(N__32459));
    LocalMux I__6292 (
            .O(N__32459),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_6 ));
    InMux I__6291 (
            .O(N__32456),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ));
    InMux I__6290 (
            .O(N__32453),
            .I(N__32450));
    LocalMux I__6289 (
            .O(N__32450),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_7 ));
    InMux I__6288 (
            .O(N__32447),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ));
    InMux I__6287 (
            .O(N__32444),
            .I(N__32441));
    LocalMux I__6286 (
            .O(N__32441),
            .I(\phase_controller_inst1.stoper_hc.un1_startlt8 ));
    CascadeMux I__6285 (
            .O(N__32438),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8_cascade_ ));
    InMux I__6284 (
            .O(N__32435),
            .I(N__32432));
    LocalMux I__6283 (
            .O(N__32432),
            .I(N__32429));
    Odrv4 I__6282 (
            .O(N__32429),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_10 ));
    InMux I__6281 (
            .O(N__32426),
            .I(N__32423));
    LocalMux I__6280 (
            .O(N__32423),
            .I(N__32420));
    Span4Mux_v I__6279 (
            .O(N__32420),
            .I(N__32417));
    Odrv4 I__6278 (
            .O(N__32417),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_13 ));
    IoInMux I__6277 (
            .O(N__32414),
            .I(N__32411));
    LocalMux I__6276 (
            .O(N__32411),
            .I(N__32408));
    Span4Mux_s0_v I__6275 (
            .O(N__32408),
            .I(N__32405));
    Sp12to4 I__6274 (
            .O(N__32405),
            .I(N__32402));
    Span12Mux_h I__6273 (
            .O(N__32402),
            .I(N__32399));
    Span12Mux_v I__6272 (
            .O(N__32399),
            .I(N__32396));
    Odrv12 I__6271 (
            .O(N__32396),
            .I(\current_shift_inst.timer_s1.N_187_i ));
    InMux I__6270 (
            .O(N__32393),
            .I(N__32389));
    CascadeMux I__6269 (
            .O(N__32392),
            .I(N__32386));
    LocalMux I__6268 (
            .O(N__32389),
            .I(N__32382));
    InMux I__6267 (
            .O(N__32386),
            .I(N__32375));
    InMux I__6266 (
            .O(N__32385),
            .I(N__32375));
    Span4Mux_h I__6265 (
            .O(N__32382),
            .I(N__32372));
    InMux I__6264 (
            .O(N__32381),
            .I(N__32367));
    InMux I__6263 (
            .O(N__32380),
            .I(N__32367));
    LocalMux I__6262 (
            .O(N__32375),
            .I(N__32362));
    Span4Mux_h I__6261 (
            .O(N__32372),
            .I(N__32362));
    LocalMux I__6260 (
            .O(N__32367),
            .I(\current_shift_inst.phase_validZ0 ));
    Odrv4 I__6259 (
            .O(N__32362),
            .I(\current_shift_inst.phase_validZ0 ));
    CascadeMux I__6258 (
            .O(N__32357),
            .I(N__32353));
    CascadeMux I__6257 (
            .O(N__32356),
            .I(N__32347));
    InMux I__6256 (
            .O(N__32353),
            .I(N__32342));
    InMux I__6255 (
            .O(N__32352),
            .I(N__32342));
    InMux I__6254 (
            .O(N__32351),
            .I(N__32335));
    InMux I__6253 (
            .O(N__32350),
            .I(N__32335));
    InMux I__6252 (
            .O(N__32347),
            .I(N__32335));
    LocalMux I__6251 (
            .O(N__32342),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    LocalMux I__6250 (
            .O(N__32335),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    InMux I__6249 (
            .O(N__32330),
            .I(N__32324));
    InMux I__6248 (
            .O(N__32329),
            .I(N__32321));
    InMux I__6247 (
            .O(N__32328),
            .I(N__32316));
    InMux I__6246 (
            .O(N__32327),
            .I(N__32316));
    LocalMux I__6245 (
            .O(N__32324),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__6244 (
            .O(N__32321),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__6243 (
            .O(N__32316),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    CascadeMux I__6242 (
            .O(N__32309),
            .I(N__32301));
    InMux I__6241 (
            .O(N__32308),
            .I(N__32293));
    InMux I__6240 (
            .O(N__32307),
            .I(N__32293));
    InMux I__6239 (
            .O(N__32306),
            .I(N__32293));
    InMux I__6238 (
            .O(N__32305),
            .I(N__32288));
    InMux I__6237 (
            .O(N__32304),
            .I(N__32288));
    InMux I__6236 (
            .O(N__32301),
            .I(N__32283));
    InMux I__6235 (
            .O(N__32300),
            .I(N__32283));
    LocalMux I__6234 (
            .O(N__32293),
            .I(\current_shift_inst.meas_stateZ0Z_0 ));
    LocalMux I__6233 (
            .O(N__32288),
            .I(\current_shift_inst.meas_stateZ0Z_0 ));
    LocalMux I__6232 (
            .O(N__32283),
            .I(\current_shift_inst.meas_stateZ0Z_0 ));
    CascadeMux I__6231 (
            .O(N__32276),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto5Z0Z_3_cascade_ ));
    IoInMux I__6230 (
            .O(N__32273),
            .I(N__32270));
    LocalMux I__6229 (
            .O(N__32270),
            .I(N__32267));
    Span4Mux_s0_v I__6228 (
            .O(N__32267),
            .I(N__32264));
    Span4Mux_v I__6227 (
            .O(N__32264),
            .I(N__32261));
    Odrv4 I__6226 (
            .O(N__32261),
            .I(\delay_measurement_inst.delay_hc_timer.N_321_i ));
    CascadeMux I__6225 (
            .O(N__32258),
            .I(\current_shift_inst.N_199_cascade_ ));
    InMux I__6224 (
            .O(N__32255),
            .I(N__32252));
    LocalMux I__6223 (
            .O(N__32252),
            .I(N__32247));
    CascadeMux I__6222 (
            .O(N__32251),
            .I(N__32243));
    InMux I__6221 (
            .O(N__32250),
            .I(N__32240));
    Span4Mux_v I__6220 (
            .O(N__32247),
            .I(N__32237));
    InMux I__6219 (
            .O(N__32246),
            .I(N__32234));
    InMux I__6218 (
            .O(N__32243),
            .I(N__32231));
    LocalMux I__6217 (
            .O(N__32240),
            .I(N__32228));
    Odrv4 I__6216 (
            .O(N__32237),
            .I(\phase_controller_slave.stateZ0Z_1 ));
    LocalMux I__6215 (
            .O(N__32234),
            .I(\phase_controller_slave.stateZ0Z_1 ));
    LocalMux I__6214 (
            .O(N__32231),
            .I(\phase_controller_slave.stateZ0Z_1 ));
    Odrv4 I__6213 (
            .O(N__32228),
            .I(\phase_controller_slave.stateZ0Z_1 ));
    InMux I__6212 (
            .O(N__32219),
            .I(N__32214));
    InMux I__6211 (
            .O(N__32218),
            .I(N__32211));
    InMux I__6210 (
            .O(N__32217),
            .I(N__32208));
    LocalMux I__6209 (
            .O(N__32214),
            .I(N__32203));
    LocalMux I__6208 (
            .O(N__32211),
            .I(N__32203));
    LocalMux I__6207 (
            .O(N__32208),
            .I(N__32200));
    Span4Mux_h I__6206 (
            .O(N__32203),
            .I(N__32197));
    Span4Mux_h I__6205 (
            .O(N__32200),
            .I(N__32194));
    Span4Mux_v I__6204 (
            .O(N__32197),
            .I(N__32191));
    Span4Mux_v I__6203 (
            .O(N__32194),
            .I(N__32188));
    Sp12to4 I__6202 (
            .O(N__32191),
            .I(N__32185));
    Span4Mux_v I__6201 (
            .O(N__32188),
            .I(N__32182));
    Span12Mux_v I__6200 (
            .O(N__32185),
            .I(N__32179));
    Span4Mux_v I__6199 (
            .O(N__32182),
            .I(N__32176));
    Odrv12 I__6198 (
            .O(N__32179),
            .I(il_min_comp2_D2));
    Odrv4 I__6197 (
            .O(N__32176),
            .I(il_min_comp2_D2));
    CascadeMux I__6196 (
            .O(N__32171),
            .I(N__32168));
    InMux I__6195 (
            .O(N__32168),
            .I(N__32163));
    InMux I__6194 (
            .O(N__32167),
            .I(N__32158));
    InMux I__6193 (
            .O(N__32166),
            .I(N__32158));
    LocalMux I__6192 (
            .O(N__32163),
            .I(il_max_comp2_D2));
    LocalMux I__6191 (
            .O(N__32158),
            .I(il_max_comp2_D2));
    InMux I__6190 (
            .O(N__32153),
            .I(N__32145));
    InMux I__6189 (
            .O(N__32152),
            .I(N__32145));
    InMux I__6188 (
            .O(N__32151),
            .I(N__32140));
    InMux I__6187 (
            .O(N__32150),
            .I(N__32140));
    LocalMux I__6186 (
            .O(N__32145),
            .I(\phase_controller_slave.stateZ0Z_3 ));
    LocalMux I__6185 (
            .O(N__32140),
            .I(\phase_controller_slave.stateZ0Z_3 ));
    CEMux I__6184 (
            .O(N__32135),
            .I(N__32130));
    CEMux I__6183 (
            .O(N__32134),
            .I(N__32127));
    CEMux I__6182 (
            .O(N__32133),
            .I(N__32123));
    LocalMux I__6181 (
            .O(N__32130),
            .I(N__32120));
    LocalMux I__6180 (
            .O(N__32127),
            .I(N__32117));
    CEMux I__6179 (
            .O(N__32126),
            .I(N__32114));
    LocalMux I__6178 (
            .O(N__32123),
            .I(N__32111));
    Span4Mux_v I__6177 (
            .O(N__32120),
            .I(N__32106));
    Span4Mux_v I__6176 (
            .O(N__32117),
            .I(N__32106));
    LocalMux I__6175 (
            .O(N__32114),
            .I(N__32103));
    Span4Mux_v I__6174 (
            .O(N__32111),
            .I(N__32098));
    Span4Mux_h I__6173 (
            .O(N__32106),
            .I(N__32098));
    Span4Mux_h I__6172 (
            .O(N__32103),
            .I(N__32095));
    Odrv4 I__6171 (
            .O(N__32098),
            .I(\current_shift_inst.timer_phase.N_192_i ));
    Odrv4 I__6170 (
            .O(N__32095),
            .I(\current_shift_inst.timer_phase.N_192_i ));
    InMux I__6169 (
            .O(N__32090),
            .I(N__32056));
    InMux I__6168 (
            .O(N__32089),
            .I(N__32056));
    InMux I__6167 (
            .O(N__32088),
            .I(N__32047));
    InMux I__6166 (
            .O(N__32087),
            .I(N__32047));
    InMux I__6165 (
            .O(N__32086),
            .I(N__32047));
    InMux I__6164 (
            .O(N__32085),
            .I(N__32047));
    InMux I__6163 (
            .O(N__32084),
            .I(N__32038));
    InMux I__6162 (
            .O(N__32083),
            .I(N__32038));
    InMux I__6161 (
            .O(N__32082),
            .I(N__32038));
    InMux I__6160 (
            .O(N__32081),
            .I(N__32038));
    InMux I__6159 (
            .O(N__32080),
            .I(N__32029));
    InMux I__6158 (
            .O(N__32079),
            .I(N__32029));
    InMux I__6157 (
            .O(N__32078),
            .I(N__32029));
    InMux I__6156 (
            .O(N__32077),
            .I(N__32029));
    InMux I__6155 (
            .O(N__32076),
            .I(N__32020));
    InMux I__6154 (
            .O(N__32075),
            .I(N__32020));
    InMux I__6153 (
            .O(N__32074),
            .I(N__32020));
    InMux I__6152 (
            .O(N__32073),
            .I(N__32020));
    InMux I__6151 (
            .O(N__32072),
            .I(N__32011));
    InMux I__6150 (
            .O(N__32071),
            .I(N__32011));
    InMux I__6149 (
            .O(N__32070),
            .I(N__32011));
    InMux I__6148 (
            .O(N__32069),
            .I(N__32011));
    InMux I__6147 (
            .O(N__32068),
            .I(N__32002));
    InMux I__6146 (
            .O(N__32067),
            .I(N__32002));
    InMux I__6145 (
            .O(N__32066),
            .I(N__32002));
    InMux I__6144 (
            .O(N__32065),
            .I(N__32002));
    InMux I__6143 (
            .O(N__32064),
            .I(N__31993));
    InMux I__6142 (
            .O(N__32063),
            .I(N__31993));
    InMux I__6141 (
            .O(N__32062),
            .I(N__31993));
    InMux I__6140 (
            .O(N__32061),
            .I(N__31993));
    LocalMux I__6139 (
            .O(N__32056),
            .I(N__31988));
    LocalMux I__6138 (
            .O(N__32047),
            .I(N__31988));
    LocalMux I__6137 (
            .O(N__32038),
            .I(N__31983));
    LocalMux I__6136 (
            .O(N__32029),
            .I(N__31983));
    LocalMux I__6135 (
            .O(N__32020),
            .I(N__31978));
    LocalMux I__6134 (
            .O(N__32011),
            .I(N__31978));
    LocalMux I__6133 (
            .O(N__32002),
            .I(N__31973));
    LocalMux I__6132 (
            .O(N__31993),
            .I(N__31973));
    Span4Mux_h I__6131 (
            .O(N__31988),
            .I(N__31970));
    Span4Mux_h I__6130 (
            .O(N__31983),
            .I(N__31967));
    Span4Mux_h I__6129 (
            .O(N__31978),
            .I(N__31964));
    Odrv4 I__6128 (
            .O(N__31973),
            .I(\current_shift_inst.timer_phase.running_i ));
    Odrv4 I__6127 (
            .O(N__31970),
            .I(\current_shift_inst.timer_phase.running_i ));
    Odrv4 I__6126 (
            .O(N__31967),
            .I(\current_shift_inst.timer_phase.running_i ));
    Odrv4 I__6125 (
            .O(N__31964),
            .I(\current_shift_inst.timer_phase.running_i ));
    InMux I__6124 (
            .O(N__31955),
            .I(N__31952));
    LocalMux I__6123 (
            .O(N__31952),
            .I(N__31949));
    Glb2LocalMux I__6122 (
            .O(N__31949),
            .I(N__31946));
    GlobalMux I__6121 (
            .O(N__31946),
            .I(clk_12mhz));
    IoInMux I__6120 (
            .O(N__31943),
            .I(N__31940));
    LocalMux I__6119 (
            .O(N__31940),
            .I(N__31937));
    Span12Mux_s0_v I__6118 (
            .O(N__31937),
            .I(N__31934));
    Odrv12 I__6117 (
            .O(N__31934),
            .I(GB_BUFFER_clk_12mhz_THRU_CO));
    CascadeMux I__6116 (
            .O(N__31931),
            .I(N__31928));
    InMux I__6115 (
            .O(N__31928),
            .I(N__31925));
    LocalMux I__6114 (
            .O(N__31925),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1Z0Z_6 ));
    CascadeMux I__6113 (
            .O(N__31922),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1Z0Z_6_cascade_ ));
    CascadeMux I__6112 (
            .O(N__31919),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6_cascade_ ));
    CascadeMux I__6111 (
            .O(N__31916),
            .I(\phase_controller_slave.start_timer_hc_0_sqmuxa_cascade_ ));
    IoInMux I__6110 (
            .O(N__31913),
            .I(N__31910));
    LocalMux I__6109 (
            .O(N__31910),
            .I(N__31907));
    IoSpan4Mux I__6108 (
            .O(N__31907),
            .I(N__31904));
    Span4Mux_s3_v I__6107 (
            .O(N__31904),
            .I(N__31900));
    InMux I__6106 (
            .O(N__31903),
            .I(N__31897));
    Span4Mux_v I__6105 (
            .O(N__31900),
            .I(N__31894));
    LocalMux I__6104 (
            .O(N__31897),
            .I(N__31891));
    Odrv4 I__6103 (
            .O(N__31894),
            .I(s3_phy_c));
    Odrv12 I__6102 (
            .O(N__31891),
            .I(s3_phy_c));
    CascadeMux I__6101 (
            .O(N__31886),
            .I(N__31883));
    InMux I__6100 (
            .O(N__31883),
            .I(N__31880));
    LocalMux I__6099 (
            .O(N__31880),
            .I(N__31877));
    Span4Mux_h I__6098 (
            .O(N__31877),
            .I(N__31874));
    Odrv4 I__6097 (
            .O(N__31874),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI1C4K_24 ));
    CascadeMux I__6096 (
            .O(N__31871),
            .I(N__31868));
    InMux I__6095 (
            .O(N__31868),
            .I(N__31863));
    InMux I__6094 (
            .O(N__31867),
            .I(N__31860));
    InMux I__6093 (
            .O(N__31866),
            .I(N__31856));
    LocalMux I__6092 (
            .O(N__31863),
            .I(N__31853));
    LocalMux I__6091 (
            .O(N__31860),
            .I(N__31850));
    InMux I__6090 (
            .O(N__31859),
            .I(N__31847));
    LocalMux I__6089 (
            .O(N__31856),
            .I(N__31842));
    Span12Mux_h I__6088 (
            .O(N__31853),
            .I(N__31842));
    Span4Mux_h I__6087 (
            .O(N__31850),
            .I(N__31837));
    LocalMux I__6086 (
            .O(N__31847),
            .I(N__31837));
    Odrv12 I__6085 (
            .O(N__31842),
            .I(\current_shift_inst.elapsed_time_ns_phase_26 ));
    Odrv4 I__6084 (
            .O(N__31837),
            .I(\current_shift_inst.elapsed_time_ns_phase_26 ));
    CascadeMux I__6083 (
            .O(N__31832),
            .I(N__31829));
    InMux I__6082 (
            .O(N__31829),
            .I(N__31826));
    LocalMux I__6081 (
            .O(N__31826),
            .I(N__31820));
    InMux I__6080 (
            .O(N__31825),
            .I(N__31817));
    CascadeMux I__6079 (
            .O(N__31824),
            .I(N__31814));
    InMux I__6078 (
            .O(N__31823),
            .I(N__31811));
    Span4Mux_h I__6077 (
            .O(N__31820),
            .I(N__31806));
    LocalMux I__6076 (
            .O(N__31817),
            .I(N__31806));
    InMux I__6075 (
            .O(N__31814),
            .I(N__31803));
    LocalMux I__6074 (
            .O(N__31811),
            .I(\current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0 ));
    Odrv4 I__6073 (
            .O(N__31806),
            .I(\current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0 ));
    LocalMux I__6072 (
            .O(N__31803),
            .I(\current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0 ));
    InMux I__6071 (
            .O(N__31796),
            .I(N__31793));
    LocalMux I__6070 (
            .O(N__31793),
            .I(N__31790));
    Span4Mux_h I__6069 (
            .O(N__31790),
            .I(N__31787));
    Odrv4 I__6068 (
            .O(N__31787),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIB4C81_25 ));
    InMux I__6067 (
            .O(N__31784),
            .I(N__31779));
    InMux I__6066 (
            .O(N__31783),
            .I(N__31774));
    InMux I__6065 (
            .O(N__31782),
            .I(N__31774));
    LocalMux I__6064 (
            .O(N__31779),
            .I(N__31769));
    LocalMux I__6063 (
            .O(N__31774),
            .I(N__31769));
    Span4Mux_h I__6062 (
            .O(N__31769),
            .I(N__31765));
    InMux I__6061 (
            .O(N__31768),
            .I(N__31762));
    Span4Mux_v I__6060 (
            .O(N__31765),
            .I(N__31759));
    LocalMux I__6059 (
            .O(N__31762),
            .I(N__31756));
    Odrv4 I__6058 (
            .O(N__31759),
            .I(\current_shift_inst.elapsed_time_ns_phase_25 ));
    Odrv4 I__6057 (
            .O(N__31756),
            .I(\current_shift_inst.elapsed_time_ns_phase_25 ));
    InMux I__6056 (
            .O(N__31751),
            .I(N__31743));
    InMux I__6055 (
            .O(N__31750),
            .I(N__31743));
    InMux I__6054 (
            .O(N__31749),
            .I(N__31740));
    InMux I__6053 (
            .O(N__31748),
            .I(N__31737));
    LocalMux I__6052 (
            .O(N__31743),
            .I(\current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0 ));
    LocalMux I__6051 (
            .O(N__31740),
            .I(\current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0 ));
    LocalMux I__6050 (
            .O(N__31737),
            .I(\current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0 ));
    CascadeMux I__6049 (
            .O(N__31730),
            .I(N__31727));
    InMux I__6048 (
            .O(N__31727),
            .I(N__31724));
    LocalMux I__6047 (
            .O(N__31724),
            .I(N__31721));
    Span4Mux_v I__6046 (
            .O(N__31721),
            .I(N__31718));
    Span4Mux_h I__6045 (
            .O(N__31718),
            .I(N__31715));
    Odrv4 I__6044 (
            .O(N__31715),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI4G5K_25 ));
    InMux I__6043 (
            .O(N__31712),
            .I(N__31709));
    LocalMux I__6042 (
            .O(N__31709),
            .I(N__31706));
    Span4Mux_v I__6041 (
            .O(N__31706),
            .I(N__31701));
    InMux I__6040 (
            .O(N__31705),
            .I(N__31698));
    InMux I__6039 (
            .O(N__31704),
            .I(N__31695));
    Span4Mux_h I__6038 (
            .O(N__31701),
            .I(N__31692));
    LocalMux I__6037 (
            .O(N__31698),
            .I(N__31689));
    LocalMux I__6036 (
            .O(N__31695),
            .I(N__31686));
    Odrv4 I__6035 (
            .O(N__31692),
            .I(\current_shift_inst.elapsed_time_ns_phase_29 ));
    Odrv12 I__6034 (
            .O(N__31689),
            .I(\current_shift_inst.elapsed_time_ns_phase_29 ));
    Odrv4 I__6033 (
            .O(N__31686),
            .I(\current_shift_inst.elapsed_time_ns_phase_29 ));
    InMux I__6032 (
            .O(N__31679),
            .I(N__31676));
    LocalMux I__6031 (
            .O(N__31676),
            .I(N__31672));
    InMux I__6030 (
            .O(N__31675),
            .I(N__31668));
    Span4Mux_h I__6029 (
            .O(N__31672),
            .I(N__31665));
    InMux I__6028 (
            .O(N__31671),
            .I(N__31662));
    LocalMux I__6027 (
            .O(N__31668),
            .I(\current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0 ));
    Odrv4 I__6026 (
            .O(N__31665),
            .I(\current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0 ));
    LocalMux I__6025 (
            .O(N__31662),
            .I(\current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0 ));
    InMux I__6024 (
            .O(N__31655),
            .I(N__31651));
    CascadeMux I__6023 (
            .O(N__31654),
            .I(N__31648));
    LocalMux I__6022 (
            .O(N__31651),
            .I(N__31645));
    InMux I__6021 (
            .O(N__31648),
            .I(N__31642));
    Span4Mux_v I__6020 (
            .O(N__31645),
            .I(N__31639));
    LocalMux I__6019 (
            .O(N__31642),
            .I(N__31636));
    Span4Mux_h I__6018 (
            .O(N__31639),
            .I(N__31631));
    Span4Mux_v I__6017 (
            .O(N__31636),
            .I(N__31631));
    Odrv4 I__6016 (
            .O(N__31631),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI7OAK_29 ));
    InMux I__6015 (
            .O(N__31628),
            .I(N__31623));
    InMux I__6014 (
            .O(N__31627),
            .I(N__31617));
    InMux I__6013 (
            .O(N__31626),
            .I(N__31617));
    LocalMux I__6012 (
            .O(N__31623),
            .I(N__31614));
    InMux I__6011 (
            .O(N__31622),
            .I(N__31611));
    LocalMux I__6010 (
            .O(N__31617),
            .I(N__31608));
    Span4Mux_v I__6009 (
            .O(N__31614),
            .I(N__31603));
    LocalMux I__6008 (
            .O(N__31611),
            .I(N__31603));
    Span12Mux_v I__6007 (
            .O(N__31608),
            .I(N__31600));
    Span4Mux_v I__6006 (
            .O(N__31603),
            .I(N__31597));
    Odrv12 I__6005 (
            .O(N__31600),
            .I(\current_shift_inst.elapsed_time_ns_phase_24 ));
    Odrv4 I__6004 (
            .O(N__31597),
            .I(\current_shift_inst.elapsed_time_ns_phase_24 ));
    InMux I__6003 (
            .O(N__31592),
            .I(N__31589));
    LocalMux I__6002 (
            .O(N__31589),
            .I(N__31584));
    InMux I__6001 (
            .O(N__31588),
            .I(N__31581));
    InMux I__6000 (
            .O(N__31587),
            .I(N__31578));
    Span4Mux_h I__5999 (
            .O(N__31584),
            .I(N__31573));
    LocalMux I__5998 (
            .O(N__31581),
            .I(N__31573));
    LocalMux I__5997 (
            .O(N__31578),
            .I(N__31569));
    Span4Mux_v I__5996 (
            .O(N__31573),
            .I(N__31566));
    InMux I__5995 (
            .O(N__31572),
            .I(N__31563));
    Odrv4 I__5994 (
            .O(N__31569),
            .I(\current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0 ));
    Odrv4 I__5993 (
            .O(N__31566),
            .I(\current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0 ));
    LocalMux I__5992 (
            .O(N__31563),
            .I(\current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0 ));
    CascadeMux I__5991 (
            .O(N__31556),
            .I(N__31553));
    InMux I__5990 (
            .O(N__31553),
            .I(N__31550));
    LocalMux I__5989 (
            .O(N__31550),
            .I(N__31545));
    InMux I__5988 (
            .O(N__31549),
            .I(N__31541));
    InMux I__5987 (
            .O(N__31548),
            .I(N__31538));
    Span4Mux_v I__5986 (
            .O(N__31545),
            .I(N__31535));
    InMux I__5985 (
            .O(N__31544),
            .I(N__31532));
    LocalMux I__5984 (
            .O(N__31541),
            .I(N__31529));
    LocalMux I__5983 (
            .O(N__31538),
            .I(N__31526));
    Span4Mux_h I__5982 (
            .O(N__31535),
            .I(N__31521));
    LocalMux I__5981 (
            .O(N__31532),
            .I(N__31521));
    Span4Mux_v I__5980 (
            .O(N__31529),
            .I(N__31518));
    Span4Mux_v I__5979 (
            .O(N__31526),
            .I(N__31515));
    Odrv4 I__5978 (
            .O(N__31521),
            .I(\current_shift_inst.elapsed_time_ns_phase_23 ));
    Odrv4 I__5977 (
            .O(N__31518),
            .I(\current_shift_inst.elapsed_time_ns_phase_23 ));
    Odrv4 I__5976 (
            .O(N__31515),
            .I(\current_shift_inst.elapsed_time_ns_phase_23 ));
    CascadeMux I__5975 (
            .O(N__31508),
            .I(N__31504));
    CascadeMux I__5974 (
            .O(N__31507),
            .I(N__31499));
    InMux I__5973 (
            .O(N__31504),
            .I(N__31496));
    InMux I__5972 (
            .O(N__31503),
            .I(N__31491));
    InMux I__5971 (
            .O(N__31502),
            .I(N__31491));
    InMux I__5970 (
            .O(N__31499),
            .I(N__31488));
    LocalMux I__5969 (
            .O(N__31496),
            .I(\current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0 ));
    LocalMux I__5968 (
            .O(N__31491),
            .I(\current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0 ));
    LocalMux I__5967 (
            .O(N__31488),
            .I(\current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0 ));
    InMux I__5966 (
            .O(N__31481),
            .I(N__31478));
    LocalMux I__5965 (
            .O(N__31478),
            .I(N__31475));
    Span4Mux_h I__5964 (
            .O(N__31475),
            .I(N__31472));
    Odrv4 I__5963 (
            .O(N__31472),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIVJ781_23 ));
    CascadeMux I__5962 (
            .O(N__31469),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3_cascade_ ));
    InMux I__5961 (
            .O(N__31466),
            .I(N__31463));
    LocalMux I__5960 (
            .O(N__31463),
            .I(\current_shift_inst.un4_control_input_axb_27 ));
    InMux I__5959 (
            .O(N__31460),
            .I(N__31457));
    LocalMux I__5958 (
            .O(N__31457),
            .I(\current_shift_inst.un4_control_input_axb_30 ));
    InMux I__5957 (
            .O(N__31454),
            .I(N__31451));
    LocalMux I__5956 (
            .O(N__31451),
            .I(\current_shift_inst.un4_control_input_axb_21 ));
    InMux I__5955 (
            .O(N__31448),
            .I(N__31445));
    LocalMux I__5954 (
            .O(N__31445),
            .I(\current_shift_inst.un4_control_input_axb_25 ));
    InMux I__5953 (
            .O(N__31442),
            .I(N__31439));
    LocalMux I__5952 (
            .O(N__31439),
            .I(\current_shift_inst.un4_control_input_axb_20 ));
    InMux I__5951 (
            .O(N__31436),
            .I(N__31432));
    InMux I__5950 (
            .O(N__31435),
            .I(N__31429));
    LocalMux I__5949 (
            .O(N__31432),
            .I(N__31426));
    LocalMux I__5948 (
            .O(N__31429),
            .I(N__31423));
    Odrv4 I__5947 (
            .O(N__31426),
            .I(\current_shift_inst.z_31 ));
    Odrv4 I__5946 (
            .O(N__31423),
            .I(\current_shift_inst.z_31 ));
    InMux I__5945 (
            .O(N__31418),
            .I(N__31414));
    CascadeMux I__5944 (
            .O(N__31417),
            .I(N__31411));
    LocalMux I__5943 (
            .O(N__31414),
            .I(N__31408));
    InMux I__5942 (
            .O(N__31411),
            .I(N__31405));
    Sp12to4 I__5941 (
            .O(N__31408),
            .I(N__31400));
    LocalMux I__5940 (
            .O(N__31405),
            .I(N__31400));
    Odrv12 I__5939 (
            .O(N__31400),
            .I(\current_shift_inst.z_i_31 ));
    InMux I__5938 (
            .O(N__31397),
            .I(N__31394));
    LocalMux I__5937 (
            .O(N__31394),
            .I(\current_shift_inst.un4_control_input_axb_28 ));
    InMux I__5936 (
            .O(N__31391),
            .I(N__31388));
    LocalMux I__5935 (
            .O(N__31388),
            .I(\current_shift_inst.un4_control_input_axb_11 ));
    CascadeMux I__5934 (
            .O(N__31385),
            .I(N__31382));
    InMux I__5933 (
            .O(N__31382),
            .I(N__31379));
    LocalMux I__5932 (
            .O(N__31379),
            .I(\current_shift_inst.un4_control_input_axb_19 ));
    InMux I__5931 (
            .O(N__31376),
            .I(N__31373));
    LocalMux I__5930 (
            .O(N__31373),
            .I(\current_shift_inst.un4_control_input_axb_10 ));
    InMux I__5929 (
            .O(N__31370),
            .I(N__31367));
    LocalMux I__5928 (
            .O(N__31367),
            .I(\current_shift_inst.un4_control_input_axb_12 ));
    InMux I__5927 (
            .O(N__31364),
            .I(N__31361));
    LocalMux I__5926 (
            .O(N__31361),
            .I(\current_shift_inst.un4_control_input_axb_14 ));
    InMux I__5925 (
            .O(N__31358),
            .I(N__31355));
    LocalMux I__5924 (
            .O(N__31355),
            .I(\current_shift_inst.un4_control_input_axb_18 ));
    InMux I__5923 (
            .O(N__31352),
            .I(N__31349));
    LocalMux I__5922 (
            .O(N__31349),
            .I(\current_shift_inst.un4_control_input_axb_29 ));
    InMux I__5921 (
            .O(N__31346),
            .I(N__31343));
    LocalMux I__5920 (
            .O(N__31343),
            .I(\current_shift_inst.un4_control_input_axb_22 ));
    InMux I__5919 (
            .O(N__31340),
            .I(N__31337));
    LocalMux I__5918 (
            .O(N__31337),
            .I(\current_shift_inst.un4_control_input_axb_26 ));
    InMux I__5917 (
            .O(N__31334),
            .I(N__31331));
    LocalMux I__5916 (
            .O(N__31331),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_1 ));
    InMux I__5915 (
            .O(N__31328),
            .I(N__31325));
    LocalMux I__5914 (
            .O(N__31325),
            .I(\current_shift_inst.un4_control_input_axb_1 ));
    InMux I__5913 (
            .O(N__31322),
            .I(N__31319));
    LocalMux I__5912 (
            .O(N__31319),
            .I(\current_shift_inst.timer_s1.elapsed_time_ns_s1_2 ));
    InMux I__5911 (
            .O(N__31316),
            .I(N__31313));
    LocalMux I__5910 (
            .O(N__31313),
            .I(\current_shift_inst.un4_control_input_axb_2 ));
    InMux I__5909 (
            .O(N__31310),
            .I(N__31307));
    LocalMux I__5908 (
            .O(N__31307),
            .I(\current_shift_inst.un4_control_input_axb_24 ));
    InMux I__5907 (
            .O(N__31304),
            .I(N__31301));
    LocalMux I__5906 (
            .O(N__31301),
            .I(\current_shift_inst.un4_control_input_axb_15 ));
    InMux I__5905 (
            .O(N__31298),
            .I(N__31295));
    LocalMux I__5904 (
            .O(N__31295),
            .I(N__31292));
    Odrv4 I__5903 (
            .O(N__31292),
            .I(\current_shift_inst.un4_control_input_axb_5 ));
    CascadeMux I__5902 (
            .O(N__31289),
            .I(N__31286));
    InMux I__5901 (
            .O(N__31286),
            .I(N__31283));
    LocalMux I__5900 (
            .O(N__31283),
            .I(N__31280));
    Odrv4 I__5899 (
            .O(N__31280),
            .I(\current_shift_inst.un4_control_input_axb_6 ));
    InMux I__5898 (
            .O(N__31277),
            .I(N__31274));
    LocalMux I__5897 (
            .O(N__31274),
            .I(N__31271));
    Odrv4 I__5896 (
            .O(N__31271),
            .I(\current_shift_inst.un4_control_input_axb_7 ));
    CascadeMux I__5895 (
            .O(N__31268),
            .I(N__31265));
    InMux I__5894 (
            .O(N__31265),
            .I(N__31262));
    LocalMux I__5893 (
            .O(N__31262),
            .I(N__31259));
    Odrv12 I__5892 (
            .O(N__31259),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ));
    CascadeMux I__5891 (
            .O(N__31256),
            .I(N__31253));
    InMux I__5890 (
            .O(N__31253),
            .I(N__31250));
    LocalMux I__5889 (
            .O(N__31250),
            .I(N__31247));
    Odrv12 I__5888 (
            .O(N__31247),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ));
    CascadeMux I__5887 (
            .O(N__31244),
            .I(N__31241));
    InMux I__5886 (
            .O(N__31241),
            .I(N__31238));
    LocalMux I__5885 (
            .O(N__31238),
            .I(N__31235));
    Span4Mux_h I__5884 (
            .O(N__31235),
            .I(N__31232));
    Odrv4 I__5883 (
            .O(N__31232),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ));
    CEMux I__5882 (
            .O(N__31229),
            .I(N__31221));
    CEMux I__5881 (
            .O(N__31228),
            .I(N__31218));
    CEMux I__5880 (
            .O(N__31227),
            .I(N__31215));
    CEMux I__5879 (
            .O(N__31226),
            .I(N__31212));
    CEMux I__5878 (
            .O(N__31225),
            .I(N__31209));
    CEMux I__5877 (
            .O(N__31224),
            .I(N__31206));
    LocalMux I__5876 (
            .O(N__31221),
            .I(N__31203));
    LocalMux I__5875 (
            .O(N__31218),
            .I(N__31200));
    LocalMux I__5874 (
            .O(N__31215),
            .I(N__31197));
    LocalMux I__5873 (
            .O(N__31212),
            .I(N__31194));
    LocalMux I__5872 (
            .O(N__31209),
            .I(N__31191));
    LocalMux I__5871 (
            .O(N__31206),
            .I(N__31188));
    Span4Mux_h I__5870 (
            .O(N__31203),
            .I(N__31185));
    Span4Mux_h I__5869 (
            .O(N__31200),
            .I(N__31180));
    Span4Mux_v I__5868 (
            .O(N__31197),
            .I(N__31180));
    Span4Mux_h I__5867 (
            .O(N__31194),
            .I(N__31177));
    Span4Mux_h I__5866 (
            .O(N__31191),
            .I(N__31174));
    Odrv12 I__5865 (
            .O(N__31188),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ));
    Odrv4 I__5864 (
            .O(N__31185),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ));
    Odrv4 I__5863 (
            .O(N__31180),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ));
    Odrv4 I__5862 (
            .O(N__31177),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ));
    Odrv4 I__5861 (
            .O(N__31174),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ));
    CascadeMux I__5860 (
            .O(N__31163),
            .I(N__31160));
    InMux I__5859 (
            .O(N__31160),
            .I(N__31157));
    LocalMux I__5858 (
            .O(N__31157),
            .I(\current_shift_inst.un4_control_input_axb_3 ));
    InMux I__5857 (
            .O(N__31154),
            .I(N__31151));
    LocalMux I__5856 (
            .O(N__31151),
            .I(\current_shift_inst.un4_control_input_axb_4 ));
    InMux I__5855 (
            .O(N__31148),
            .I(N__31145));
    LocalMux I__5854 (
            .O(N__31145),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9 ));
    InMux I__5853 (
            .O(N__31142),
            .I(N__31139));
    LocalMux I__5852 (
            .O(N__31139),
            .I(N__31135));
    InMux I__5851 (
            .O(N__31138),
            .I(N__31132));
    Span4Mux_v I__5850 (
            .O(N__31135),
            .I(N__31129));
    LocalMux I__5849 (
            .O(N__31132),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    Odrv4 I__5848 (
            .O(N__31129),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    CascadeMux I__5847 (
            .O(N__31124),
            .I(\phase_controller_inst1.start_timer_hc_0_sqmuxa_cascade_ ));
    InMux I__5846 (
            .O(N__31121),
            .I(N__31118));
    LocalMux I__5845 (
            .O(N__31118),
            .I(\phase_controller_inst1.N_88 ));
    InMux I__5844 (
            .O(N__31115),
            .I(N__31112));
    LocalMux I__5843 (
            .O(N__31112),
            .I(N__31107));
    InMux I__5842 (
            .O(N__31111),
            .I(N__31101));
    InMux I__5841 (
            .O(N__31110),
            .I(N__31101));
    Span4Mux_h I__5840 (
            .O(N__31107),
            .I(N__31098));
    InMux I__5839 (
            .O(N__31106),
            .I(N__31095));
    LocalMux I__5838 (
            .O(N__31101),
            .I(N__31092));
    Odrv4 I__5837 (
            .O(N__31098),
            .I(\phase_controller_inst1.hc_time_passed ));
    LocalMux I__5836 (
            .O(N__31095),
            .I(\phase_controller_inst1.hc_time_passed ));
    Odrv4 I__5835 (
            .O(N__31092),
            .I(\phase_controller_inst1.hc_time_passed ));
    InMux I__5834 (
            .O(N__31085),
            .I(N__31082));
    LocalMux I__5833 (
            .O(N__31082),
            .I(N__31079));
    Odrv4 I__5832 (
            .O(N__31079),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIDR081_20 ));
    CascadeMux I__5831 (
            .O(N__31076),
            .I(N__31073));
    InMux I__5830 (
            .O(N__31073),
            .I(N__31067));
    InMux I__5829 (
            .O(N__31072),
            .I(N__31062));
    InMux I__5828 (
            .O(N__31071),
            .I(N__31062));
    CascadeMux I__5827 (
            .O(N__31070),
            .I(N__31059));
    LocalMux I__5826 (
            .O(N__31067),
            .I(N__31054));
    LocalMux I__5825 (
            .O(N__31062),
            .I(N__31054));
    InMux I__5824 (
            .O(N__31059),
            .I(N__31051));
    Odrv4 I__5823 (
            .O(N__31054),
            .I(\current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0 ));
    LocalMux I__5822 (
            .O(N__31051),
            .I(\current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0 ));
    CascadeMux I__5821 (
            .O(N__31046),
            .I(N__31042));
    InMux I__5820 (
            .O(N__31045),
            .I(N__31034));
    InMux I__5819 (
            .O(N__31042),
            .I(N__31034));
    InMux I__5818 (
            .O(N__31041),
            .I(N__31034));
    LocalMux I__5817 (
            .O(N__31034),
            .I(N__31030));
    InMux I__5816 (
            .O(N__31033),
            .I(N__31027));
    Span4Mux_h I__5815 (
            .O(N__31030),
            .I(N__31022));
    LocalMux I__5814 (
            .O(N__31027),
            .I(N__31022));
    Odrv4 I__5813 (
            .O(N__31022),
            .I(\current_shift_inst.elapsed_time_ns_phase_20 ));
    CascadeMux I__5812 (
            .O(N__31019),
            .I(N__31016));
    InMux I__5811 (
            .O(N__31016),
            .I(N__31013));
    LocalMux I__5810 (
            .O(N__31013),
            .I(N__31010));
    Odrv4 I__5809 (
            .O(N__31010),
            .I(\current_shift_inst.elapsed_time_ns_1_RNILRVJ_20 ));
    CascadeMux I__5808 (
            .O(N__31007),
            .I(N__31004));
    InMux I__5807 (
            .O(N__31004),
            .I(N__30999));
    InMux I__5806 (
            .O(N__31003),
            .I(N__30996));
    InMux I__5805 (
            .O(N__31002),
            .I(N__30993));
    LocalMux I__5804 (
            .O(N__30999),
            .I(N__30989));
    LocalMux I__5803 (
            .O(N__30996),
            .I(N__30984));
    LocalMux I__5802 (
            .O(N__30993),
            .I(N__30984));
    InMux I__5801 (
            .O(N__30992),
            .I(N__30981));
    Span4Mux_v I__5800 (
            .O(N__30989),
            .I(N__30978));
    Span4Mux_h I__5799 (
            .O(N__30984),
            .I(N__30973));
    LocalMux I__5798 (
            .O(N__30981),
            .I(N__30973));
    Odrv4 I__5797 (
            .O(N__30978),
            .I(\current_shift_inst.elapsed_time_ns_phase_21 ));
    Odrv4 I__5796 (
            .O(N__30973),
            .I(\current_shift_inst.elapsed_time_ns_phase_21 ));
    InMux I__5795 (
            .O(N__30968),
            .I(N__30965));
    LocalMux I__5794 (
            .O(N__30965),
            .I(N__30960));
    InMux I__5793 (
            .O(N__30964),
            .I(N__30955));
    InMux I__5792 (
            .O(N__30963),
            .I(N__30955));
    Span4Mux_v I__5791 (
            .O(N__30960),
            .I(N__30951));
    LocalMux I__5790 (
            .O(N__30955),
            .I(N__30948));
    InMux I__5789 (
            .O(N__30954),
            .I(N__30945));
    Odrv4 I__5788 (
            .O(N__30951),
            .I(\current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0 ));
    Odrv4 I__5787 (
            .O(N__30948),
            .I(\current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0 ));
    LocalMux I__5786 (
            .O(N__30945),
            .I(\current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0 ));
    CascadeMux I__5785 (
            .O(N__30938),
            .I(N__30935));
    InMux I__5784 (
            .O(N__30935),
            .I(N__30932));
    LocalMux I__5783 (
            .O(N__30932),
            .I(N__30929));
    Span4Mux_h I__5782 (
            .O(N__30929),
            .I(N__30926));
    Odrv4 I__5781 (
            .O(N__30926),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIOV0K_21 ));
    CascadeMux I__5780 (
            .O(N__30923),
            .I(N__30920));
    InMux I__5779 (
            .O(N__30920),
            .I(N__30917));
    LocalMux I__5778 (
            .O(N__30917),
            .I(N__30914));
    Odrv12 I__5777 (
            .O(N__30914),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIU73K_23 ));
    CascadeMux I__5776 (
            .O(N__30911),
            .I(N__30908));
    InMux I__5775 (
            .O(N__30908),
            .I(N__30905));
    LocalMux I__5774 (
            .O(N__30905),
            .I(N__30902));
    Odrv12 I__5773 (
            .O(N__30902),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI7K6K_26 ));
    InMux I__5772 (
            .O(N__30899),
            .I(N__30896));
    LocalMux I__5771 (
            .O(N__30896),
            .I(N__30893));
    Span12Mux_v I__5770 (
            .O(N__30893),
            .I(N__30890));
    Span12Mux_v I__5769 (
            .O(N__30890),
            .I(N__30887));
    Odrv12 I__5768 (
            .O(N__30887),
            .I(il_max_comp2_D1));
    InMux I__5767 (
            .O(N__30884),
            .I(N__30880));
    InMux I__5766 (
            .O(N__30883),
            .I(N__30876));
    LocalMux I__5765 (
            .O(N__30880),
            .I(N__30873));
    InMux I__5764 (
            .O(N__30879),
            .I(N__30870));
    LocalMux I__5763 (
            .O(N__30876),
            .I(N__30864));
    Span4Mux_h I__5762 (
            .O(N__30873),
            .I(N__30864));
    LocalMux I__5761 (
            .O(N__30870),
            .I(N__30861));
    InMux I__5760 (
            .O(N__30869),
            .I(N__30858));
    Span4Mux_v I__5759 (
            .O(N__30864),
            .I(N__30855));
    Span4Mux_v I__5758 (
            .O(N__30861),
            .I(N__30852));
    LocalMux I__5757 (
            .O(N__30858),
            .I(N__30849));
    Odrv4 I__5756 (
            .O(N__30855),
            .I(\current_shift_inst.elapsed_time_ns_phase_28 ));
    Odrv4 I__5755 (
            .O(N__30852),
            .I(\current_shift_inst.elapsed_time_ns_phase_28 ));
    Odrv4 I__5754 (
            .O(N__30849),
            .I(\current_shift_inst.elapsed_time_ns_phase_28 ));
    CascadeMux I__5753 (
            .O(N__30842),
            .I(N__30839));
    InMux I__5752 (
            .O(N__30839),
            .I(N__30835));
    InMux I__5751 (
            .O(N__30838),
            .I(N__30832));
    LocalMux I__5750 (
            .O(N__30835),
            .I(N__30828));
    LocalMux I__5749 (
            .O(N__30832),
            .I(N__30824));
    CascadeMux I__5748 (
            .O(N__30831),
            .I(N__30821));
    Span4Mux_v I__5747 (
            .O(N__30828),
            .I(N__30818));
    InMux I__5746 (
            .O(N__30827),
            .I(N__30815));
    Span4Mux_h I__5745 (
            .O(N__30824),
            .I(N__30812));
    InMux I__5744 (
            .O(N__30821),
            .I(N__30809));
    Odrv4 I__5743 (
            .O(N__30818),
            .I(\current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0 ));
    LocalMux I__5742 (
            .O(N__30815),
            .I(\current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0 ));
    Odrv4 I__5741 (
            .O(N__30812),
            .I(\current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0 ));
    LocalMux I__5740 (
            .O(N__30809),
            .I(\current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0 ));
    CascadeMux I__5739 (
            .O(N__30800),
            .I(N__30797));
    InMux I__5738 (
            .O(N__30797),
            .I(N__30794));
    LocalMux I__5737 (
            .O(N__30794),
            .I(N__30791));
    Span4Mux_v I__5736 (
            .O(N__30791),
            .I(N__30788));
    Odrv4 I__5735 (
            .O(N__30788),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIDS8K_28 ));
    InMux I__5734 (
            .O(N__30785),
            .I(N__30782));
    LocalMux I__5733 (
            .O(N__30782),
            .I(N__30779));
    Span4Mux_h I__5732 (
            .O(N__30779),
            .I(N__30776));
    Odrv4 I__5731 (
            .O(N__30776),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5S981_24 ));
    CascadeMux I__5730 (
            .O(N__30773),
            .I(N__30768));
    InMux I__5729 (
            .O(N__30772),
            .I(N__30763));
    InMux I__5728 (
            .O(N__30771),
            .I(N__30763));
    InMux I__5727 (
            .O(N__30768),
            .I(N__30759));
    LocalMux I__5726 (
            .O(N__30763),
            .I(N__30756));
    InMux I__5725 (
            .O(N__30762),
            .I(N__30753));
    LocalMux I__5724 (
            .O(N__30759),
            .I(N__30750));
    Span4Mux_h I__5723 (
            .O(N__30756),
            .I(N__30745));
    LocalMux I__5722 (
            .O(N__30753),
            .I(N__30745));
    Odrv12 I__5721 (
            .O(N__30750),
            .I(\current_shift_inst.elapsed_time_ns_phase_11 ));
    Odrv4 I__5720 (
            .O(N__30745),
            .I(\current_shift_inst.elapsed_time_ns_phase_11 ));
    InMux I__5719 (
            .O(N__30740),
            .I(N__30730));
    InMux I__5718 (
            .O(N__30739),
            .I(N__30730));
    InMux I__5717 (
            .O(N__30738),
            .I(N__30730));
    CascadeMux I__5716 (
            .O(N__30737),
            .I(N__30727));
    LocalMux I__5715 (
            .O(N__30730),
            .I(N__30724));
    InMux I__5714 (
            .O(N__30727),
            .I(N__30721));
    Odrv4 I__5713 (
            .O(N__30724),
            .I(\current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0 ));
    LocalMux I__5712 (
            .O(N__30721),
            .I(\current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0 ));
    CascadeMux I__5711 (
            .O(N__30716),
            .I(N__30712));
    InMux I__5710 (
            .O(N__30715),
            .I(N__30709));
    InMux I__5709 (
            .O(N__30712),
            .I(N__30704));
    LocalMux I__5708 (
            .O(N__30709),
            .I(N__30701));
    InMux I__5707 (
            .O(N__30708),
            .I(N__30698));
    CascadeMux I__5706 (
            .O(N__30707),
            .I(N__30695));
    LocalMux I__5705 (
            .O(N__30704),
            .I(N__30688));
    Span4Mux_h I__5704 (
            .O(N__30701),
            .I(N__30688));
    LocalMux I__5703 (
            .O(N__30698),
            .I(N__30688));
    InMux I__5702 (
            .O(N__30695),
            .I(N__30685));
    Odrv4 I__5701 (
            .O(N__30688),
            .I(\current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0 ));
    LocalMux I__5700 (
            .O(N__30685),
            .I(\current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0 ));
    CascadeMux I__5699 (
            .O(N__30680),
            .I(N__30676));
    CascadeMux I__5698 (
            .O(N__30679),
            .I(N__30673));
    InMux I__5697 (
            .O(N__30676),
            .I(N__30669));
    InMux I__5696 (
            .O(N__30673),
            .I(N__30664));
    InMux I__5695 (
            .O(N__30672),
            .I(N__30664));
    LocalMux I__5694 (
            .O(N__30669),
            .I(N__30658));
    LocalMux I__5693 (
            .O(N__30664),
            .I(N__30658));
    InMux I__5692 (
            .O(N__30663),
            .I(N__30655));
    Span4Mux_h I__5691 (
            .O(N__30658),
            .I(N__30650));
    LocalMux I__5690 (
            .O(N__30655),
            .I(N__30650));
    Odrv4 I__5689 (
            .O(N__30650),
            .I(\current_shift_inst.elapsed_time_ns_phase_12 ));
    InMux I__5688 (
            .O(N__30647),
            .I(N__30644));
    LocalMux I__5687 (
            .O(N__30644),
            .I(N__30641));
    Odrv4 I__5686 (
            .O(N__30641),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIDLO51_11 ));
    InMux I__5685 (
            .O(N__30638),
            .I(N__30635));
    LocalMux I__5684 (
            .O(N__30635),
            .I(N__30632));
    Span4Mux_v I__5683 (
            .O(N__30632),
            .I(N__30627));
    InMux I__5682 (
            .O(N__30631),
            .I(N__30624));
    InMux I__5681 (
            .O(N__30630),
            .I(N__30621));
    Span4Mux_v I__5680 (
            .O(N__30627),
            .I(N__30618));
    LocalMux I__5679 (
            .O(N__30624),
            .I(N__30615));
    LocalMux I__5678 (
            .O(N__30621),
            .I(N__30612));
    Odrv4 I__5677 (
            .O(N__30618),
            .I(\current_shift_inst.elapsed_time_ns_phase_30 ));
    Odrv12 I__5676 (
            .O(N__30615),
            .I(\current_shift_inst.elapsed_time_ns_phase_30 ));
    Odrv4 I__5675 (
            .O(N__30612),
            .I(\current_shift_inst.elapsed_time_ns_phase_30 ));
    CascadeMux I__5674 (
            .O(N__30605),
            .I(N__30600));
    CascadeMux I__5673 (
            .O(N__30604),
            .I(N__30595));
    CascadeMux I__5672 (
            .O(N__30603),
            .I(N__30591));
    InMux I__5671 (
            .O(N__30600),
            .I(N__30587));
    InMux I__5670 (
            .O(N__30599),
            .I(N__30584));
    InMux I__5669 (
            .O(N__30598),
            .I(N__30575));
    InMux I__5668 (
            .O(N__30595),
            .I(N__30575));
    InMux I__5667 (
            .O(N__30594),
            .I(N__30575));
    InMux I__5666 (
            .O(N__30591),
            .I(N__30575));
    InMux I__5665 (
            .O(N__30590),
            .I(N__30571));
    LocalMux I__5664 (
            .O(N__30587),
            .I(N__30564));
    LocalMux I__5663 (
            .O(N__30584),
            .I(N__30564));
    LocalMux I__5662 (
            .O(N__30575),
            .I(N__30564));
    InMux I__5661 (
            .O(N__30574),
            .I(N__30561));
    LocalMux I__5660 (
            .O(N__30571),
            .I(N__30557));
    Span4Mux_h I__5659 (
            .O(N__30564),
            .I(N__30554));
    LocalMux I__5658 (
            .O(N__30561),
            .I(N__30551));
    InMux I__5657 (
            .O(N__30560),
            .I(N__30548));
    Span4Mux_v I__5656 (
            .O(N__30557),
            .I(N__30539));
    Span4Mux_h I__5655 (
            .O(N__30554),
            .I(N__30539));
    Span4Mux_h I__5654 (
            .O(N__30551),
            .I(N__30539));
    LocalMux I__5653 (
            .O(N__30548),
            .I(N__30539));
    Span4Mux_v I__5652 (
            .O(N__30539),
            .I(N__30536));
    Odrv4 I__5651 (
            .O(N__30536),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    CascadeMux I__5650 (
            .O(N__30533),
            .I(N__30530));
    InMux I__5649 (
            .O(N__30530),
            .I(N__30526));
    CascadeMux I__5648 (
            .O(N__30529),
            .I(N__30523));
    LocalMux I__5647 (
            .O(N__30526),
            .I(N__30520));
    InMux I__5646 (
            .O(N__30523),
            .I(N__30517));
    Span4Mux_h I__5645 (
            .O(N__30520),
            .I(N__30514));
    LocalMux I__5644 (
            .O(N__30517),
            .I(N__30511));
    Span4Mux_v I__5643 (
            .O(N__30514),
            .I(N__30508));
    Span4Mux_v I__5642 (
            .O(N__30511),
            .I(N__30505));
    Odrv4 I__5641 (
            .O(N__30508),
            .I(\current_shift_inst.elapsed_time_ns_phase_31 ));
    Odrv4 I__5640 (
            .O(N__30505),
            .I(\current_shift_inst.elapsed_time_ns_phase_31 ));
    InMux I__5639 (
            .O(N__30500),
            .I(N__30496));
    InMux I__5638 (
            .O(N__30499),
            .I(N__30493));
    LocalMux I__5637 (
            .O(N__30496),
            .I(N__30490));
    LocalMux I__5636 (
            .O(N__30493),
            .I(N__30484));
    Span4Mux_h I__5635 (
            .O(N__30490),
            .I(N__30484));
    InMux I__5634 (
            .O(N__30489),
            .I(N__30481));
    Odrv4 I__5633 (
            .O(N__30484),
            .I(\current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0 ));
    LocalMux I__5632 (
            .O(N__30481),
            .I(\current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0 ));
    InMux I__5631 (
            .O(N__30476),
            .I(N__30473));
    LocalMux I__5630 (
            .O(N__30473),
            .I(N__30470));
    Span4Mux_h I__5629 (
            .O(N__30470),
            .I(N__30467));
    Odrv4 I__5628 (
            .O(N__30467),
            .I(\current_shift_inst.un38_control_input_0_axb_31 ));
    InMux I__5627 (
            .O(N__30464),
            .I(N__30459));
    InMux I__5626 (
            .O(N__30463),
            .I(N__30456));
    InMux I__5625 (
            .O(N__30462),
            .I(N__30453));
    LocalMux I__5624 (
            .O(N__30459),
            .I(N__30449));
    LocalMux I__5623 (
            .O(N__30456),
            .I(N__30446));
    LocalMux I__5622 (
            .O(N__30453),
            .I(N__30443));
    InMux I__5621 (
            .O(N__30452),
            .I(N__30440));
    Span4Mux_h I__5620 (
            .O(N__30449),
            .I(N__30435));
    Span4Mux_v I__5619 (
            .O(N__30446),
            .I(N__30435));
    Span4Mux_v I__5618 (
            .O(N__30443),
            .I(N__30430));
    LocalMux I__5617 (
            .O(N__30440),
            .I(N__30430));
    Odrv4 I__5616 (
            .O(N__30435),
            .I(\current_shift_inst.elapsed_time_ns_phase_19 ));
    Odrv4 I__5615 (
            .O(N__30430),
            .I(\current_shift_inst.elapsed_time_ns_phase_19 ));
    CascadeMux I__5614 (
            .O(N__30425),
            .I(N__30421));
    InMux I__5613 (
            .O(N__30424),
            .I(N__30418));
    InMux I__5612 (
            .O(N__30421),
            .I(N__30413));
    LocalMux I__5611 (
            .O(N__30418),
            .I(N__30410));
    InMux I__5610 (
            .O(N__30417),
            .I(N__30407));
    CascadeMux I__5609 (
            .O(N__30416),
            .I(N__30404));
    LocalMux I__5608 (
            .O(N__30413),
            .I(N__30401));
    Span4Mux_v I__5607 (
            .O(N__30410),
            .I(N__30398));
    LocalMux I__5606 (
            .O(N__30407),
            .I(N__30395));
    InMux I__5605 (
            .O(N__30404),
            .I(N__30392));
    Odrv12 I__5604 (
            .O(N__30401),
            .I(\current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0 ));
    Odrv4 I__5603 (
            .O(N__30398),
            .I(\current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0 ));
    Odrv4 I__5602 (
            .O(N__30395),
            .I(\current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0 ));
    LocalMux I__5601 (
            .O(N__30392),
            .I(\current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0 ));
    InMux I__5600 (
            .O(N__30383),
            .I(N__30380));
    LocalMux I__5599 (
            .O(N__30380),
            .I(N__30377));
    Odrv12 I__5598 (
            .O(N__30377),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPC571_19 ));
    CascadeMux I__5597 (
            .O(N__30374),
            .I(N__30371));
    InMux I__5596 (
            .O(N__30371),
            .I(N__30368));
    LocalMux I__5595 (
            .O(N__30368),
            .I(N__30365));
    Span4Mux_h I__5594 (
            .O(N__30365),
            .I(N__30362));
    Odrv4 I__5593 (
            .O(N__30362),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI190J_15 ));
    InMux I__5592 (
            .O(N__30359),
            .I(N__30354));
    CascadeMux I__5591 (
            .O(N__30358),
            .I(N__30351));
    CascadeMux I__5590 (
            .O(N__30357),
            .I(N__30347));
    LocalMux I__5589 (
            .O(N__30354),
            .I(N__30344));
    InMux I__5588 (
            .O(N__30351),
            .I(N__30341));
    InMux I__5587 (
            .O(N__30350),
            .I(N__30338));
    InMux I__5586 (
            .O(N__30347),
            .I(N__30335));
    Span4Mux_v I__5585 (
            .O(N__30344),
            .I(N__30332));
    LocalMux I__5584 (
            .O(N__30341),
            .I(N__30325));
    LocalMux I__5583 (
            .O(N__30338),
            .I(N__30325));
    LocalMux I__5582 (
            .O(N__30335),
            .I(N__30325));
    Odrv4 I__5581 (
            .O(N__30332),
            .I(\current_shift_inst.elapsed_time_ns_phase_16 ));
    Odrv4 I__5580 (
            .O(N__30325),
            .I(\current_shift_inst.elapsed_time_ns_phase_16 ));
    InMux I__5579 (
            .O(N__30320),
            .I(N__30316));
    InMux I__5578 (
            .O(N__30319),
            .I(N__30313));
    LocalMux I__5577 (
            .O(N__30316),
            .I(N__30307));
    LocalMux I__5576 (
            .O(N__30313),
            .I(N__30307));
    InMux I__5575 (
            .O(N__30312),
            .I(N__30304));
    Span4Mux_v I__5574 (
            .O(N__30307),
            .I(N__30300));
    LocalMux I__5573 (
            .O(N__30304),
            .I(N__30297));
    InMux I__5572 (
            .O(N__30303),
            .I(N__30294));
    Odrv4 I__5571 (
            .O(N__30300),
            .I(\current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0 ));
    Odrv12 I__5570 (
            .O(N__30297),
            .I(\current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0 ));
    LocalMux I__5569 (
            .O(N__30294),
            .I(\current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0 ));
    InMux I__5568 (
            .O(N__30287),
            .I(N__30284));
    LocalMux I__5567 (
            .O(N__30284),
            .I(N__30281));
    Odrv4 I__5566 (
            .O(N__30281),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5M161_15 ));
    InMux I__5565 (
            .O(N__30278),
            .I(N__30275));
    LocalMux I__5564 (
            .O(N__30275),
            .I(N__30272));
    Span4Mux_h I__5563 (
            .O(N__30272),
            .I(N__30266));
    InMux I__5562 (
            .O(N__30271),
            .I(N__30263));
    InMux I__5561 (
            .O(N__30270),
            .I(N__30260));
    InMux I__5560 (
            .O(N__30269),
            .I(N__30257));
    Span4Mux_h I__5559 (
            .O(N__30266),
            .I(N__30254));
    LocalMux I__5558 (
            .O(N__30263),
            .I(N__30251));
    LocalMux I__5557 (
            .O(N__30260),
            .I(N__30246));
    LocalMux I__5556 (
            .O(N__30257),
            .I(N__30246));
    Odrv4 I__5555 (
            .O(N__30254),
            .I(\current_shift_inst.elapsed_time_ns_phase_14 ));
    Odrv12 I__5554 (
            .O(N__30251),
            .I(\current_shift_inst.elapsed_time_ns_phase_14 ));
    Odrv4 I__5553 (
            .O(N__30246),
            .I(\current_shift_inst.elapsed_time_ns_phase_14 ));
    CascadeMux I__5552 (
            .O(N__30239),
            .I(N__30236));
    InMux I__5551 (
            .O(N__30236),
            .I(N__30226));
    InMux I__5550 (
            .O(N__30235),
            .I(N__30226));
    InMux I__5549 (
            .O(N__30234),
            .I(N__30226));
    CascadeMux I__5548 (
            .O(N__30233),
            .I(N__30223));
    LocalMux I__5547 (
            .O(N__30226),
            .I(N__30220));
    InMux I__5546 (
            .O(N__30223),
            .I(N__30217));
    Odrv12 I__5545 (
            .O(N__30220),
            .I(\current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0 ));
    LocalMux I__5544 (
            .O(N__30217),
            .I(\current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0 ));
    CascadeMux I__5543 (
            .O(N__30212),
            .I(N__30208));
    InMux I__5542 (
            .O(N__30211),
            .I(N__30204));
    InMux I__5541 (
            .O(N__30208),
            .I(N__30201));
    InMux I__5540 (
            .O(N__30207),
            .I(N__30198));
    LocalMux I__5539 (
            .O(N__30204),
            .I(N__30194));
    LocalMux I__5538 (
            .O(N__30201),
            .I(N__30191));
    LocalMux I__5537 (
            .O(N__30198),
            .I(N__30188));
    CascadeMux I__5536 (
            .O(N__30197),
            .I(N__30185));
    Span4Mux_v I__5535 (
            .O(N__30194),
            .I(N__30182));
    Span4Mux_v I__5534 (
            .O(N__30191),
            .I(N__30177));
    Span4Mux_h I__5533 (
            .O(N__30188),
            .I(N__30177));
    InMux I__5532 (
            .O(N__30185),
            .I(N__30174));
    Odrv4 I__5531 (
            .O(N__30182),
            .I(\current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0 ));
    Odrv4 I__5530 (
            .O(N__30177),
            .I(\current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0 ));
    LocalMux I__5529 (
            .O(N__30174),
            .I(\current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0 ));
    InMux I__5528 (
            .O(N__30167),
            .I(N__30157));
    InMux I__5527 (
            .O(N__30166),
            .I(N__30157));
    InMux I__5526 (
            .O(N__30165),
            .I(N__30157));
    InMux I__5525 (
            .O(N__30164),
            .I(N__30154));
    LocalMux I__5524 (
            .O(N__30157),
            .I(N__30151));
    LocalMux I__5523 (
            .O(N__30154),
            .I(N__30148));
    Span4Mux_v I__5522 (
            .O(N__30151),
            .I(N__30145));
    Span4Mux_v I__5521 (
            .O(N__30148),
            .I(N__30142));
    Odrv4 I__5520 (
            .O(N__30145),
            .I(\current_shift_inst.elapsed_time_ns_phase_15 ));
    Odrv4 I__5519 (
            .O(N__30142),
            .I(\current_shift_inst.elapsed_time_ns_phase_15 ));
    InMux I__5518 (
            .O(N__30137),
            .I(N__30134));
    LocalMux I__5517 (
            .O(N__30134),
            .I(N__30131));
    Odrv4 I__5516 (
            .O(N__30131),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIVDV51_14 ));
    CascadeMux I__5515 (
            .O(N__30128),
            .I(N__30125));
    InMux I__5514 (
            .O(N__30125),
            .I(N__30122));
    LocalMux I__5513 (
            .O(N__30122),
            .I(N__30117));
    InMux I__5512 (
            .O(N__30121),
            .I(N__30112));
    InMux I__5511 (
            .O(N__30120),
            .I(N__30112));
    Span4Mux_h I__5510 (
            .O(N__30117),
            .I(N__30108));
    LocalMux I__5509 (
            .O(N__30112),
            .I(N__30105));
    CascadeMux I__5508 (
            .O(N__30111),
            .I(N__30102));
    Sp12to4 I__5507 (
            .O(N__30108),
            .I(N__30099));
    Span4Mux_h I__5506 (
            .O(N__30105),
            .I(N__30096));
    InMux I__5505 (
            .O(N__30102),
            .I(N__30093));
    Odrv12 I__5504 (
            .O(N__30099),
            .I(\current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0 ));
    Odrv4 I__5503 (
            .O(N__30096),
            .I(\current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0 ));
    LocalMux I__5502 (
            .O(N__30093),
            .I(\current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0 ));
    InMux I__5501 (
            .O(N__30086),
            .I(\current_shift_inst.un4_control_input_cry_27 ));
    InMux I__5500 (
            .O(N__30083),
            .I(\current_shift_inst.un4_control_input_cry_28 ));
    InMux I__5499 (
            .O(N__30080),
            .I(\current_shift_inst.un4_control_input_cry_29 ));
    InMux I__5498 (
            .O(N__30077),
            .I(\current_shift_inst.un4_control_input_cry_30 ));
    InMux I__5497 (
            .O(N__30074),
            .I(N__30070));
    InMux I__5496 (
            .O(N__30073),
            .I(N__30066));
    LocalMux I__5495 (
            .O(N__30070),
            .I(N__30062));
    InMux I__5494 (
            .O(N__30069),
            .I(N__30059));
    LocalMux I__5493 (
            .O(N__30066),
            .I(N__30056));
    InMux I__5492 (
            .O(N__30065),
            .I(N__30053));
    Span4Mux_h I__5491 (
            .O(N__30062),
            .I(N__30044));
    LocalMux I__5490 (
            .O(N__30059),
            .I(N__30044));
    Span4Mux_h I__5489 (
            .O(N__30056),
            .I(N__30044));
    LocalMux I__5488 (
            .O(N__30053),
            .I(N__30044));
    Odrv4 I__5487 (
            .O(N__30044),
            .I(\current_shift_inst.elapsed_time_ns_phase_9 ));
    CascadeMux I__5486 (
            .O(N__30041),
            .I(N__30038));
    InMux I__5485 (
            .O(N__30038),
            .I(N__30034));
    InMux I__5484 (
            .O(N__30037),
            .I(N__30031));
    LocalMux I__5483 (
            .O(N__30034),
            .I(N__30024));
    LocalMux I__5482 (
            .O(N__30031),
            .I(N__30024));
    InMux I__5481 (
            .O(N__30030),
            .I(N__30021));
    CascadeMux I__5480 (
            .O(N__30029),
            .I(N__30018));
    Span4Mux_v I__5479 (
            .O(N__30024),
            .I(N__30015));
    LocalMux I__5478 (
            .O(N__30021),
            .I(N__30012));
    InMux I__5477 (
            .O(N__30018),
            .I(N__30009));
    Odrv4 I__5476 (
            .O(N__30015),
            .I(\current_shift_inst.un4_control_input_cry_9_c_RNIALDJZ0 ));
    Odrv12 I__5475 (
            .O(N__30012),
            .I(\current_shift_inst.un4_control_input_cry_9_c_RNIALDJZ0 ));
    LocalMux I__5474 (
            .O(N__30009),
            .I(\current_shift_inst.un4_control_input_cry_9_c_RNIALDJZ0 ));
    InMux I__5473 (
            .O(N__30002),
            .I(N__29999));
    LocalMux I__5472 (
            .O(N__29999),
            .I(N__29996));
    Odrv12 I__5471 (
            .O(N__29996),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIO0U12_8 ));
    CascadeMux I__5470 (
            .O(N__29993),
            .I(N__29990));
    InMux I__5469 (
            .O(N__29990),
            .I(N__29987));
    LocalMux I__5468 (
            .O(N__29987),
            .I(N__29984));
    Odrv12 I__5467 (
            .O(N__29984),
            .I(\current_shift_inst.elapsed_time_ns_1_RNILORI_11 ));
    CascadeMux I__5466 (
            .O(N__29981),
            .I(N__29978));
    InMux I__5465 (
            .O(N__29978),
            .I(N__29975));
    LocalMux I__5464 (
            .O(N__29975),
            .I(N__29972));
    Odrv4 I__5463 (
            .O(N__29972),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIOSSI_12 ));
    InMux I__5462 (
            .O(N__29969),
            .I(N__29964));
    InMux I__5461 (
            .O(N__29968),
            .I(N__29961));
    InMux I__5460 (
            .O(N__29967),
            .I(N__29958));
    LocalMux I__5459 (
            .O(N__29964),
            .I(N__29952));
    LocalMux I__5458 (
            .O(N__29961),
            .I(N__29952));
    LocalMux I__5457 (
            .O(N__29958),
            .I(N__29949));
    InMux I__5456 (
            .O(N__29957),
            .I(N__29946));
    Span4Mux_v I__5455 (
            .O(N__29952),
            .I(N__29943));
    Span4Mux_h I__5454 (
            .O(N__29949),
            .I(N__29938));
    LocalMux I__5453 (
            .O(N__29946),
            .I(N__29938));
    Odrv4 I__5452 (
            .O(N__29943),
            .I(\current_shift_inst.elapsed_time_ns_phase_13 ));
    Odrv4 I__5451 (
            .O(N__29938),
            .I(\current_shift_inst.elapsed_time_ns_phase_13 ));
    CascadeMux I__5450 (
            .O(N__29933),
            .I(N__29930));
    InMux I__5449 (
            .O(N__29930),
            .I(N__29926));
    InMux I__5448 (
            .O(N__29929),
            .I(N__29922));
    LocalMux I__5447 (
            .O(N__29926),
            .I(N__29918));
    InMux I__5446 (
            .O(N__29925),
            .I(N__29915));
    LocalMux I__5445 (
            .O(N__29922),
            .I(N__29912));
    CascadeMux I__5444 (
            .O(N__29921),
            .I(N__29909));
    Span4Mux_h I__5443 (
            .O(N__29918),
            .I(N__29904));
    LocalMux I__5442 (
            .O(N__29915),
            .I(N__29904));
    Span4Mux_v I__5441 (
            .O(N__29912),
            .I(N__29901));
    InMux I__5440 (
            .O(N__29909),
            .I(N__29898));
    Odrv4 I__5439 (
            .O(N__29904),
            .I(\current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0 ));
    Odrv4 I__5438 (
            .O(N__29901),
            .I(\current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0 ));
    LocalMux I__5437 (
            .O(N__29898),
            .I(\current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0 ));
    InMux I__5436 (
            .O(N__29891),
            .I(N__29888));
    LocalMux I__5435 (
            .O(N__29888),
            .I(N__29885));
    Odrv12 I__5434 (
            .O(N__29885),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJTQ51_12 ));
    InMux I__5433 (
            .O(N__29882),
            .I(N__29877));
    InMux I__5432 (
            .O(N__29881),
            .I(N__29874));
    InMux I__5431 (
            .O(N__29880),
            .I(N__29870));
    LocalMux I__5430 (
            .O(N__29877),
            .I(N__29865));
    LocalMux I__5429 (
            .O(N__29874),
            .I(N__29865));
    InMux I__5428 (
            .O(N__29873),
            .I(N__29862));
    LocalMux I__5427 (
            .O(N__29870),
            .I(N__29859));
    Span4Mux_v I__5426 (
            .O(N__29865),
            .I(N__29856));
    LocalMux I__5425 (
            .O(N__29862),
            .I(N__29853));
    Odrv4 I__5424 (
            .O(N__29859),
            .I(\current_shift_inst.elapsed_time_ns_phase_8 ));
    Odrv4 I__5423 (
            .O(N__29856),
            .I(\current_shift_inst.elapsed_time_ns_phase_8 ));
    Odrv4 I__5422 (
            .O(N__29853),
            .I(\current_shift_inst.elapsed_time_ns_phase_8 ));
    InMux I__5421 (
            .O(N__29846),
            .I(N__29842));
    CascadeMux I__5420 (
            .O(N__29845),
            .I(N__29839));
    LocalMux I__5419 (
            .O(N__29842),
            .I(N__29834));
    InMux I__5418 (
            .O(N__29839),
            .I(N__29831));
    InMux I__5417 (
            .O(N__29838),
            .I(N__29828));
    CascadeMux I__5416 (
            .O(N__29837),
            .I(N__29825));
    Span4Mux_v I__5415 (
            .O(N__29834),
            .I(N__29822));
    LocalMux I__5414 (
            .O(N__29831),
            .I(N__29817));
    LocalMux I__5413 (
            .O(N__29828),
            .I(N__29817));
    InMux I__5412 (
            .O(N__29825),
            .I(N__29814));
    Odrv4 I__5411 (
            .O(N__29822),
            .I(\current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0 ));
    Odrv12 I__5410 (
            .O(N__29817),
            .I(\current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0 ));
    LocalMux I__5409 (
            .O(N__29814),
            .I(\current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0 ));
    CascadeMux I__5408 (
            .O(N__29807),
            .I(N__29804));
    InMux I__5407 (
            .O(N__29804),
            .I(N__29801));
    LocalMux I__5406 (
            .O(N__29801),
            .I(N__29798));
    Odrv4 I__5405 (
            .O(N__29798),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIN7DV_8 ));
    InMux I__5404 (
            .O(N__29795),
            .I(\current_shift_inst.un4_control_input_cry_18 ));
    InMux I__5403 (
            .O(N__29792),
            .I(\current_shift_inst.un4_control_input_cry_19 ));
    InMux I__5402 (
            .O(N__29789),
            .I(\current_shift_inst.un4_control_input_cry_20 ));
    InMux I__5401 (
            .O(N__29786),
            .I(\current_shift_inst.un4_control_input_cry_21 ));
    CascadeMux I__5400 (
            .O(N__29783),
            .I(N__29780));
    InMux I__5399 (
            .O(N__29780),
            .I(N__29771));
    InMux I__5398 (
            .O(N__29779),
            .I(N__29771));
    InMux I__5397 (
            .O(N__29778),
            .I(N__29771));
    LocalMux I__5396 (
            .O(N__29771),
            .I(N__29767));
    CascadeMux I__5395 (
            .O(N__29770),
            .I(N__29764));
    Span4Mux_v I__5394 (
            .O(N__29767),
            .I(N__29761));
    InMux I__5393 (
            .O(N__29764),
            .I(N__29758));
    Odrv4 I__5392 (
            .O(N__29761),
            .I(\current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0 ));
    LocalMux I__5391 (
            .O(N__29758),
            .I(\current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0 ));
    InMux I__5390 (
            .O(N__29753),
            .I(\current_shift_inst.un4_control_input_cry_22 ));
    InMux I__5389 (
            .O(N__29750),
            .I(\current_shift_inst.un4_control_input_cry_23 ));
    InMux I__5388 (
            .O(N__29747),
            .I(bfn_11_17_0_));
    InMux I__5387 (
            .O(N__29744),
            .I(\current_shift_inst.un4_control_input_cry_25 ));
    InMux I__5386 (
            .O(N__29741),
            .I(\current_shift_inst.un4_control_input_cry_26 ));
    InMux I__5385 (
            .O(N__29738),
            .I(N__29733));
    InMux I__5384 (
            .O(N__29737),
            .I(N__29728));
    InMux I__5383 (
            .O(N__29736),
            .I(N__29728));
    LocalMux I__5382 (
            .O(N__29733),
            .I(N__29725));
    LocalMux I__5381 (
            .O(N__29728),
            .I(N__29722));
    Span4Mux_v I__5380 (
            .O(N__29725),
            .I(N__29718));
    Span4Mux_h I__5379 (
            .O(N__29722),
            .I(N__29715));
    InMux I__5378 (
            .O(N__29721),
            .I(N__29712));
    Odrv4 I__5377 (
            .O(N__29718),
            .I(\current_shift_inst.un4_control_input_cry_10_c_RNIJLTGZ0 ));
    Odrv4 I__5376 (
            .O(N__29715),
            .I(\current_shift_inst.un4_control_input_cry_10_c_RNIJLTGZ0 ));
    LocalMux I__5375 (
            .O(N__29712),
            .I(\current_shift_inst.un4_control_input_cry_10_c_RNIJLTGZ0 ));
    InMux I__5374 (
            .O(N__29705),
            .I(\current_shift_inst.un4_control_input_cry_10 ));
    InMux I__5373 (
            .O(N__29702),
            .I(\current_shift_inst.un4_control_input_cry_11 ));
    InMux I__5372 (
            .O(N__29699),
            .I(\current_shift_inst.un4_control_input_cry_12 ));
    InMux I__5371 (
            .O(N__29696),
            .I(\current_shift_inst.un4_control_input_cry_13 ));
    InMux I__5370 (
            .O(N__29693),
            .I(\current_shift_inst.un4_control_input_cry_14 ));
    InMux I__5369 (
            .O(N__29690),
            .I(\current_shift_inst.un4_control_input_cry_15 ));
    InMux I__5368 (
            .O(N__29687),
            .I(bfn_11_16_0_));
    CascadeMux I__5367 (
            .O(N__29684),
            .I(N__29681));
    InMux I__5366 (
            .O(N__29681),
            .I(N__29676));
    InMux I__5365 (
            .O(N__29680),
            .I(N__29671));
    InMux I__5364 (
            .O(N__29679),
            .I(N__29671));
    LocalMux I__5363 (
            .O(N__29676),
            .I(N__29667));
    LocalMux I__5362 (
            .O(N__29671),
            .I(N__29664));
    CascadeMux I__5361 (
            .O(N__29670),
            .I(N__29661));
    Span4Mux_h I__5360 (
            .O(N__29667),
            .I(N__29656));
    Span4Mux_v I__5359 (
            .O(N__29664),
            .I(N__29656));
    InMux I__5358 (
            .O(N__29661),
            .I(N__29653));
    Odrv4 I__5357 (
            .O(N__29656),
            .I(\current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0 ));
    LocalMux I__5356 (
            .O(N__29653),
            .I(\current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0 ));
    InMux I__5355 (
            .O(N__29648),
            .I(\current_shift_inst.un4_control_input_cry_17 ));
    InMux I__5354 (
            .O(N__29645),
            .I(N__29642));
    LocalMux I__5353 (
            .O(N__29642),
            .I(N__29637));
    InMux I__5352 (
            .O(N__29641),
            .I(N__29632));
    InMux I__5351 (
            .O(N__29640),
            .I(N__29632));
    Span4Mux_v I__5350 (
            .O(N__29637),
            .I(N__29628));
    LocalMux I__5349 (
            .O(N__29632),
            .I(N__29625));
    InMux I__5348 (
            .O(N__29631),
            .I(N__29622));
    Odrv4 I__5347 (
            .O(N__29628),
            .I(\current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0 ));
    Odrv4 I__5346 (
            .O(N__29625),
            .I(\current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0 ));
    LocalMux I__5345 (
            .O(N__29622),
            .I(\current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0 ));
    CascadeMux I__5344 (
            .O(N__29615),
            .I(N__29611));
    InMux I__5343 (
            .O(N__29614),
            .I(N__29608));
    InMux I__5342 (
            .O(N__29611),
            .I(N__29605));
    LocalMux I__5341 (
            .O(N__29608),
            .I(N__29599));
    LocalMux I__5340 (
            .O(N__29605),
            .I(N__29599));
    CascadeMux I__5339 (
            .O(N__29604),
            .I(N__29596));
    Span4Mux_v I__5338 (
            .O(N__29599),
            .I(N__29593));
    InMux I__5337 (
            .O(N__29596),
            .I(N__29590));
    Odrv4 I__5336 (
            .O(N__29593),
            .I(\current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0 ));
    LocalMux I__5335 (
            .O(N__29590),
            .I(\current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0 ));
    InMux I__5334 (
            .O(N__29585),
            .I(\current_shift_inst.un4_control_input_cry_1 ));
    InMux I__5333 (
            .O(N__29582),
            .I(N__29578));
    InMux I__5332 (
            .O(N__29581),
            .I(N__29575));
    LocalMux I__5331 (
            .O(N__29578),
            .I(N__29570));
    LocalMux I__5330 (
            .O(N__29575),
            .I(N__29570));
    Span4Mux_h I__5329 (
            .O(N__29570),
            .I(N__29566));
    InMux I__5328 (
            .O(N__29569),
            .I(N__29563));
    Odrv4 I__5327 (
            .O(N__29566),
            .I(\current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0 ));
    LocalMux I__5326 (
            .O(N__29563),
            .I(\current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0 ));
    InMux I__5325 (
            .O(N__29558),
            .I(\current_shift_inst.un4_control_input_cry_2 ));
    InMux I__5324 (
            .O(N__29555),
            .I(N__29552));
    LocalMux I__5323 (
            .O(N__29552),
            .I(N__29549));
    Span4Mux_h I__5322 (
            .O(N__29549),
            .I(N__29545));
    InMux I__5321 (
            .O(N__29548),
            .I(N__29542));
    Odrv4 I__5320 (
            .O(N__29545),
            .I(\current_shift_inst.un4_control_input_cry_3_c_RNINL4GZ0 ));
    LocalMux I__5319 (
            .O(N__29542),
            .I(\current_shift_inst.un4_control_input_cry_3_c_RNINL4GZ0 ));
    InMux I__5318 (
            .O(N__29537),
            .I(\current_shift_inst.un4_control_input_cry_3 ));
    CascadeMux I__5317 (
            .O(N__29534),
            .I(N__29531));
    InMux I__5316 (
            .O(N__29531),
            .I(N__29526));
    InMux I__5315 (
            .O(N__29530),
            .I(N__29523));
    InMux I__5314 (
            .O(N__29529),
            .I(N__29520));
    LocalMux I__5313 (
            .O(N__29526),
            .I(N__29514));
    LocalMux I__5312 (
            .O(N__29523),
            .I(N__29514));
    LocalMux I__5311 (
            .O(N__29520),
            .I(N__29511));
    CascadeMux I__5310 (
            .O(N__29519),
            .I(N__29508));
    Span4Mux_h I__5309 (
            .O(N__29514),
            .I(N__29505));
    Span4Mux_h I__5308 (
            .O(N__29511),
            .I(N__29502));
    InMux I__5307 (
            .O(N__29508),
            .I(N__29499));
    Odrv4 I__5306 (
            .O(N__29505),
            .I(\current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0 ));
    Odrv4 I__5305 (
            .O(N__29502),
            .I(\current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0 ));
    LocalMux I__5304 (
            .O(N__29499),
            .I(\current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0 ));
    InMux I__5303 (
            .O(N__29492),
            .I(\current_shift_inst.un4_control_input_cry_4 ));
    InMux I__5302 (
            .O(N__29489),
            .I(N__29484));
    InMux I__5301 (
            .O(N__29488),
            .I(N__29479));
    InMux I__5300 (
            .O(N__29487),
            .I(N__29479));
    LocalMux I__5299 (
            .O(N__29484),
            .I(N__29476));
    LocalMux I__5298 (
            .O(N__29479),
            .I(N__29473));
    Span4Mux_v I__5297 (
            .O(N__29476),
            .I(N__29469));
    Span4Mux_h I__5296 (
            .O(N__29473),
            .I(N__29466));
    InMux I__5295 (
            .O(N__29472),
            .I(N__29463));
    Odrv4 I__5294 (
            .O(N__29469),
            .I(\current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0 ));
    Odrv4 I__5293 (
            .O(N__29466),
            .I(\current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0 ));
    LocalMux I__5292 (
            .O(N__29463),
            .I(\current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0 ));
    InMux I__5291 (
            .O(N__29456),
            .I(\current_shift_inst.un4_control_input_cry_5 ));
    InMux I__5290 (
            .O(N__29453),
            .I(N__29448));
    InMux I__5289 (
            .O(N__29452),
            .I(N__29443));
    InMux I__5288 (
            .O(N__29451),
            .I(N__29443));
    LocalMux I__5287 (
            .O(N__29448),
            .I(N__29439));
    LocalMux I__5286 (
            .O(N__29443),
            .I(N__29436));
    CascadeMux I__5285 (
            .O(N__29442),
            .I(N__29433));
    Span4Mux_h I__5284 (
            .O(N__29439),
            .I(N__29430));
    Span4Mux_v I__5283 (
            .O(N__29436),
            .I(N__29427));
    InMux I__5282 (
            .O(N__29433),
            .I(N__29424));
    Odrv4 I__5281 (
            .O(N__29430),
            .I(\current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0 ));
    Odrv4 I__5280 (
            .O(N__29427),
            .I(\current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0 ));
    LocalMux I__5279 (
            .O(N__29424),
            .I(\current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0 ));
    InMux I__5278 (
            .O(N__29417),
            .I(\current_shift_inst.un4_control_input_cry_6 ));
    CascadeMux I__5277 (
            .O(N__29414),
            .I(N__29411));
    InMux I__5276 (
            .O(N__29411),
            .I(N__29408));
    LocalMux I__5275 (
            .O(N__29408),
            .I(N__29404));
    CascadeMux I__5274 (
            .O(N__29407),
            .I(N__29400));
    Span4Mux_h I__5273 (
            .O(N__29404),
            .I(N__29397));
    InMux I__5272 (
            .O(N__29403),
            .I(N__29392));
    InMux I__5271 (
            .O(N__29400),
            .I(N__29392));
    Sp12to4 I__5270 (
            .O(N__29397),
            .I(N__29388));
    LocalMux I__5269 (
            .O(N__29392),
            .I(N__29385));
    CascadeMux I__5268 (
            .O(N__29391),
            .I(N__29382));
    Span12Mux_v I__5267 (
            .O(N__29388),
            .I(N__29379));
    Span4Mux_v I__5266 (
            .O(N__29385),
            .I(N__29376));
    InMux I__5265 (
            .O(N__29382),
            .I(N__29373));
    Odrv12 I__5264 (
            .O(N__29379),
            .I(\current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0 ));
    Odrv4 I__5263 (
            .O(N__29376),
            .I(\current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0 ));
    LocalMux I__5262 (
            .O(N__29373),
            .I(\current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0 ));
    InMux I__5261 (
            .O(N__29366),
            .I(\current_shift_inst.un4_control_input_cry_7 ));
    InMux I__5260 (
            .O(N__29363),
            .I(bfn_11_15_0_));
    InMux I__5259 (
            .O(N__29360),
            .I(\current_shift_inst.un4_control_input_cry_9 ));
    CascadeMux I__5258 (
            .O(N__29357),
            .I(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6_cascade_ ));
    CascadeMux I__5257 (
            .O(N__29354),
            .I(N__29351));
    InMux I__5256 (
            .O(N__29351),
            .I(N__29348));
    LocalMux I__5255 (
            .O(N__29348),
            .I(N__29345));
    Odrv4 I__5254 (
            .O(N__29345),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ));
    CascadeMux I__5253 (
            .O(N__29342),
            .I(N__29339));
    InMux I__5252 (
            .O(N__29339),
            .I(N__29336));
    LocalMux I__5251 (
            .O(N__29336),
            .I(N__29333));
    Span4Mux_h I__5250 (
            .O(N__29333),
            .I(N__29330));
    Odrv4 I__5249 (
            .O(N__29330),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ));
    CascadeMux I__5248 (
            .O(N__29327),
            .I(N__29322));
    InMux I__5247 (
            .O(N__29326),
            .I(N__29319));
    InMux I__5246 (
            .O(N__29325),
            .I(N__29316));
    InMux I__5245 (
            .O(N__29322),
            .I(N__29313));
    LocalMux I__5244 (
            .O(N__29319),
            .I(\current_shift_inst.elapsed_time_ns_1_fast_31 ));
    LocalMux I__5243 (
            .O(N__29316),
            .I(\current_shift_inst.elapsed_time_ns_1_fast_31 ));
    LocalMux I__5242 (
            .O(N__29313),
            .I(\current_shift_inst.elapsed_time_ns_1_fast_31 ));
    CascadeMux I__5241 (
            .O(N__29306),
            .I(N__29303));
    InMux I__5240 (
            .O(N__29303),
            .I(N__29300));
    LocalMux I__5239 (
            .O(N__29300),
            .I(N__29297));
    Span4Mux_v I__5238 (
            .O(N__29297),
            .I(N__29294));
    Span4Mux_h I__5237 (
            .O(N__29294),
            .I(N__29290));
    InMux I__5236 (
            .O(N__29293),
            .I(N__29287));
    Odrv4 I__5235 (
            .O(N__29290),
            .I(\current_shift_inst.un38_control_input_0 ));
    LocalMux I__5234 (
            .O(N__29287),
            .I(\current_shift_inst.un38_control_input_0 ));
    InMux I__5233 (
            .O(N__29282),
            .I(N__29279));
    LocalMux I__5232 (
            .O(N__29279),
            .I(N__29275));
    InMux I__5231 (
            .O(N__29278),
            .I(N__29272));
    Span4Mux_h I__5230 (
            .O(N__29275),
            .I(N__29269));
    LocalMux I__5229 (
            .O(N__29272),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    Odrv4 I__5228 (
            .O(N__29269),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__5227 (
            .O(N__29264),
            .I(N__29261));
    LocalMux I__5226 (
            .O(N__29261),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13 ));
    InMux I__5225 (
            .O(N__29258),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ));
    InMux I__5224 (
            .O(N__29255),
            .I(N__29251));
    InMux I__5223 (
            .O(N__29254),
            .I(N__29248));
    LocalMux I__5222 (
            .O(N__29251),
            .I(N__29245));
    LocalMux I__5221 (
            .O(N__29248),
            .I(N__29242));
    Odrv12 I__5220 (
            .O(N__29245),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    Odrv4 I__5219 (
            .O(N__29242),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    InMux I__5218 (
            .O(N__29237),
            .I(N__29234));
    LocalMux I__5217 (
            .O(N__29234),
            .I(N__29231));
    Odrv4 I__5216 (
            .O(N__29231),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14 ));
    InMux I__5215 (
            .O(N__29228),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ));
    InMux I__5214 (
            .O(N__29225),
            .I(N__29222));
    LocalMux I__5213 (
            .O(N__29222),
            .I(N__29218));
    InMux I__5212 (
            .O(N__29221),
            .I(N__29215));
    Span4Mux_v I__5211 (
            .O(N__29218),
            .I(N__29212));
    LocalMux I__5210 (
            .O(N__29215),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    Odrv4 I__5209 (
            .O(N__29212),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__5208 (
            .O(N__29207),
            .I(N__29204));
    LocalMux I__5207 (
            .O(N__29204),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15 ));
    InMux I__5206 (
            .O(N__29201),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ));
    InMux I__5205 (
            .O(N__29198),
            .I(N__29195));
    LocalMux I__5204 (
            .O(N__29195),
            .I(N__29191));
    InMux I__5203 (
            .O(N__29194),
            .I(N__29188));
    Span4Mux_h I__5202 (
            .O(N__29191),
            .I(N__29185));
    LocalMux I__5201 (
            .O(N__29188),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    Odrv4 I__5200 (
            .O(N__29185),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    InMux I__5199 (
            .O(N__29180),
            .I(N__29177));
    LocalMux I__5198 (
            .O(N__29177),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16 ));
    InMux I__5197 (
            .O(N__29174),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ));
    InMux I__5196 (
            .O(N__29171),
            .I(N__29168));
    LocalMux I__5195 (
            .O(N__29168),
            .I(N__29164));
    InMux I__5194 (
            .O(N__29167),
            .I(N__29161));
    Span4Mux_h I__5193 (
            .O(N__29164),
            .I(N__29158));
    LocalMux I__5192 (
            .O(N__29161),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    Odrv4 I__5191 (
            .O(N__29158),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    InMux I__5190 (
            .O(N__29153),
            .I(N__29150));
    LocalMux I__5189 (
            .O(N__29150),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17 ));
    InMux I__5188 (
            .O(N__29147),
            .I(bfn_11_10_0_));
    InMux I__5187 (
            .O(N__29144),
            .I(N__29141));
    LocalMux I__5186 (
            .O(N__29141),
            .I(N__29137));
    InMux I__5185 (
            .O(N__29140),
            .I(N__29134));
    Span4Mux_v I__5184 (
            .O(N__29137),
            .I(N__29131));
    LocalMux I__5183 (
            .O(N__29134),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    Odrv4 I__5182 (
            .O(N__29131),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__5181 (
            .O(N__29126),
            .I(N__29123));
    LocalMux I__5180 (
            .O(N__29123),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18 ));
    InMux I__5179 (
            .O(N__29120),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ));
    InMux I__5178 (
            .O(N__29117),
            .I(N__29114));
    LocalMux I__5177 (
            .O(N__29114),
            .I(N__29110));
    InMux I__5176 (
            .O(N__29113),
            .I(N__29107));
    Span4Mux_h I__5175 (
            .O(N__29110),
            .I(N__29104));
    LocalMux I__5174 (
            .O(N__29107),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    Odrv4 I__5173 (
            .O(N__29104),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__5172 (
            .O(N__29099),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17 ));
    InMux I__5171 (
            .O(N__29096),
            .I(N__29093));
    LocalMux I__5170 (
            .O(N__29093),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19 ));
    InMux I__5169 (
            .O(N__29090),
            .I(N__29087));
    LocalMux I__5168 (
            .O(N__29087),
            .I(N__29084));
    Odrv12 I__5167 (
            .O(N__29084),
            .I(il_min_comp1_D1));
    InMux I__5166 (
            .O(N__29081),
            .I(N__29078));
    LocalMux I__5165 (
            .O(N__29078),
            .I(N__29075));
    Span4Mux_v I__5164 (
            .O(N__29075),
            .I(N__29071));
    InMux I__5163 (
            .O(N__29074),
            .I(N__29068));
    Odrv4 I__5162 (
            .O(N__29071),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    LocalMux I__5161 (
            .O(N__29068),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    InMux I__5160 (
            .O(N__29063),
            .I(N__29060));
    LocalMux I__5159 (
            .O(N__29060),
            .I(N__29057));
    Span4Mux_h I__5158 (
            .O(N__29057),
            .I(N__29054));
    Odrv4 I__5157 (
            .O(N__29054),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5 ));
    InMux I__5156 (
            .O(N__29051),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ));
    InMux I__5155 (
            .O(N__29048),
            .I(N__29045));
    LocalMux I__5154 (
            .O(N__29045),
            .I(N__29042));
    Span4Mux_h I__5153 (
            .O(N__29042),
            .I(N__29038));
    InMux I__5152 (
            .O(N__29041),
            .I(N__29035));
    Odrv4 I__5151 (
            .O(N__29038),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    LocalMux I__5150 (
            .O(N__29035),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    InMux I__5149 (
            .O(N__29030),
            .I(N__29027));
    LocalMux I__5148 (
            .O(N__29027),
            .I(N__29024));
    Span4Mux_h I__5147 (
            .O(N__29024),
            .I(N__29021));
    Odrv4 I__5146 (
            .O(N__29021),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6 ));
    InMux I__5145 (
            .O(N__29018),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ));
    InMux I__5144 (
            .O(N__29015),
            .I(N__29012));
    LocalMux I__5143 (
            .O(N__29012),
            .I(N__29009));
    Span4Mux_h I__5142 (
            .O(N__29009),
            .I(N__29005));
    InMux I__5141 (
            .O(N__29008),
            .I(N__29002));
    Odrv4 I__5140 (
            .O(N__29005),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    LocalMux I__5139 (
            .O(N__29002),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    InMux I__5138 (
            .O(N__28997),
            .I(N__28994));
    LocalMux I__5137 (
            .O(N__28994),
            .I(N__28991));
    Span4Mux_h I__5136 (
            .O(N__28991),
            .I(N__28988));
    Odrv4 I__5135 (
            .O(N__28988),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7 ));
    InMux I__5134 (
            .O(N__28985),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ));
    InMux I__5133 (
            .O(N__28982),
            .I(N__28979));
    LocalMux I__5132 (
            .O(N__28979),
            .I(N__28975));
    InMux I__5131 (
            .O(N__28978),
            .I(N__28972));
    Span4Mux_h I__5130 (
            .O(N__28975),
            .I(N__28967));
    LocalMux I__5129 (
            .O(N__28972),
            .I(N__28967));
    Odrv4 I__5128 (
            .O(N__28967),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    InMux I__5127 (
            .O(N__28964),
            .I(N__28961));
    LocalMux I__5126 (
            .O(N__28961),
            .I(N__28958));
    Span4Mux_h I__5125 (
            .O(N__28958),
            .I(N__28955));
    Odrv4 I__5124 (
            .O(N__28955),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8 ));
    InMux I__5123 (
            .O(N__28952),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ));
    InMux I__5122 (
            .O(N__28949),
            .I(bfn_11_9_0_));
    InMux I__5121 (
            .O(N__28946),
            .I(N__28942));
    InMux I__5120 (
            .O(N__28945),
            .I(N__28939));
    LocalMux I__5119 (
            .O(N__28942),
            .I(N__28936));
    LocalMux I__5118 (
            .O(N__28939),
            .I(N__28933));
    Odrv4 I__5117 (
            .O(N__28936),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    Odrv4 I__5116 (
            .O(N__28933),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    InMux I__5115 (
            .O(N__28928),
            .I(N__28925));
    LocalMux I__5114 (
            .O(N__28925),
            .I(N__28922));
    Odrv12 I__5113 (
            .O(N__28922),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10 ));
    InMux I__5112 (
            .O(N__28919),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ));
    InMux I__5111 (
            .O(N__28916),
            .I(N__28912));
    CascadeMux I__5110 (
            .O(N__28915),
            .I(N__28909));
    LocalMux I__5109 (
            .O(N__28912),
            .I(N__28906));
    InMux I__5108 (
            .O(N__28909),
            .I(N__28903));
    Span4Mux_v I__5107 (
            .O(N__28906),
            .I(N__28900));
    LocalMux I__5106 (
            .O(N__28903),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    Odrv4 I__5105 (
            .O(N__28900),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    InMux I__5104 (
            .O(N__28895),
            .I(N__28892));
    LocalMux I__5103 (
            .O(N__28892),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11 ));
    InMux I__5102 (
            .O(N__28889),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ));
    InMux I__5101 (
            .O(N__28886),
            .I(N__28882));
    CascadeMux I__5100 (
            .O(N__28885),
            .I(N__28879));
    LocalMux I__5099 (
            .O(N__28882),
            .I(N__28876));
    InMux I__5098 (
            .O(N__28879),
            .I(N__28873));
    Span4Mux_h I__5097 (
            .O(N__28876),
            .I(N__28870));
    LocalMux I__5096 (
            .O(N__28873),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    Odrv4 I__5095 (
            .O(N__28870),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__5094 (
            .O(N__28865),
            .I(N__28862));
    LocalMux I__5093 (
            .O(N__28862),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12 ));
    InMux I__5092 (
            .O(N__28859),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ));
    InMux I__5091 (
            .O(N__28856),
            .I(N__28824));
    InMux I__5090 (
            .O(N__28855),
            .I(N__28810));
    InMux I__5089 (
            .O(N__28854),
            .I(N__28810));
    InMux I__5088 (
            .O(N__28853),
            .I(N__28810));
    InMux I__5087 (
            .O(N__28852),
            .I(N__28801));
    InMux I__5086 (
            .O(N__28851),
            .I(N__28801));
    InMux I__5085 (
            .O(N__28850),
            .I(N__28801));
    InMux I__5084 (
            .O(N__28849),
            .I(N__28801));
    CascadeMux I__5083 (
            .O(N__28848),
            .I(N__28797));
    CascadeMux I__5082 (
            .O(N__28847),
            .I(N__28793));
    CascadeMux I__5081 (
            .O(N__28846),
            .I(N__28789));
    CascadeMux I__5080 (
            .O(N__28845),
            .I(N__28786));
    CascadeMux I__5079 (
            .O(N__28844),
            .I(N__28783));
    CascadeMux I__5078 (
            .O(N__28843),
            .I(N__28780));
    CascadeMux I__5077 (
            .O(N__28842),
            .I(N__28777));
    CascadeMux I__5076 (
            .O(N__28841),
            .I(N__28774));
    CascadeMux I__5075 (
            .O(N__28840),
            .I(N__28771));
    CascadeMux I__5074 (
            .O(N__28839),
            .I(N__28768));
    CascadeMux I__5073 (
            .O(N__28838),
            .I(N__28765));
    CascadeMux I__5072 (
            .O(N__28837),
            .I(N__28762));
    CascadeMux I__5071 (
            .O(N__28836),
            .I(N__28759));
    CascadeMux I__5070 (
            .O(N__28835),
            .I(N__28756));
    CascadeMux I__5069 (
            .O(N__28834),
            .I(N__28753));
    CascadeMux I__5068 (
            .O(N__28833),
            .I(N__28750));
    CascadeMux I__5067 (
            .O(N__28832),
            .I(N__28747));
    CascadeMux I__5066 (
            .O(N__28831),
            .I(N__28744));
    CascadeMux I__5065 (
            .O(N__28830),
            .I(N__28741));
    CascadeMux I__5064 (
            .O(N__28829),
            .I(N__28738));
    CascadeMux I__5063 (
            .O(N__28828),
            .I(N__28735));
    CascadeMux I__5062 (
            .O(N__28827),
            .I(N__28732));
    LocalMux I__5061 (
            .O(N__28824),
            .I(N__28728));
    InMux I__5060 (
            .O(N__28823),
            .I(N__28721));
    InMux I__5059 (
            .O(N__28822),
            .I(N__28721));
    InMux I__5058 (
            .O(N__28821),
            .I(N__28721));
    InMux I__5057 (
            .O(N__28820),
            .I(N__28712));
    InMux I__5056 (
            .O(N__28819),
            .I(N__28712));
    InMux I__5055 (
            .O(N__28818),
            .I(N__28712));
    InMux I__5054 (
            .O(N__28817),
            .I(N__28712));
    LocalMux I__5053 (
            .O(N__28810),
            .I(N__28707));
    LocalMux I__5052 (
            .O(N__28801),
            .I(N__28707));
    InMux I__5051 (
            .O(N__28800),
            .I(N__28700));
    InMux I__5050 (
            .O(N__28797),
            .I(N__28700));
    InMux I__5049 (
            .O(N__28796),
            .I(N__28700));
    InMux I__5048 (
            .O(N__28793),
            .I(N__28682));
    InMux I__5047 (
            .O(N__28792),
            .I(N__28682));
    InMux I__5046 (
            .O(N__28789),
            .I(N__28682));
    InMux I__5045 (
            .O(N__28786),
            .I(N__28682));
    InMux I__5044 (
            .O(N__28783),
            .I(N__28682));
    InMux I__5043 (
            .O(N__28780),
            .I(N__28675));
    InMux I__5042 (
            .O(N__28777),
            .I(N__28675));
    InMux I__5041 (
            .O(N__28774),
            .I(N__28675));
    InMux I__5040 (
            .O(N__28771),
            .I(N__28666));
    InMux I__5039 (
            .O(N__28768),
            .I(N__28666));
    InMux I__5038 (
            .O(N__28765),
            .I(N__28666));
    InMux I__5037 (
            .O(N__28762),
            .I(N__28666));
    InMux I__5036 (
            .O(N__28759),
            .I(N__28657));
    InMux I__5035 (
            .O(N__28756),
            .I(N__28657));
    InMux I__5034 (
            .O(N__28753),
            .I(N__28657));
    InMux I__5033 (
            .O(N__28750),
            .I(N__28657));
    InMux I__5032 (
            .O(N__28747),
            .I(N__28649));
    InMux I__5031 (
            .O(N__28744),
            .I(N__28649));
    InMux I__5030 (
            .O(N__28741),
            .I(N__28649));
    InMux I__5029 (
            .O(N__28738),
            .I(N__28642));
    InMux I__5028 (
            .O(N__28735),
            .I(N__28642));
    InMux I__5027 (
            .O(N__28732),
            .I(N__28642));
    InMux I__5026 (
            .O(N__28731),
            .I(N__28639));
    Span4Mux_v I__5025 (
            .O(N__28728),
            .I(N__28632));
    LocalMux I__5024 (
            .O(N__28721),
            .I(N__28632));
    LocalMux I__5023 (
            .O(N__28712),
            .I(N__28632));
    Span4Mux_s2_h I__5022 (
            .O(N__28707),
            .I(N__28627));
    LocalMux I__5021 (
            .O(N__28700),
            .I(N__28627));
    CascadeMux I__5020 (
            .O(N__28699),
            .I(N__28624));
    CascadeMux I__5019 (
            .O(N__28698),
            .I(N__28621));
    CascadeMux I__5018 (
            .O(N__28697),
            .I(N__28618));
    CascadeMux I__5017 (
            .O(N__28696),
            .I(N__28615));
    CascadeMux I__5016 (
            .O(N__28695),
            .I(N__28612));
    CascadeMux I__5015 (
            .O(N__28694),
            .I(N__28609));
    CascadeMux I__5014 (
            .O(N__28693),
            .I(N__28606));
    LocalMux I__5013 (
            .O(N__28682),
            .I(N__28603));
    LocalMux I__5012 (
            .O(N__28675),
            .I(N__28600));
    LocalMux I__5011 (
            .O(N__28666),
            .I(N__28595));
    LocalMux I__5010 (
            .O(N__28657),
            .I(N__28595));
    InMux I__5009 (
            .O(N__28656),
            .I(N__28592));
    LocalMux I__5008 (
            .O(N__28649),
            .I(N__28587));
    LocalMux I__5007 (
            .O(N__28642),
            .I(N__28587));
    LocalMux I__5006 (
            .O(N__28639),
            .I(N__28582));
    Span4Mux_v I__5005 (
            .O(N__28632),
            .I(N__28582));
    Sp12to4 I__5004 (
            .O(N__28627),
            .I(N__28579));
    InMux I__5003 (
            .O(N__28624),
            .I(N__28572));
    InMux I__5002 (
            .O(N__28621),
            .I(N__28572));
    InMux I__5001 (
            .O(N__28618),
            .I(N__28572));
    InMux I__5000 (
            .O(N__28615),
            .I(N__28563));
    InMux I__4999 (
            .O(N__28612),
            .I(N__28563));
    InMux I__4998 (
            .O(N__28609),
            .I(N__28563));
    InMux I__4997 (
            .O(N__28606),
            .I(N__28563));
    Span4Mux_v I__4996 (
            .O(N__28603),
            .I(N__28558));
    Span4Mux_v I__4995 (
            .O(N__28600),
            .I(N__28558));
    Span4Mux_v I__4994 (
            .O(N__28595),
            .I(N__28555));
    LocalMux I__4993 (
            .O(N__28592),
            .I(N__28552));
    Span4Mux_h I__4992 (
            .O(N__28587),
            .I(N__28549));
    Span4Mux_h I__4991 (
            .O(N__28582),
            .I(N__28544));
    Span12Mux_v I__4990 (
            .O(N__28579),
            .I(N__28537));
    LocalMux I__4989 (
            .O(N__28572),
            .I(N__28537));
    LocalMux I__4988 (
            .O(N__28563),
            .I(N__28537));
    Span4Mux_v I__4987 (
            .O(N__28558),
            .I(N__28532));
    Span4Mux_v I__4986 (
            .O(N__28555),
            .I(N__28532));
    Span4Mux_v I__4985 (
            .O(N__28552),
            .I(N__28529));
    Span4Mux_v I__4984 (
            .O(N__28549),
            .I(N__28525));
    InMux I__4983 (
            .O(N__28548),
            .I(N__28522));
    InMux I__4982 (
            .O(N__28547),
            .I(N__28519));
    Sp12to4 I__4981 (
            .O(N__28544),
            .I(N__28516));
    Span12Mux_h I__4980 (
            .O(N__28537),
            .I(N__28513));
    Span4Mux_v I__4979 (
            .O(N__28532),
            .I(N__28510));
    Sp12to4 I__4978 (
            .O(N__28529),
            .I(N__28507));
    InMux I__4977 (
            .O(N__28528),
            .I(N__28504));
    Span4Mux_v I__4976 (
            .O(N__28525),
            .I(N__28501));
    LocalMux I__4975 (
            .O(N__28522),
            .I(N__28496));
    LocalMux I__4974 (
            .O(N__28519),
            .I(N__28496));
    Span12Mux_v I__4973 (
            .O(N__28516),
            .I(N__28493));
    Span12Mux_v I__4972 (
            .O(N__28513),
            .I(N__28486));
    Sp12to4 I__4971 (
            .O(N__28510),
            .I(N__28486));
    Span12Mux_s11_h I__4970 (
            .O(N__28507),
            .I(N__28486));
    LocalMux I__4969 (
            .O(N__28504),
            .I(N__28483));
    Span4Mux_h I__4968 (
            .O(N__28501),
            .I(N__28478));
    Span4Mux_h I__4967 (
            .O(N__28496),
            .I(N__28478));
    Odrv12 I__4966 (
            .O(N__28493),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__4965 (
            .O(N__28486),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__4964 (
            .O(N__28483),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__4963 (
            .O(N__28478),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__4962 (
            .O(N__28469),
            .I(N__28466));
    InMux I__4961 (
            .O(N__28466),
            .I(N__28463));
    LocalMux I__4960 (
            .O(N__28463),
            .I(N__28460));
    Span4Mux_h I__4959 (
            .O(N__28460),
            .I(N__28457));
    Odrv4 I__4958 (
            .O(N__28457),
            .I(\current_shift_inst.z_5_30 ));
    InMux I__4957 (
            .O(N__28454),
            .I(\current_shift_inst.z_5_cry_29 ));
    InMux I__4956 (
            .O(N__28451),
            .I(\current_shift_inst.z_5_cry_30 ));
    InMux I__4955 (
            .O(N__28448),
            .I(N__28445));
    LocalMux I__4954 (
            .O(N__28445),
            .I(N__28442));
    Span4Mux_v I__4953 (
            .O(N__28442),
            .I(N__28439));
    Odrv4 I__4952 (
            .O(N__28439),
            .I(\current_shift_inst.z_5_cry_30_THRU_CO ));
    IoInMux I__4951 (
            .O(N__28436),
            .I(N__28433));
    LocalMux I__4950 (
            .O(N__28433),
            .I(N__28430));
    IoSpan4Mux I__4949 (
            .O(N__28430),
            .I(N__28427));
    Span4Mux_s2_v I__4948 (
            .O(N__28427),
            .I(N__28424));
    Odrv4 I__4947 (
            .O(N__28424),
            .I(s4_phy_c));
    InMux I__4946 (
            .O(N__28421),
            .I(N__28418));
    LocalMux I__4945 (
            .O(N__28418),
            .I(N__28415));
    Span4Mux_h I__4944 (
            .O(N__28415),
            .I(N__28412));
    Span4Mux_v I__4943 (
            .O(N__28412),
            .I(N__28409));
    Odrv4 I__4942 (
            .O(N__28409),
            .I(il_min_comp1_c));
    InMux I__4941 (
            .O(N__28406),
            .I(N__28403));
    LocalMux I__4940 (
            .O(N__28403),
            .I(N__28400));
    Span4Mux_h I__4939 (
            .O(N__28400),
            .I(N__28397));
    Span4Mux_v I__4938 (
            .O(N__28397),
            .I(N__28394));
    Odrv4 I__4937 (
            .O(N__28394),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0 ));
    CascadeMux I__4936 (
            .O(N__28391),
            .I(N__28388));
    InMux I__4935 (
            .O(N__28388),
            .I(N__28384));
    InMux I__4934 (
            .O(N__28387),
            .I(N__28381));
    LocalMux I__4933 (
            .O(N__28384),
            .I(N__28378));
    LocalMux I__4932 (
            .O(N__28381),
            .I(N__28374));
    Span4Mux_h I__4931 (
            .O(N__28378),
            .I(N__28371));
    InMux I__4930 (
            .O(N__28377),
            .I(N__28368));
    Odrv4 I__4929 (
            .O(N__28374),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__4928 (
            .O(N__28371),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__4927 (
            .O(N__28368),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    InMux I__4926 (
            .O(N__28361),
            .I(N__28358));
    LocalMux I__4925 (
            .O(N__28358),
            .I(N__28355));
    Span4Mux_h I__4924 (
            .O(N__28355),
            .I(N__28351));
    InMux I__4923 (
            .O(N__28354),
            .I(N__28348));
    Odrv4 I__4922 (
            .O(N__28351),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    LocalMux I__4921 (
            .O(N__28348),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    InMux I__4920 (
            .O(N__28343),
            .I(N__28340));
    LocalMux I__4919 (
            .O(N__28340),
            .I(N__28337));
    Span4Mux_h I__4918 (
            .O(N__28337),
            .I(N__28334));
    Odrv4 I__4917 (
            .O(N__28334),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2 ));
    InMux I__4916 (
            .O(N__28331),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ));
    InMux I__4915 (
            .O(N__28328),
            .I(N__28325));
    LocalMux I__4914 (
            .O(N__28325),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0 ));
    CascadeMux I__4913 (
            .O(N__28322),
            .I(N__28319));
    InMux I__4912 (
            .O(N__28319),
            .I(N__28316));
    LocalMux I__4911 (
            .O(N__28316),
            .I(N__28313));
    Span4Mux_h I__4910 (
            .O(N__28313),
            .I(N__28309));
    InMux I__4909 (
            .O(N__28312),
            .I(N__28306));
    Odrv4 I__4908 (
            .O(N__28309),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    LocalMux I__4907 (
            .O(N__28306),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    InMux I__4906 (
            .O(N__28301),
            .I(N__28298));
    LocalMux I__4905 (
            .O(N__28298),
            .I(N__28295));
    Span4Mux_v I__4904 (
            .O(N__28295),
            .I(N__28292));
    Odrv4 I__4903 (
            .O(N__28292),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3 ));
    InMux I__4902 (
            .O(N__28289),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ));
    InMux I__4901 (
            .O(N__28286),
            .I(N__28283));
    LocalMux I__4900 (
            .O(N__28283),
            .I(N__28280));
    Span4Mux_v I__4899 (
            .O(N__28280),
            .I(N__28276));
    InMux I__4898 (
            .O(N__28279),
            .I(N__28273));
    Odrv4 I__4897 (
            .O(N__28276),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    LocalMux I__4896 (
            .O(N__28273),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    InMux I__4895 (
            .O(N__28268),
            .I(N__28265));
    LocalMux I__4894 (
            .O(N__28265),
            .I(N__28262));
    Span4Mux_v I__4893 (
            .O(N__28262),
            .I(N__28259));
    Odrv4 I__4892 (
            .O(N__28259),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4 ));
    InMux I__4891 (
            .O(N__28256),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ));
    InMux I__4890 (
            .O(N__28253),
            .I(\current_shift_inst.z_5_cry_20 ));
    InMux I__4889 (
            .O(N__28250),
            .I(N__28240));
    InMux I__4888 (
            .O(N__28249),
            .I(N__28240));
    InMux I__4887 (
            .O(N__28248),
            .I(N__28240));
    InMux I__4886 (
            .O(N__28247),
            .I(N__28237));
    LocalMux I__4885 (
            .O(N__28240),
            .I(N__28234));
    LocalMux I__4884 (
            .O(N__28237),
            .I(N__28231));
    Odrv4 I__4883 (
            .O(N__28234),
            .I(\current_shift_inst.elapsed_time_ns_phase_22 ));
    Odrv4 I__4882 (
            .O(N__28231),
            .I(\current_shift_inst.elapsed_time_ns_phase_22 ));
    InMux I__4881 (
            .O(N__28226),
            .I(N__28223));
    LocalMux I__4880 (
            .O(N__28223),
            .I(N__28220));
    Span4Mux_h I__4879 (
            .O(N__28220),
            .I(N__28217));
    Odrv4 I__4878 (
            .O(N__28217),
            .I(\current_shift_inst.z_5_22 ));
    InMux I__4877 (
            .O(N__28214),
            .I(\current_shift_inst.z_5_cry_21 ));
    CascadeMux I__4876 (
            .O(N__28211),
            .I(N__28208));
    InMux I__4875 (
            .O(N__28208),
            .I(N__28205));
    LocalMux I__4874 (
            .O(N__28205),
            .I(N__28202));
    Span4Mux_v I__4873 (
            .O(N__28202),
            .I(N__28199));
    Odrv4 I__4872 (
            .O(N__28199),
            .I(\current_shift_inst.z_5_23 ));
    InMux I__4871 (
            .O(N__28196),
            .I(\current_shift_inst.z_5_cry_22 ));
    InMux I__4870 (
            .O(N__28193),
            .I(N__28190));
    LocalMux I__4869 (
            .O(N__28190),
            .I(N__28187));
    Span4Mux_h I__4868 (
            .O(N__28187),
            .I(N__28184));
    Odrv4 I__4867 (
            .O(N__28184),
            .I(\current_shift_inst.z_5_24 ));
    InMux I__4866 (
            .O(N__28181),
            .I(\current_shift_inst.z_5_cry_23 ));
    CascadeMux I__4865 (
            .O(N__28178),
            .I(N__28175));
    InMux I__4864 (
            .O(N__28175),
            .I(N__28172));
    LocalMux I__4863 (
            .O(N__28172),
            .I(N__28169));
    Span4Mux_h I__4862 (
            .O(N__28169),
            .I(N__28166));
    Odrv4 I__4861 (
            .O(N__28166),
            .I(\current_shift_inst.z_5_25 ));
    InMux I__4860 (
            .O(N__28163),
            .I(bfn_10_21_0_));
    InMux I__4859 (
            .O(N__28160),
            .I(N__28157));
    LocalMux I__4858 (
            .O(N__28157),
            .I(N__28154));
    Span4Mux_h I__4857 (
            .O(N__28154),
            .I(N__28151));
    Odrv4 I__4856 (
            .O(N__28151),
            .I(\current_shift_inst.z_5_26 ));
    InMux I__4855 (
            .O(N__28148),
            .I(\current_shift_inst.z_5_cry_25 ));
    CascadeMux I__4854 (
            .O(N__28145),
            .I(N__28141));
    InMux I__4853 (
            .O(N__28144),
            .I(N__28136));
    InMux I__4852 (
            .O(N__28141),
            .I(N__28131));
    InMux I__4851 (
            .O(N__28140),
            .I(N__28131));
    InMux I__4850 (
            .O(N__28139),
            .I(N__28128));
    LocalMux I__4849 (
            .O(N__28136),
            .I(N__28123));
    LocalMux I__4848 (
            .O(N__28131),
            .I(N__28123));
    LocalMux I__4847 (
            .O(N__28128),
            .I(N__28120));
    Span4Mux_v I__4846 (
            .O(N__28123),
            .I(N__28115));
    Span4Mux_h I__4845 (
            .O(N__28120),
            .I(N__28115));
    Odrv4 I__4844 (
            .O(N__28115),
            .I(\current_shift_inst.elapsed_time_ns_phase_27 ));
    InMux I__4843 (
            .O(N__28112),
            .I(N__28109));
    LocalMux I__4842 (
            .O(N__28109),
            .I(N__28106));
    Span4Mux_h I__4841 (
            .O(N__28106),
            .I(N__28103));
    Odrv4 I__4840 (
            .O(N__28103),
            .I(\current_shift_inst.z_5_27 ));
    InMux I__4839 (
            .O(N__28100),
            .I(\current_shift_inst.z_5_cry_26 ));
    InMux I__4838 (
            .O(N__28097),
            .I(N__28094));
    LocalMux I__4837 (
            .O(N__28094),
            .I(N__28091));
    Span4Mux_h I__4836 (
            .O(N__28091),
            .I(N__28088));
    Odrv4 I__4835 (
            .O(N__28088),
            .I(\current_shift_inst.z_5_28 ));
    InMux I__4834 (
            .O(N__28085),
            .I(\current_shift_inst.z_5_cry_27 ));
    CascadeMux I__4833 (
            .O(N__28082),
            .I(N__28079));
    InMux I__4832 (
            .O(N__28079),
            .I(N__28076));
    LocalMux I__4831 (
            .O(N__28076),
            .I(N__28073));
    Span4Mux_h I__4830 (
            .O(N__28073),
            .I(N__28070));
    Odrv4 I__4829 (
            .O(N__28070),
            .I(\current_shift_inst.z_5_29 ));
    InMux I__4828 (
            .O(N__28067),
            .I(\current_shift_inst.z_5_cry_28 ));
    InMux I__4827 (
            .O(N__28064),
            .I(N__28061));
    LocalMux I__4826 (
            .O(N__28061),
            .I(N__28058));
    Span4Mux_h I__4825 (
            .O(N__28058),
            .I(N__28055));
    Odrv4 I__4824 (
            .O(N__28055),
            .I(\current_shift_inst.z_5_13 ));
    InMux I__4823 (
            .O(N__28052),
            .I(\current_shift_inst.z_5_cry_12 ));
    InMux I__4822 (
            .O(N__28049),
            .I(N__28046));
    LocalMux I__4821 (
            .O(N__28046),
            .I(N__28043));
    Span4Mux_h I__4820 (
            .O(N__28043),
            .I(N__28040));
    Odrv4 I__4819 (
            .O(N__28040),
            .I(\current_shift_inst.z_5_14 ));
    InMux I__4818 (
            .O(N__28037),
            .I(\current_shift_inst.z_5_cry_13 ));
    InMux I__4817 (
            .O(N__28034),
            .I(N__28031));
    LocalMux I__4816 (
            .O(N__28031),
            .I(N__28028));
    Span4Mux_v I__4815 (
            .O(N__28028),
            .I(N__28025));
    Odrv4 I__4814 (
            .O(N__28025),
            .I(\current_shift_inst.z_5_15 ));
    InMux I__4813 (
            .O(N__28022),
            .I(\current_shift_inst.z_5_cry_14 ));
    CascadeMux I__4812 (
            .O(N__28019),
            .I(N__28016));
    InMux I__4811 (
            .O(N__28016),
            .I(N__28013));
    LocalMux I__4810 (
            .O(N__28013),
            .I(N__28010));
    Span4Mux_v I__4809 (
            .O(N__28010),
            .I(N__28007));
    Odrv4 I__4808 (
            .O(N__28007),
            .I(\current_shift_inst.z_5_16 ));
    InMux I__4807 (
            .O(N__28004),
            .I(\current_shift_inst.z_5_cry_15 ));
    InMux I__4806 (
            .O(N__28001),
            .I(N__27997));
    CascadeMux I__4805 (
            .O(N__28000),
            .I(N__27994));
    LocalMux I__4804 (
            .O(N__27997),
            .I(N__27989));
    InMux I__4803 (
            .O(N__27994),
            .I(N__27984));
    InMux I__4802 (
            .O(N__27993),
            .I(N__27984));
    InMux I__4801 (
            .O(N__27992),
            .I(N__27981));
    Span12Mux_s9_h I__4800 (
            .O(N__27989),
            .I(N__27976));
    LocalMux I__4799 (
            .O(N__27984),
            .I(N__27976));
    LocalMux I__4798 (
            .O(N__27981),
            .I(N__27973));
    Odrv12 I__4797 (
            .O(N__27976),
            .I(\current_shift_inst.elapsed_time_ns_phase_17 ));
    Odrv4 I__4796 (
            .O(N__27973),
            .I(\current_shift_inst.elapsed_time_ns_phase_17 ));
    InMux I__4795 (
            .O(N__27968),
            .I(N__27965));
    LocalMux I__4794 (
            .O(N__27965),
            .I(N__27962));
    Span4Mux_v I__4793 (
            .O(N__27962),
            .I(N__27959));
    Odrv4 I__4792 (
            .O(N__27959),
            .I(\current_shift_inst.z_5_17 ));
    InMux I__4791 (
            .O(N__27956),
            .I(bfn_10_20_0_));
    CascadeMux I__4790 (
            .O(N__27953),
            .I(N__27950));
    InMux I__4789 (
            .O(N__27950),
            .I(N__27945));
    InMux I__4788 (
            .O(N__27949),
            .I(N__27940));
    InMux I__4787 (
            .O(N__27948),
            .I(N__27940));
    LocalMux I__4786 (
            .O(N__27945),
            .I(N__27934));
    LocalMux I__4785 (
            .O(N__27940),
            .I(N__27934));
    InMux I__4784 (
            .O(N__27939),
            .I(N__27931));
    Span4Mux_v I__4783 (
            .O(N__27934),
            .I(N__27928));
    LocalMux I__4782 (
            .O(N__27931),
            .I(N__27925));
    Odrv4 I__4781 (
            .O(N__27928),
            .I(\current_shift_inst.elapsed_time_ns_phase_18 ));
    Odrv4 I__4780 (
            .O(N__27925),
            .I(\current_shift_inst.elapsed_time_ns_phase_18 ));
    CascadeMux I__4779 (
            .O(N__27920),
            .I(N__27917));
    InMux I__4778 (
            .O(N__27917),
            .I(N__27914));
    LocalMux I__4777 (
            .O(N__27914),
            .I(N__27911));
    Span4Mux_h I__4776 (
            .O(N__27911),
            .I(N__27908));
    Odrv4 I__4775 (
            .O(N__27908),
            .I(\current_shift_inst.z_5_18 ));
    InMux I__4774 (
            .O(N__27905),
            .I(\current_shift_inst.z_5_cry_17 ));
    InMux I__4773 (
            .O(N__27902),
            .I(N__27899));
    LocalMux I__4772 (
            .O(N__27899),
            .I(N__27896));
    Span4Mux_h I__4771 (
            .O(N__27896),
            .I(N__27893));
    Odrv4 I__4770 (
            .O(N__27893),
            .I(\current_shift_inst.z_5_19 ));
    InMux I__4769 (
            .O(N__27890),
            .I(\current_shift_inst.z_5_cry_18 ));
    InMux I__4768 (
            .O(N__27887),
            .I(N__27884));
    LocalMux I__4767 (
            .O(N__27884),
            .I(N__27881));
    Span4Mux_v I__4766 (
            .O(N__27881),
            .I(N__27878));
    Odrv4 I__4765 (
            .O(N__27878),
            .I(\current_shift_inst.z_5_20 ));
    InMux I__4764 (
            .O(N__27875),
            .I(\current_shift_inst.z_5_cry_19 ));
    CascadeMux I__4763 (
            .O(N__27872),
            .I(N__27869));
    InMux I__4762 (
            .O(N__27869),
            .I(N__27866));
    LocalMux I__4761 (
            .O(N__27866),
            .I(N__27863));
    Span4Mux_h I__4760 (
            .O(N__27863),
            .I(N__27860));
    Odrv4 I__4759 (
            .O(N__27860),
            .I(\current_shift_inst.z_5_21 ));
    CascadeMux I__4758 (
            .O(N__27857),
            .I(N__27854));
    InMux I__4757 (
            .O(N__27854),
            .I(N__27849));
    InMux I__4756 (
            .O(N__27853),
            .I(N__27846));
    InMux I__4755 (
            .O(N__27852),
            .I(N__27843));
    LocalMux I__4754 (
            .O(N__27849),
            .I(N__27835));
    LocalMux I__4753 (
            .O(N__27846),
            .I(N__27835));
    LocalMux I__4752 (
            .O(N__27843),
            .I(N__27835));
    InMux I__4751 (
            .O(N__27842),
            .I(N__27832));
    Span4Mux_v I__4750 (
            .O(N__27835),
            .I(N__27829));
    LocalMux I__4749 (
            .O(N__27832),
            .I(N__27826));
    Odrv4 I__4748 (
            .O(N__27829),
            .I(\current_shift_inst.elapsed_time_ns_phase_5 ));
    Odrv4 I__4747 (
            .O(N__27826),
            .I(\current_shift_inst.elapsed_time_ns_phase_5 ));
    CascadeMux I__4746 (
            .O(N__27821),
            .I(N__27818));
    InMux I__4745 (
            .O(N__27818),
            .I(N__27815));
    LocalMux I__4744 (
            .O(N__27815),
            .I(N__27812));
    Span4Mux_h I__4743 (
            .O(N__27812),
            .I(N__27809));
    Odrv4 I__4742 (
            .O(N__27809),
            .I(\current_shift_inst.z_5_5 ));
    InMux I__4741 (
            .O(N__27806),
            .I(\current_shift_inst.z_5_cry_4 ));
    InMux I__4740 (
            .O(N__27803),
            .I(N__27800));
    LocalMux I__4739 (
            .O(N__27800),
            .I(N__27794));
    InMux I__4738 (
            .O(N__27799),
            .I(N__27789));
    InMux I__4737 (
            .O(N__27798),
            .I(N__27789));
    InMux I__4736 (
            .O(N__27797),
            .I(N__27786));
    Span4Mux_v I__4735 (
            .O(N__27794),
            .I(N__27783));
    LocalMux I__4734 (
            .O(N__27789),
            .I(N__27778));
    LocalMux I__4733 (
            .O(N__27786),
            .I(N__27778));
    Odrv4 I__4732 (
            .O(N__27783),
            .I(\current_shift_inst.elapsed_time_ns_phase_6 ));
    Odrv4 I__4731 (
            .O(N__27778),
            .I(\current_shift_inst.elapsed_time_ns_phase_6 ));
    InMux I__4730 (
            .O(N__27773),
            .I(N__27770));
    LocalMux I__4729 (
            .O(N__27770),
            .I(N__27767));
    Span4Mux_h I__4728 (
            .O(N__27767),
            .I(N__27764));
    Odrv4 I__4727 (
            .O(N__27764),
            .I(\current_shift_inst.z_5_6 ));
    InMux I__4726 (
            .O(N__27761),
            .I(\current_shift_inst.z_5_cry_5 ));
    CascadeMux I__4725 (
            .O(N__27758),
            .I(N__27753));
    InMux I__4724 (
            .O(N__27757),
            .I(N__27749));
    InMux I__4723 (
            .O(N__27756),
            .I(N__27746));
    InMux I__4722 (
            .O(N__27753),
            .I(N__27741));
    InMux I__4721 (
            .O(N__27752),
            .I(N__27741));
    LocalMux I__4720 (
            .O(N__27749),
            .I(N__27738));
    LocalMux I__4719 (
            .O(N__27746),
            .I(N__27735));
    LocalMux I__4718 (
            .O(N__27741),
            .I(N__27732));
    Span4Mux_v I__4717 (
            .O(N__27738),
            .I(N__27729));
    Odrv12 I__4716 (
            .O(N__27735),
            .I(\current_shift_inst.elapsed_time_ns_phase_7 ));
    Odrv4 I__4715 (
            .O(N__27732),
            .I(\current_shift_inst.elapsed_time_ns_phase_7 ));
    Odrv4 I__4714 (
            .O(N__27729),
            .I(\current_shift_inst.elapsed_time_ns_phase_7 ));
    InMux I__4713 (
            .O(N__27722),
            .I(N__27719));
    LocalMux I__4712 (
            .O(N__27719),
            .I(N__27716));
    Span4Mux_v I__4711 (
            .O(N__27716),
            .I(N__27713));
    Odrv4 I__4710 (
            .O(N__27713),
            .I(\current_shift_inst.z_5_7 ));
    InMux I__4709 (
            .O(N__27710),
            .I(\current_shift_inst.z_5_cry_6 ));
    InMux I__4708 (
            .O(N__27707),
            .I(N__27704));
    LocalMux I__4707 (
            .O(N__27704),
            .I(N__27701));
    Span4Mux_v I__4706 (
            .O(N__27701),
            .I(N__27698));
    Odrv4 I__4705 (
            .O(N__27698),
            .I(\current_shift_inst.z_5_8 ));
    InMux I__4704 (
            .O(N__27695),
            .I(\current_shift_inst.z_5_cry_7 ));
    InMux I__4703 (
            .O(N__27692),
            .I(N__27689));
    LocalMux I__4702 (
            .O(N__27689),
            .I(N__27686));
    Span4Mux_v I__4701 (
            .O(N__27686),
            .I(N__27683));
    Odrv4 I__4700 (
            .O(N__27683),
            .I(\current_shift_inst.z_5_9 ));
    InMux I__4699 (
            .O(N__27680),
            .I(bfn_10_19_0_));
    InMux I__4698 (
            .O(N__27677),
            .I(N__27669));
    InMux I__4697 (
            .O(N__27676),
            .I(N__27669));
    InMux I__4696 (
            .O(N__27675),
            .I(N__27666));
    InMux I__4695 (
            .O(N__27674),
            .I(N__27663));
    LocalMux I__4694 (
            .O(N__27669),
            .I(N__27660));
    LocalMux I__4693 (
            .O(N__27666),
            .I(N__27655));
    LocalMux I__4692 (
            .O(N__27663),
            .I(N__27655));
    Odrv12 I__4691 (
            .O(N__27660),
            .I(\current_shift_inst.elapsed_time_ns_phase_10 ));
    Odrv4 I__4690 (
            .O(N__27655),
            .I(\current_shift_inst.elapsed_time_ns_phase_10 ));
    CascadeMux I__4689 (
            .O(N__27650),
            .I(N__27647));
    InMux I__4688 (
            .O(N__27647),
            .I(N__27644));
    LocalMux I__4687 (
            .O(N__27644),
            .I(N__27641));
    Span4Mux_h I__4686 (
            .O(N__27641),
            .I(N__27638));
    Odrv4 I__4685 (
            .O(N__27638),
            .I(\current_shift_inst.z_5_10 ));
    InMux I__4684 (
            .O(N__27635),
            .I(\current_shift_inst.z_5_cry_9 ));
    InMux I__4683 (
            .O(N__27632),
            .I(N__27629));
    LocalMux I__4682 (
            .O(N__27629),
            .I(N__27626));
    Span4Mux_h I__4681 (
            .O(N__27626),
            .I(N__27623));
    Odrv4 I__4680 (
            .O(N__27623),
            .I(\current_shift_inst.z_5_11 ));
    InMux I__4679 (
            .O(N__27620),
            .I(\current_shift_inst.z_5_cry_10 ));
    InMux I__4678 (
            .O(N__27617),
            .I(N__27614));
    LocalMux I__4677 (
            .O(N__27614),
            .I(N__27611));
    Span4Mux_h I__4676 (
            .O(N__27611),
            .I(N__27608));
    Odrv4 I__4675 (
            .O(N__27608),
            .I(\current_shift_inst.z_5_12 ));
    InMux I__4674 (
            .O(N__27605),
            .I(\current_shift_inst.z_5_cry_11 ));
    InMux I__4673 (
            .O(N__27602),
            .I(\current_shift_inst.z_cry_30 ));
    InMux I__4672 (
            .O(N__27599),
            .I(N__27592));
    InMux I__4671 (
            .O(N__27598),
            .I(N__27582));
    InMux I__4670 (
            .O(N__27597),
            .I(N__27582));
    InMux I__4669 (
            .O(N__27596),
            .I(N__27582));
    InMux I__4668 (
            .O(N__27595),
            .I(N__27582));
    LocalMux I__4667 (
            .O(N__27592),
            .I(N__27579));
    InMux I__4666 (
            .O(N__27591),
            .I(N__27576));
    LocalMux I__4665 (
            .O(N__27582),
            .I(\current_shift_inst.elapsed_time_ns_phase_1 ));
    Odrv4 I__4664 (
            .O(N__27579),
            .I(\current_shift_inst.elapsed_time_ns_phase_1 ));
    LocalMux I__4663 (
            .O(N__27576),
            .I(\current_shift_inst.elapsed_time_ns_phase_1 ));
    CascadeMux I__4662 (
            .O(N__27569),
            .I(N__27565));
    InMux I__4661 (
            .O(N__27568),
            .I(N__27560));
    InMux I__4660 (
            .O(N__27565),
            .I(N__27555));
    InMux I__4659 (
            .O(N__27564),
            .I(N__27555));
    InMux I__4658 (
            .O(N__27563),
            .I(N__27552));
    LocalMux I__4657 (
            .O(N__27560),
            .I(\current_shift_inst.elapsed_time_ns_phase_2 ));
    LocalMux I__4656 (
            .O(N__27555),
            .I(\current_shift_inst.elapsed_time_ns_phase_2 ));
    LocalMux I__4655 (
            .O(N__27552),
            .I(\current_shift_inst.elapsed_time_ns_phase_2 ));
    CascadeMux I__4654 (
            .O(N__27545),
            .I(N__27542));
    InMux I__4653 (
            .O(N__27542),
            .I(N__27539));
    LocalMux I__4652 (
            .O(N__27539),
            .I(N__27536));
    Span4Mux_h I__4651 (
            .O(N__27536),
            .I(N__27533));
    Odrv4 I__4650 (
            .O(N__27533),
            .I(\current_shift_inst.z_5_2 ));
    InMux I__4649 (
            .O(N__27530),
            .I(\current_shift_inst.z_5_cry_1 ));
    InMux I__4648 (
            .O(N__27527),
            .I(N__27521));
    InMux I__4647 (
            .O(N__27526),
            .I(N__27521));
    LocalMux I__4646 (
            .O(N__27521),
            .I(N__27517));
    InMux I__4645 (
            .O(N__27520),
            .I(N__27514));
    Span4Mux_h I__4644 (
            .O(N__27517),
            .I(N__27509));
    LocalMux I__4643 (
            .O(N__27514),
            .I(N__27509));
    Odrv4 I__4642 (
            .O(N__27509),
            .I(\current_shift_inst.elapsed_time_ns_phase_3 ));
    CascadeMux I__4641 (
            .O(N__27506),
            .I(N__27503));
    InMux I__4640 (
            .O(N__27503),
            .I(N__27500));
    LocalMux I__4639 (
            .O(N__27500),
            .I(N__27497));
    Span4Mux_h I__4638 (
            .O(N__27497),
            .I(N__27494));
    Odrv4 I__4637 (
            .O(N__27494),
            .I(\current_shift_inst.z_5_3 ));
    InMux I__4636 (
            .O(N__27491),
            .I(\current_shift_inst.z_5_cry_2 ));
    InMux I__4635 (
            .O(N__27488),
            .I(N__27480));
    InMux I__4634 (
            .O(N__27487),
            .I(N__27480));
    InMux I__4633 (
            .O(N__27486),
            .I(N__27477));
    InMux I__4632 (
            .O(N__27485),
            .I(N__27474));
    LocalMux I__4631 (
            .O(N__27480),
            .I(N__27469));
    LocalMux I__4630 (
            .O(N__27477),
            .I(N__27469));
    LocalMux I__4629 (
            .O(N__27474),
            .I(N__27466));
    Span4Mux_v I__4628 (
            .O(N__27469),
            .I(N__27461));
    Span4Mux_h I__4627 (
            .O(N__27466),
            .I(N__27461));
    Odrv4 I__4626 (
            .O(N__27461),
            .I(\current_shift_inst.elapsed_time_ns_phase_4 ));
    InMux I__4625 (
            .O(N__27458),
            .I(N__27455));
    LocalMux I__4624 (
            .O(N__27455),
            .I(N__27452));
    Span4Mux_h I__4623 (
            .O(N__27452),
            .I(N__27449));
    Odrv4 I__4622 (
            .O(N__27449),
            .I(\current_shift_inst.z_5_4 ));
    InMux I__4621 (
            .O(N__27446),
            .I(\current_shift_inst.z_5_cry_3 ));
    InMux I__4620 (
            .O(N__27443),
            .I(N__27440));
    LocalMux I__4619 (
            .O(N__27440),
            .I(G_406));
    CascadeMux I__4618 (
            .O(N__27437),
            .I(N__27434));
    InMux I__4617 (
            .O(N__27434),
            .I(N__27431));
    LocalMux I__4616 (
            .O(N__27431),
            .I(N__27428));
    Span4Mux_h I__4615 (
            .O(N__27428),
            .I(N__27425));
    Odrv4 I__4614 (
            .O(N__27425),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ));
    CascadeMux I__4613 (
            .O(N__27422),
            .I(N__27419));
    InMux I__4612 (
            .O(N__27419),
            .I(N__27416));
    LocalMux I__4611 (
            .O(N__27416),
            .I(N__27413));
    Odrv4 I__4610 (
            .O(N__27413),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ));
    CascadeMux I__4609 (
            .O(N__27410),
            .I(N__27407));
    InMux I__4608 (
            .O(N__27407),
            .I(N__27404));
    LocalMux I__4607 (
            .O(N__27404),
            .I(N__27401));
    Odrv4 I__4606 (
            .O(N__27401),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ));
    InMux I__4605 (
            .O(N__27398),
            .I(N__27394));
    InMux I__4604 (
            .O(N__27397),
            .I(N__27390));
    LocalMux I__4603 (
            .O(N__27394),
            .I(N__27386));
    InMux I__4602 (
            .O(N__27393),
            .I(N__27383));
    LocalMux I__4601 (
            .O(N__27390),
            .I(N__27380));
    InMux I__4600 (
            .O(N__27389),
            .I(N__27377));
    Odrv4 I__4599 (
            .O(N__27386),
            .I(\phase_controller_inst1.stoper_hc.time_passed11 ));
    LocalMux I__4598 (
            .O(N__27383),
            .I(\phase_controller_inst1.stoper_hc.time_passed11 ));
    Odrv12 I__4597 (
            .O(N__27380),
            .I(\phase_controller_inst1.stoper_hc.time_passed11 ));
    LocalMux I__4596 (
            .O(N__27377),
            .I(\phase_controller_inst1.stoper_hc.time_passed11 ));
    CascadeMux I__4595 (
            .O(N__27368),
            .I(N__27365));
    InMux I__4594 (
            .O(N__27365),
            .I(N__27362));
    LocalMux I__4593 (
            .O(N__27362),
            .I(N__27359));
    Odrv4 I__4592 (
            .O(N__27359),
            .I(\phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa ));
    CascadeMux I__4591 (
            .O(N__27356),
            .I(N__27353));
    InMux I__4590 (
            .O(N__27353),
            .I(N__27350));
    LocalMux I__4589 (
            .O(N__27350),
            .I(G_407));
    InMux I__4588 (
            .O(N__27347),
            .I(N__27342));
    InMux I__4587 (
            .O(N__27346),
            .I(N__27339));
    InMux I__4586 (
            .O(N__27345),
            .I(N__27336));
    LocalMux I__4585 (
            .O(N__27342),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    LocalMux I__4584 (
            .O(N__27339),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    LocalMux I__4583 (
            .O(N__27336),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    InMux I__4582 (
            .O(N__27329),
            .I(\pwm_generator_inst.counter_cry_5 ));
    InMux I__4581 (
            .O(N__27326),
            .I(N__27321));
    InMux I__4580 (
            .O(N__27325),
            .I(N__27318));
    InMux I__4579 (
            .O(N__27324),
            .I(N__27315));
    LocalMux I__4578 (
            .O(N__27321),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    LocalMux I__4577 (
            .O(N__27318),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    LocalMux I__4576 (
            .O(N__27315),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    InMux I__4575 (
            .O(N__27308),
            .I(\pwm_generator_inst.counter_cry_6 ));
    InMux I__4574 (
            .O(N__27305),
            .I(N__27300));
    InMux I__4573 (
            .O(N__27304),
            .I(N__27297));
    InMux I__4572 (
            .O(N__27303),
            .I(N__27294));
    LocalMux I__4571 (
            .O(N__27300),
            .I(N__27291));
    LocalMux I__4570 (
            .O(N__27297),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    LocalMux I__4569 (
            .O(N__27294),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    Odrv4 I__4568 (
            .O(N__27291),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    InMux I__4567 (
            .O(N__27284),
            .I(bfn_10_10_0_));
    InMux I__4566 (
            .O(N__27281),
            .I(N__27269));
    InMux I__4565 (
            .O(N__27280),
            .I(N__27266));
    InMux I__4564 (
            .O(N__27279),
            .I(N__27257));
    InMux I__4563 (
            .O(N__27278),
            .I(N__27257));
    InMux I__4562 (
            .O(N__27277),
            .I(N__27257));
    InMux I__4561 (
            .O(N__27276),
            .I(N__27257));
    InMux I__4560 (
            .O(N__27275),
            .I(N__27248));
    InMux I__4559 (
            .O(N__27274),
            .I(N__27248));
    InMux I__4558 (
            .O(N__27273),
            .I(N__27248));
    InMux I__4557 (
            .O(N__27272),
            .I(N__27248));
    LocalMux I__4556 (
            .O(N__27269),
            .I(N__27245));
    LocalMux I__4555 (
            .O(N__27266),
            .I(N__27242));
    LocalMux I__4554 (
            .O(N__27257),
            .I(\pwm_generator_inst.un1_counter_0 ));
    LocalMux I__4553 (
            .O(N__27248),
            .I(\pwm_generator_inst.un1_counter_0 ));
    Odrv12 I__4552 (
            .O(N__27245),
            .I(\pwm_generator_inst.un1_counter_0 ));
    Odrv4 I__4551 (
            .O(N__27242),
            .I(\pwm_generator_inst.un1_counter_0 ));
    InMux I__4550 (
            .O(N__27233),
            .I(\pwm_generator_inst.counter_cry_8 ));
    InMux I__4549 (
            .O(N__27230),
            .I(N__27225));
    InMux I__4548 (
            .O(N__27229),
            .I(N__27222));
    InMux I__4547 (
            .O(N__27228),
            .I(N__27219));
    LocalMux I__4546 (
            .O(N__27225),
            .I(N__27216));
    LocalMux I__4545 (
            .O(N__27222),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    LocalMux I__4544 (
            .O(N__27219),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    Odrv4 I__4543 (
            .O(N__27216),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    CascadeMux I__4542 (
            .O(N__27209),
            .I(\pwm_generator_inst.un1_counterlto2_0_cascade_ ));
    CascadeMux I__4541 (
            .O(N__27206),
            .I(\pwm_generator_inst.un1_counterlt9_cascade_ ));
    InMux I__4540 (
            .O(N__27203),
            .I(N__27200));
    LocalMux I__4539 (
            .O(N__27200),
            .I(\pwm_generator_inst.un1_counterlto9_2 ));
    InMux I__4538 (
            .O(N__27197),
            .I(N__27192));
    InMux I__4537 (
            .O(N__27196),
            .I(N__27189));
    InMux I__4536 (
            .O(N__27195),
            .I(N__27186));
    LocalMux I__4535 (
            .O(N__27192),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    LocalMux I__4534 (
            .O(N__27189),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    LocalMux I__4533 (
            .O(N__27186),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    InMux I__4532 (
            .O(N__27179),
            .I(bfn_10_9_0_));
    InMux I__4531 (
            .O(N__27176),
            .I(N__27171));
    InMux I__4530 (
            .O(N__27175),
            .I(N__27168));
    InMux I__4529 (
            .O(N__27174),
            .I(N__27165));
    LocalMux I__4528 (
            .O(N__27171),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    LocalMux I__4527 (
            .O(N__27168),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    LocalMux I__4526 (
            .O(N__27165),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    InMux I__4525 (
            .O(N__27158),
            .I(\pwm_generator_inst.counter_cry_0 ));
    InMux I__4524 (
            .O(N__27155),
            .I(N__27150));
    InMux I__4523 (
            .O(N__27154),
            .I(N__27147));
    InMux I__4522 (
            .O(N__27153),
            .I(N__27144));
    LocalMux I__4521 (
            .O(N__27150),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    LocalMux I__4520 (
            .O(N__27147),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    LocalMux I__4519 (
            .O(N__27144),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    InMux I__4518 (
            .O(N__27137),
            .I(\pwm_generator_inst.counter_cry_1 ));
    InMux I__4517 (
            .O(N__27134),
            .I(N__27129));
    InMux I__4516 (
            .O(N__27133),
            .I(N__27126));
    InMux I__4515 (
            .O(N__27132),
            .I(N__27123));
    LocalMux I__4514 (
            .O(N__27129),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    LocalMux I__4513 (
            .O(N__27126),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    LocalMux I__4512 (
            .O(N__27123),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    InMux I__4511 (
            .O(N__27116),
            .I(\pwm_generator_inst.counter_cry_2 ));
    InMux I__4510 (
            .O(N__27113),
            .I(N__27108));
    InMux I__4509 (
            .O(N__27112),
            .I(N__27105));
    InMux I__4508 (
            .O(N__27111),
            .I(N__27102));
    LocalMux I__4507 (
            .O(N__27108),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    LocalMux I__4506 (
            .O(N__27105),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    LocalMux I__4505 (
            .O(N__27102),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    InMux I__4504 (
            .O(N__27095),
            .I(\pwm_generator_inst.counter_cry_3 ));
    InMux I__4503 (
            .O(N__27092),
            .I(N__27087));
    InMux I__4502 (
            .O(N__27091),
            .I(N__27084));
    InMux I__4501 (
            .O(N__27090),
            .I(N__27081));
    LocalMux I__4500 (
            .O(N__27087),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    LocalMux I__4499 (
            .O(N__27084),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    LocalMux I__4498 (
            .O(N__27081),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    InMux I__4497 (
            .O(N__27074),
            .I(\pwm_generator_inst.counter_cry_4 ));
    InMux I__4496 (
            .O(N__27071),
            .I(N__27067));
    InMux I__4495 (
            .O(N__27070),
            .I(N__27064));
    LocalMux I__4494 (
            .O(N__27067),
            .I(N__27058));
    LocalMux I__4493 (
            .O(N__27064),
            .I(N__27058));
    InMux I__4492 (
            .O(N__27063),
            .I(N__27055));
    Span4Mux_v I__4491 (
            .O(N__27058),
            .I(N__27052));
    LocalMux I__4490 (
            .O(N__27055),
            .I(\current_shift_inst.timer_phase.counterZ0Z_24 ));
    Odrv4 I__4489 (
            .O(N__27052),
            .I(\current_shift_inst.timer_phase.counterZ0Z_24 ));
    InMux I__4488 (
            .O(N__27047),
            .I(bfn_9_28_0_));
    InMux I__4487 (
            .O(N__27044),
            .I(N__27040));
    InMux I__4486 (
            .O(N__27043),
            .I(N__27037));
    LocalMux I__4485 (
            .O(N__27040),
            .I(N__27031));
    LocalMux I__4484 (
            .O(N__27037),
            .I(N__27031));
    InMux I__4483 (
            .O(N__27036),
            .I(N__27028));
    Span4Mux_v I__4482 (
            .O(N__27031),
            .I(N__27025));
    LocalMux I__4481 (
            .O(N__27028),
            .I(\current_shift_inst.timer_phase.counterZ0Z_25 ));
    Odrv4 I__4480 (
            .O(N__27025),
            .I(\current_shift_inst.timer_phase.counterZ0Z_25 ));
    InMux I__4479 (
            .O(N__27020),
            .I(\current_shift_inst.timer_phase.counter_cry_24 ));
    CascadeMux I__4478 (
            .O(N__27017),
            .I(N__27013));
    CascadeMux I__4477 (
            .O(N__27016),
            .I(N__27010));
    InMux I__4476 (
            .O(N__27013),
            .I(N__27005));
    InMux I__4475 (
            .O(N__27010),
            .I(N__27005));
    LocalMux I__4474 (
            .O(N__27005),
            .I(N__27001));
    InMux I__4473 (
            .O(N__27004),
            .I(N__26998));
    Span4Mux_h I__4472 (
            .O(N__27001),
            .I(N__26995));
    LocalMux I__4471 (
            .O(N__26998),
            .I(\current_shift_inst.timer_phase.counterZ0Z_26 ));
    Odrv4 I__4470 (
            .O(N__26995),
            .I(\current_shift_inst.timer_phase.counterZ0Z_26 ));
    InMux I__4469 (
            .O(N__26990),
            .I(\current_shift_inst.timer_phase.counter_cry_25 ));
    CascadeMux I__4468 (
            .O(N__26987),
            .I(N__26983));
    CascadeMux I__4467 (
            .O(N__26986),
            .I(N__26980));
    InMux I__4466 (
            .O(N__26983),
            .I(N__26974));
    InMux I__4465 (
            .O(N__26980),
            .I(N__26974));
    InMux I__4464 (
            .O(N__26979),
            .I(N__26971));
    LocalMux I__4463 (
            .O(N__26974),
            .I(N__26968));
    LocalMux I__4462 (
            .O(N__26971),
            .I(\current_shift_inst.timer_phase.counterZ0Z_27 ));
    Odrv12 I__4461 (
            .O(N__26968),
            .I(\current_shift_inst.timer_phase.counterZ0Z_27 ));
    InMux I__4460 (
            .O(N__26963),
            .I(\current_shift_inst.timer_phase.counter_cry_26 ));
    InMux I__4459 (
            .O(N__26960),
            .I(N__26957));
    LocalMux I__4458 (
            .O(N__26957),
            .I(N__26953));
    InMux I__4457 (
            .O(N__26956),
            .I(N__26950));
    Span4Mux_h I__4456 (
            .O(N__26953),
            .I(N__26947));
    LocalMux I__4455 (
            .O(N__26950),
            .I(\current_shift_inst.timer_phase.counterZ0Z_28 ));
    Odrv4 I__4454 (
            .O(N__26947),
            .I(\current_shift_inst.timer_phase.counterZ0Z_28 ));
    InMux I__4453 (
            .O(N__26942),
            .I(\current_shift_inst.timer_phase.counter_cry_27 ));
    InMux I__4452 (
            .O(N__26939),
            .I(\current_shift_inst.timer_phase.counter_cry_28 ));
    InMux I__4451 (
            .O(N__26936),
            .I(N__26932));
    InMux I__4450 (
            .O(N__26935),
            .I(N__26929));
    LocalMux I__4449 (
            .O(N__26932),
            .I(N__26926));
    LocalMux I__4448 (
            .O(N__26929),
            .I(\current_shift_inst.timer_phase.counterZ0Z_29 ));
    Odrv12 I__4447 (
            .O(N__26926),
            .I(\current_shift_inst.timer_phase.counterZ0Z_29 ));
    InMux I__4446 (
            .O(N__26921),
            .I(N__26918));
    LocalMux I__4445 (
            .O(N__26918),
            .I(il_max_comp1_D1));
    InMux I__4444 (
            .O(N__26915),
            .I(N__26911));
    InMux I__4443 (
            .O(N__26914),
            .I(N__26908));
    LocalMux I__4442 (
            .O(N__26911),
            .I(N__26902));
    LocalMux I__4441 (
            .O(N__26908),
            .I(N__26902));
    InMux I__4440 (
            .O(N__26907),
            .I(N__26899));
    Span4Mux_v I__4439 (
            .O(N__26902),
            .I(N__26896));
    LocalMux I__4438 (
            .O(N__26899),
            .I(\current_shift_inst.timer_phase.counterZ0Z_16 ));
    Odrv4 I__4437 (
            .O(N__26896),
            .I(\current_shift_inst.timer_phase.counterZ0Z_16 ));
    InMux I__4436 (
            .O(N__26891),
            .I(bfn_9_27_0_));
    InMux I__4435 (
            .O(N__26888),
            .I(N__26884));
    InMux I__4434 (
            .O(N__26887),
            .I(N__26881));
    LocalMux I__4433 (
            .O(N__26884),
            .I(N__26875));
    LocalMux I__4432 (
            .O(N__26881),
            .I(N__26875));
    InMux I__4431 (
            .O(N__26880),
            .I(N__26872));
    Span4Mux_v I__4430 (
            .O(N__26875),
            .I(N__26869));
    LocalMux I__4429 (
            .O(N__26872),
            .I(\current_shift_inst.timer_phase.counterZ0Z_17 ));
    Odrv4 I__4428 (
            .O(N__26869),
            .I(\current_shift_inst.timer_phase.counterZ0Z_17 ));
    InMux I__4427 (
            .O(N__26864),
            .I(\current_shift_inst.timer_phase.counter_cry_16 ));
    CascadeMux I__4426 (
            .O(N__26861),
            .I(N__26857));
    CascadeMux I__4425 (
            .O(N__26860),
            .I(N__26854));
    InMux I__4424 (
            .O(N__26857),
            .I(N__26849));
    InMux I__4423 (
            .O(N__26854),
            .I(N__26849));
    LocalMux I__4422 (
            .O(N__26849),
            .I(N__26845));
    InMux I__4421 (
            .O(N__26848),
            .I(N__26842));
    Span4Mux_h I__4420 (
            .O(N__26845),
            .I(N__26839));
    LocalMux I__4419 (
            .O(N__26842),
            .I(\current_shift_inst.timer_phase.counterZ0Z_18 ));
    Odrv4 I__4418 (
            .O(N__26839),
            .I(\current_shift_inst.timer_phase.counterZ0Z_18 ));
    InMux I__4417 (
            .O(N__26834),
            .I(\current_shift_inst.timer_phase.counter_cry_17 ));
    CascadeMux I__4416 (
            .O(N__26831),
            .I(N__26827));
    CascadeMux I__4415 (
            .O(N__26830),
            .I(N__26824));
    InMux I__4414 (
            .O(N__26827),
            .I(N__26819));
    InMux I__4413 (
            .O(N__26824),
            .I(N__26819));
    LocalMux I__4412 (
            .O(N__26819),
            .I(N__26815));
    InMux I__4411 (
            .O(N__26818),
            .I(N__26812));
    Span4Mux_h I__4410 (
            .O(N__26815),
            .I(N__26809));
    LocalMux I__4409 (
            .O(N__26812),
            .I(\current_shift_inst.timer_phase.counterZ0Z_19 ));
    Odrv4 I__4408 (
            .O(N__26809),
            .I(\current_shift_inst.timer_phase.counterZ0Z_19 ));
    InMux I__4407 (
            .O(N__26804),
            .I(\current_shift_inst.timer_phase.counter_cry_18 ));
    InMux I__4406 (
            .O(N__26801),
            .I(N__26795));
    InMux I__4405 (
            .O(N__26800),
            .I(N__26795));
    LocalMux I__4404 (
            .O(N__26795),
            .I(N__26791));
    InMux I__4403 (
            .O(N__26794),
            .I(N__26788));
    Span4Mux_h I__4402 (
            .O(N__26791),
            .I(N__26785));
    LocalMux I__4401 (
            .O(N__26788),
            .I(\current_shift_inst.timer_phase.counterZ0Z_20 ));
    Odrv4 I__4400 (
            .O(N__26785),
            .I(\current_shift_inst.timer_phase.counterZ0Z_20 ));
    InMux I__4399 (
            .O(N__26780),
            .I(\current_shift_inst.timer_phase.counter_cry_19 ));
    InMux I__4398 (
            .O(N__26777),
            .I(N__26771));
    InMux I__4397 (
            .O(N__26776),
            .I(N__26771));
    LocalMux I__4396 (
            .O(N__26771),
            .I(N__26767));
    InMux I__4395 (
            .O(N__26770),
            .I(N__26764));
    Span4Mux_h I__4394 (
            .O(N__26767),
            .I(N__26761));
    LocalMux I__4393 (
            .O(N__26764),
            .I(\current_shift_inst.timer_phase.counterZ0Z_21 ));
    Odrv4 I__4392 (
            .O(N__26761),
            .I(\current_shift_inst.timer_phase.counterZ0Z_21 ));
    InMux I__4391 (
            .O(N__26756),
            .I(\current_shift_inst.timer_phase.counter_cry_20 ));
    CascadeMux I__4390 (
            .O(N__26753),
            .I(N__26749));
    CascadeMux I__4389 (
            .O(N__26752),
            .I(N__26746));
    InMux I__4388 (
            .O(N__26749),
            .I(N__26741));
    InMux I__4387 (
            .O(N__26746),
            .I(N__26741));
    LocalMux I__4386 (
            .O(N__26741),
            .I(N__26737));
    InMux I__4385 (
            .O(N__26740),
            .I(N__26734));
    Span4Mux_v I__4384 (
            .O(N__26737),
            .I(N__26731));
    LocalMux I__4383 (
            .O(N__26734),
            .I(\current_shift_inst.timer_phase.counterZ0Z_22 ));
    Odrv4 I__4382 (
            .O(N__26731),
            .I(\current_shift_inst.timer_phase.counterZ0Z_22 ));
    InMux I__4381 (
            .O(N__26726),
            .I(\current_shift_inst.timer_phase.counter_cry_21 ));
    CascadeMux I__4380 (
            .O(N__26723),
            .I(N__26719));
    CascadeMux I__4379 (
            .O(N__26722),
            .I(N__26716));
    InMux I__4378 (
            .O(N__26719),
            .I(N__26710));
    InMux I__4377 (
            .O(N__26716),
            .I(N__26710));
    InMux I__4376 (
            .O(N__26715),
            .I(N__26707));
    LocalMux I__4375 (
            .O(N__26710),
            .I(N__26704));
    LocalMux I__4374 (
            .O(N__26707),
            .I(\current_shift_inst.timer_phase.counterZ0Z_23 ));
    Odrv12 I__4373 (
            .O(N__26704),
            .I(\current_shift_inst.timer_phase.counterZ0Z_23 ));
    InMux I__4372 (
            .O(N__26699),
            .I(\current_shift_inst.timer_phase.counter_cry_22 ));
    CascadeMux I__4371 (
            .O(N__26696),
            .I(N__26692));
    InMux I__4370 (
            .O(N__26695),
            .I(N__26689));
    InMux I__4369 (
            .O(N__26692),
            .I(N__26686));
    LocalMux I__4368 (
            .O(N__26689),
            .I(N__26680));
    LocalMux I__4367 (
            .O(N__26686),
            .I(N__26680));
    InMux I__4366 (
            .O(N__26685),
            .I(N__26677));
    Span4Mux_v I__4365 (
            .O(N__26680),
            .I(N__26674));
    LocalMux I__4364 (
            .O(N__26677),
            .I(\current_shift_inst.timer_phase.counterZ0Z_8 ));
    Odrv4 I__4363 (
            .O(N__26674),
            .I(\current_shift_inst.timer_phase.counterZ0Z_8 ));
    InMux I__4362 (
            .O(N__26669),
            .I(bfn_9_26_0_));
    InMux I__4361 (
            .O(N__26666),
            .I(N__26662));
    InMux I__4360 (
            .O(N__26665),
            .I(N__26659));
    LocalMux I__4359 (
            .O(N__26662),
            .I(N__26653));
    LocalMux I__4358 (
            .O(N__26659),
            .I(N__26653));
    InMux I__4357 (
            .O(N__26658),
            .I(N__26650));
    Span4Mux_v I__4356 (
            .O(N__26653),
            .I(N__26647));
    LocalMux I__4355 (
            .O(N__26650),
            .I(\current_shift_inst.timer_phase.counterZ0Z_9 ));
    Odrv4 I__4354 (
            .O(N__26647),
            .I(\current_shift_inst.timer_phase.counterZ0Z_9 ));
    InMux I__4353 (
            .O(N__26642),
            .I(\current_shift_inst.timer_phase.counter_cry_8 ));
    CascadeMux I__4352 (
            .O(N__26639),
            .I(N__26635));
    CascadeMux I__4351 (
            .O(N__26638),
            .I(N__26632));
    InMux I__4350 (
            .O(N__26635),
            .I(N__26627));
    InMux I__4349 (
            .O(N__26632),
            .I(N__26627));
    LocalMux I__4348 (
            .O(N__26627),
            .I(N__26623));
    InMux I__4347 (
            .O(N__26626),
            .I(N__26620));
    Span4Mux_h I__4346 (
            .O(N__26623),
            .I(N__26617));
    LocalMux I__4345 (
            .O(N__26620),
            .I(\current_shift_inst.timer_phase.counterZ0Z_10 ));
    Odrv4 I__4344 (
            .O(N__26617),
            .I(\current_shift_inst.timer_phase.counterZ0Z_10 ));
    InMux I__4343 (
            .O(N__26612),
            .I(\current_shift_inst.timer_phase.counter_cry_9 ));
    CascadeMux I__4342 (
            .O(N__26609),
            .I(N__26605));
    CascadeMux I__4341 (
            .O(N__26608),
            .I(N__26602));
    InMux I__4340 (
            .O(N__26605),
            .I(N__26596));
    InMux I__4339 (
            .O(N__26602),
            .I(N__26596));
    InMux I__4338 (
            .O(N__26601),
            .I(N__26593));
    LocalMux I__4337 (
            .O(N__26596),
            .I(N__26590));
    LocalMux I__4336 (
            .O(N__26593),
            .I(\current_shift_inst.timer_phase.counterZ0Z_11 ));
    Odrv12 I__4335 (
            .O(N__26590),
            .I(\current_shift_inst.timer_phase.counterZ0Z_11 ));
    InMux I__4334 (
            .O(N__26585),
            .I(\current_shift_inst.timer_phase.counter_cry_10 ));
    InMux I__4333 (
            .O(N__26582),
            .I(N__26575));
    InMux I__4332 (
            .O(N__26581),
            .I(N__26575));
    InMux I__4331 (
            .O(N__26580),
            .I(N__26572));
    LocalMux I__4330 (
            .O(N__26575),
            .I(N__26569));
    LocalMux I__4329 (
            .O(N__26572),
            .I(\current_shift_inst.timer_phase.counterZ0Z_12 ));
    Odrv12 I__4328 (
            .O(N__26569),
            .I(\current_shift_inst.timer_phase.counterZ0Z_12 ));
    InMux I__4327 (
            .O(N__26564),
            .I(\current_shift_inst.timer_phase.counter_cry_11 ));
    InMux I__4326 (
            .O(N__26561),
            .I(N__26555));
    InMux I__4325 (
            .O(N__26560),
            .I(N__26555));
    LocalMux I__4324 (
            .O(N__26555),
            .I(N__26551));
    InMux I__4323 (
            .O(N__26554),
            .I(N__26548));
    Span4Mux_h I__4322 (
            .O(N__26551),
            .I(N__26545));
    LocalMux I__4321 (
            .O(N__26548),
            .I(\current_shift_inst.timer_phase.counterZ0Z_13 ));
    Odrv4 I__4320 (
            .O(N__26545),
            .I(\current_shift_inst.timer_phase.counterZ0Z_13 ));
    InMux I__4319 (
            .O(N__26540),
            .I(\current_shift_inst.timer_phase.counter_cry_12 ));
    CascadeMux I__4318 (
            .O(N__26537),
            .I(N__26533));
    CascadeMux I__4317 (
            .O(N__26536),
            .I(N__26530));
    InMux I__4316 (
            .O(N__26533),
            .I(N__26524));
    InMux I__4315 (
            .O(N__26530),
            .I(N__26524));
    InMux I__4314 (
            .O(N__26529),
            .I(N__26521));
    LocalMux I__4313 (
            .O(N__26524),
            .I(N__26518));
    LocalMux I__4312 (
            .O(N__26521),
            .I(\current_shift_inst.timer_phase.counterZ0Z_14 ));
    Odrv12 I__4311 (
            .O(N__26518),
            .I(\current_shift_inst.timer_phase.counterZ0Z_14 ));
    InMux I__4310 (
            .O(N__26513),
            .I(\current_shift_inst.timer_phase.counter_cry_13 ));
    CascadeMux I__4309 (
            .O(N__26510),
            .I(N__26506));
    CascadeMux I__4308 (
            .O(N__26509),
            .I(N__26503));
    InMux I__4307 (
            .O(N__26506),
            .I(N__26498));
    InMux I__4306 (
            .O(N__26503),
            .I(N__26498));
    LocalMux I__4305 (
            .O(N__26498),
            .I(N__26494));
    InMux I__4304 (
            .O(N__26497),
            .I(N__26491));
    Span4Mux_v I__4303 (
            .O(N__26494),
            .I(N__26488));
    LocalMux I__4302 (
            .O(N__26491),
            .I(\current_shift_inst.timer_phase.counterZ0Z_15 ));
    Odrv4 I__4301 (
            .O(N__26488),
            .I(\current_shift_inst.timer_phase.counterZ0Z_15 ));
    InMux I__4300 (
            .O(N__26483),
            .I(\current_shift_inst.timer_phase.counter_cry_14 ));
    InMux I__4299 (
            .O(N__26480),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_29 ));
    CEMux I__4298 (
            .O(N__26477),
            .I(N__26462));
    CEMux I__4297 (
            .O(N__26476),
            .I(N__26462));
    CEMux I__4296 (
            .O(N__26475),
            .I(N__26462));
    CEMux I__4295 (
            .O(N__26474),
            .I(N__26462));
    CEMux I__4294 (
            .O(N__26473),
            .I(N__26462));
    GlobalMux I__4293 (
            .O(N__26462),
            .I(N__26459));
    gio2CtrlBuf I__4292 (
            .O(N__26459),
            .I(\current_shift_inst.timer_phase.N_188_i_g ));
    InMux I__4291 (
            .O(N__26456),
            .I(N__26452));
    InMux I__4290 (
            .O(N__26455),
            .I(N__26449));
    LocalMux I__4289 (
            .O(N__26452),
            .I(N__26446));
    LocalMux I__4288 (
            .O(N__26449),
            .I(N__26443));
    Span12Mux_v I__4287 (
            .O(N__26446),
            .I(N__26439));
    Span4Mux_h I__4286 (
            .O(N__26443),
            .I(N__26436));
    InMux I__4285 (
            .O(N__26442),
            .I(N__26433));
    Odrv12 I__4284 (
            .O(N__26439),
            .I(\current_shift_inst.timer_phase.counterZ0Z_0 ));
    Odrv4 I__4283 (
            .O(N__26436),
            .I(\current_shift_inst.timer_phase.counterZ0Z_0 ));
    LocalMux I__4282 (
            .O(N__26433),
            .I(\current_shift_inst.timer_phase.counterZ0Z_0 ));
    InMux I__4281 (
            .O(N__26426),
            .I(bfn_9_25_0_));
    InMux I__4280 (
            .O(N__26423),
            .I(N__26419));
    InMux I__4279 (
            .O(N__26422),
            .I(N__26416));
    LocalMux I__4278 (
            .O(N__26419),
            .I(N__26410));
    LocalMux I__4277 (
            .O(N__26416),
            .I(N__26410));
    InMux I__4276 (
            .O(N__26415),
            .I(N__26407));
    Odrv12 I__4275 (
            .O(N__26410),
            .I(\current_shift_inst.timer_phase.counterZ0Z_1 ));
    LocalMux I__4274 (
            .O(N__26407),
            .I(\current_shift_inst.timer_phase.counterZ0Z_1 ));
    InMux I__4273 (
            .O(N__26402),
            .I(\current_shift_inst.timer_phase.counter_cry_0 ));
    CascadeMux I__4272 (
            .O(N__26399),
            .I(N__26395));
    CascadeMux I__4271 (
            .O(N__26398),
            .I(N__26392));
    InMux I__4270 (
            .O(N__26395),
            .I(N__26386));
    InMux I__4269 (
            .O(N__26392),
            .I(N__26386));
    InMux I__4268 (
            .O(N__26391),
            .I(N__26383));
    LocalMux I__4267 (
            .O(N__26386),
            .I(N__26380));
    LocalMux I__4266 (
            .O(N__26383),
            .I(\current_shift_inst.timer_phase.counterZ0Z_2 ));
    Odrv12 I__4265 (
            .O(N__26380),
            .I(\current_shift_inst.timer_phase.counterZ0Z_2 ));
    InMux I__4264 (
            .O(N__26375),
            .I(\current_shift_inst.timer_phase.counter_cry_1 ));
    CascadeMux I__4263 (
            .O(N__26372),
            .I(N__26368));
    CascadeMux I__4262 (
            .O(N__26371),
            .I(N__26365));
    InMux I__4261 (
            .O(N__26368),
            .I(N__26360));
    InMux I__4260 (
            .O(N__26365),
            .I(N__26360));
    LocalMux I__4259 (
            .O(N__26360),
            .I(N__26356));
    InMux I__4258 (
            .O(N__26359),
            .I(N__26353));
    Span4Mux_h I__4257 (
            .O(N__26356),
            .I(N__26350));
    LocalMux I__4256 (
            .O(N__26353),
            .I(\current_shift_inst.timer_phase.counterZ0Z_3 ));
    Odrv4 I__4255 (
            .O(N__26350),
            .I(\current_shift_inst.timer_phase.counterZ0Z_3 ));
    InMux I__4254 (
            .O(N__26345),
            .I(\current_shift_inst.timer_phase.counter_cry_2 ));
    InMux I__4253 (
            .O(N__26342),
            .I(N__26335));
    InMux I__4252 (
            .O(N__26341),
            .I(N__26335));
    InMux I__4251 (
            .O(N__26340),
            .I(N__26332));
    LocalMux I__4250 (
            .O(N__26335),
            .I(N__26329));
    LocalMux I__4249 (
            .O(N__26332),
            .I(\current_shift_inst.timer_phase.counterZ0Z_4 ));
    Odrv12 I__4248 (
            .O(N__26329),
            .I(\current_shift_inst.timer_phase.counterZ0Z_4 ));
    InMux I__4247 (
            .O(N__26324),
            .I(\current_shift_inst.timer_phase.counter_cry_3 ));
    InMux I__4246 (
            .O(N__26321),
            .I(N__26315));
    InMux I__4245 (
            .O(N__26320),
            .I(N__26315));
    LocalMux I__4244 (
            .O(N__26315),
            .I(N__26311));
    InMux I__4243 (
            .O(N__26314),
            .I(N__26308));
    Span4Mux_h I__4242 (
            .O(N__26311),
            .I(N__26305));
    LocalMux I__4241 (
            .O(N__26308),
            .I(\current_shift_inst.timer_phase.counterZ0Z_5 ));
    Odrv4 I__4240 (
            .O(N__26305),
            .I(\current_shift_inst.timer_phase.counterZ0Z_5 ));
    InMux I__4239 (
            .O(N__26300),
            .I(\current_shift_inst.timer_phase.counter_cry_4 ));
    CascadeMux I__4238 (
            .O(N__26297),
            .I(N__26293));
    InMux I__4237 (
            .O(N__26296),
            .I(N__26290));
    InMux I__4236 (
            .O(N__26293),
            .I(N__26287));
    LocalMux I__4235 (
            .O(N__26290),
            .I(N__26283));
    LocalMux I__4234 (
            .O(N__26287),
            .I(N__26280));
    InMux I__4233 (
            .O(N__26286),
            .I(N__26277));
    Span4Mux_v I__4232 (
            .O(N__26283),
            .I(N__26272));
    Span4Mux_v I__4231 (
            .O(N__26280),
            .I(N__26272));
    LocalMux I__4230 (
            .O(N__26277),
            .I(\current_shift_inst.timer_phase.counterZ0Z_6 ));
    Odrv4 I__4229 (
            .O(N__26272),
            .I(\current_shift_inst.timer_phase.counterZ0Z_6 ));
    InMux I__4228 (
            .O(N__26267),
            .I(\current_shift_inst.timer_phase.counter_cry_5 ));
    CascadeMux I__4227 (
            .O(N__26264),
            .I(N__26260));
    CascadeMux I__4226 (
            .O(N__26263),
            .I(N__26257));
    InMux I__4225 (
            .O(N__26260),
            .I(N__26251));
    InMux I__4224 (
            .O(N__26257),
            .I(N__26251));
    InMux I__4223 (
            .O(N__26256),
            .I(N__26248));
    LocalMux I__4222 (
            .O(N__26251),
            .I(N__26245));
    LocalMux I__4221 (
            .O(N__26248),
            .I(\current_shift_inst.timer_phase.counterZ0Z_7 ));
    Odrv12 I__4220 (
            .O(N__26245),
            .I(\current_shift_inst.timer_phase.counterZ0Z_7 ));
    InMux I__4219 (
            .O(N__26240),
            .I(\current_shift_inst.timer_phase.counter_cry_6 ));
    InMux I__4218 (
            .O(N__26237),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_20 ));
    InMux I__4217 (
            .O(N__26234),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_21 ));
    InMux I__4216 (
            .O(N__26231),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_22 ));
    InMux I__4215 (
            .O(N__26228),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_23 ));
    InMux I__4214 (
            .O(N__26225),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_24 ));
    InMux I__4213 (
            .O(N__26222),
            .I(bfn_9_24_0_));
    InMux I__4212 (
            .O(N__26219),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_26 ));
    InMux I__4211 (
            .O(N__26216),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_27 ));
    InMux I__4210 (
            .O(N__26213),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_28 ));
    InMux I__4209 (
            .O(N__26210),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_11 ));
    InMux I__4208 (
            .O(N__26207),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_12 ));
    InMux I__4207 (
            .O(N__26204),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_13 ));
    InMux I__4206 (
            .O(N__26201),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_14 ));
    InMux I__4205 (
            .O(N__26198),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_15 ));
    InMux I__4204 (
            .O(N__26195),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_16 ));
    InMux I__4203 (
            .O(N__26192),
            .I(bfn_9_23_0_));
    InMux I__4202 (
            .O(N__26189),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_18 ));
    InMux I__4201 (
            .O(N__26186),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_19 ));
    InMux I__4200 (
            .O(N__26183),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_2 ));
    InMux I__4199 (
            .O(N__26180),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_3 ));
    InMux I__4198 (
            .O(N__26177),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_4 ));
    InMux I__4197 (
            .O(N__26174),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_5 ));
    InMux I__4196 (
            .O(N__26171),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_6 ));
    InMux I__4195 (
            .O(N__26168),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_7 ));
    InMux I__4194 (
            .O(N__26165),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_8 ));
    InMux I__4193 (
            .O(N__26162),
            .I(bfn_9_22_0_));
    InMux I__4192 (
            .O(N__26159),
            .I(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__4191 (
            .O(N__26156),
            .I(N__26153));
    InMux I__4190 (
            .O(N__26153),
            .I(N__26150));
    LocalMux I__4189 (
            .O(N__26150),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIR32K_22 ));
    InMux I__4188 (
            .O(N__26147),
            .I(N__26144));
    LocalMux I__4187 (
            .O(N__26144),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPB581_22 ));
    InMux I__4186 (
            .O(N__26141),
            .I(N__26138));
    LocalMux I__4185 (
            .O(N__26138),
            .I(N__26135));
    Odrv4 I__4184 (
            .O(N__26135),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJ3381_21 ));
    InMux I__4183 (
            .O(N__26132),
            .I(N__26129));
    LocalMux I__4182 (
            .O(N__26129),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIVQF91_30 ));
    CascadeMux I__4181 (
            .O(N__26126),
            .I(N__26123));
    InMux I__4180 (
            .O(N__26123),
            .I(N__26120));
    LocalMux I__4179 (
            .O(N__26120),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIAO7K_27 ));
    CascadeMux I__4178 (
            .O(N__26117),
            .I(N__26114));
    InMux I__4177 (
            .O(N__26114),
            .I(N__26111));
    LocalMux I__4176 (
            .O(N__26111),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI4D1J_16 ));
    InMux I__4175 (
            .O(N__26108),
            .I(N__26105));
    LocalMux I__4174 (
            .O(N__26105),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIKKJ81_29 ));
    InMux I__4173 (
            .O(N__26102),
            .I(N__26099));
    LocalMux I__4172 (
            .O(N__26099),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIHCE81_26 ));
    InMux I__4171 (
            .O(N__26096),
            .I(N__26093));
    LocalMux I__4170 (
            .O(N__26093),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI7DM51_10 ));
    InMux I__4169 (
            .O(N__26090),
            .I(N__26087));
    LocalMux I__4168 (
            .O(N__26087),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI53NU1_6 ));
    InMux I__4167 (
            .O(N__26084),
            .I(N__26081));
    LocalMux I__4166 (
            .O(N__26081),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI7H2J_17 ));
    CascadeMux I__4165 (
            .O(N__26078),
            .I(N__26075));
    InMux I__4164 (
            .O(N__26075),
            .I(N__26072));
    LocalMux I__4163 (
            .O(N__26072),
            .I(N__26069));
    Odrv4 I__4162 (
            .O(N__26069),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIIKQI_10 ));
    CascadeMux I__4161 (
            .O(N__26066),
            .I(N__26063));
    InMux I__4160 (
            .O(N__26063),
            .I(N__26060));
    LocalMux I__4159 (
            .O(N__26060),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIU4VI_14 ));
    InMux I__4158 (
            .O(N__26057),
            .I(N__26054));
    LocalMux I__4157 (
            .O(N__26054),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIBU361_16 ));
    InMux I__4156 (
            .O(N__26051),
            .I(N__26048));
    LocalMux I__4155 (
            .O(N__26048),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIBBPU1_7 ));
    InMux I__4154 (
            .O(N__26045),
            .I(N__26042));
    LocalMux I__4153 (
            .O(N__26042),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI1PG21_9 ));
    InMux I__4152 (
            .O(N__26039),
            .I(N__26036));
    LocalMux I__4151 (
            .O(N__26036),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINKG81_27 ));
    CascadeMux I__4150 (
            .O(N__26033),
            .I(N__26030));
    InMux I__4149 (
            .O(N__26030),
            .I(N__26027));
    LocalMux I__4148 (
            .O(N__26027),
            .I(\current_shift_inst.un38_control_input_0_cry_2_c_RNOZ0 ));
    CascadeMux I__4147 (
            .O(N__26024),
            .I(N__26021));
    InMux I__4146 (
            .O(N__26021),
            .I(N__26018));
    LocalMux I__4145 (
            .O(N__26018),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3 ));
    CascadeMux I__4144 (
            .O(N__26015),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3_cascade_ ));
    InMux I__4143 (
            .O(N__26012),
            .I(N__26009));
    LocalMux I__4142 (
            .O(N__26009),
            .I(\current_shift_inst.un38_control_input_0_cry_4_c_RNOZ0 ));
    CascadeMux I__4141 (
            .O(N__26006),
            .I(N__26003));
    InMux I__4140 (
            .O(N__26003),
            .I(N__26000));
    LocalMux I__4139 (
            .O(N__26000),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIK3CV_7 ));
    InMux I__4138 (
            .O(N__25997),
            .I(N__25994));
    LocalMux I__4137 (
            .O(N__25994),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP5T51_13 ));
    CascadeMux I__4136 (
            .O(N__25991),
            .I(N__25988));
    InMux I__4135 (
            .O(N__25988),
            .I(N__25985));
    LocalMux I__4134 (
            .O(N__25985),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIER9V_5 ));
    CascadeMux I__4133 (
            .O(N__25982),
            .I(N__25979));
    InMux I__4132 (
            .O(N__25979),
            .I(N__25976));
    LocalMux I__4131 (
            .O(N__25976),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJDBL1_10 ));
    InMux I__4130 (
            .O(N__25973),
            .I(N__25970));
    LocalMux I__4129 (
            .O(N__25970),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIE6961_18 ));
    CascadeMux I__4128 (
            .O(N__25967),
            .I(N__25964));
    InMux I__4127 (
            .O(N__25964),
            .I(N__25961));
    LocalMux I__4126 (
            .O(N__25961),
            .I(N__25958));
    Odrv4 I__4125 (
            .O(N__25958),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIHVAV_6 ));
    InMux I__4124 (
            .O(N__25955),
            .I(N__25951));
    InMux I__4123 (
            .O(N__25954),
            .I(N__25947));
    LocalMux I__4122 (
            .O(N__25951),
            .I(N__25943));
    InMux I__4121 (
            .O(N__25950),
            .I(N__25940));
    LocalMux I__4120 (
            .O(N__25947),
            .I(N__25937));
    InMux I__4119 (
            .O(N__25946),
            .I(N__25934));
    Span4Mux_h I__4118 (
            .O(N__25943),
            .I(N__25927));
    LocalMux I__4117 (
            .O(N__25940),
            .I(N__25927));
    Span4Mux_v I__4116 (
            .O(N__25937),
            .I(N__25927));
    LocalMux I__4115 (
            .O(N__25934),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    Odrv4 I__4114 (
            .O(N__25927),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    InMux I__4113 (
            .O(N__25922),
            .I(N__25919));
    LocalMux I__4112 (
            .O(N__25919),
            .I(N__25916));
    Span4Mux_h I__4111 (
            .O(N__25916),
            .I(N__25913));
    Odrv4 I__4110 (
            .O(N__25913),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ));
    InMux I__4109 (
            .O(N__25910),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ));
    InMux I__4108 (
            .O(N__25907),
            .I(N__25902));
    CascadeMux I__4107 (
            .O(N__25906),
            .I(N__25899));
    CascadeMux I__4106 (
            .O(N__25905),
            .I(N__25896));
    LocalMux I__4105 (
            .O(N__25902),
            .I(N__25893));
    InMux I__4104 (
            .O(N__25899),
            .I(N__25890));
    InMux I__4103 (
            .O(N__25896),
            .I(N__25887));
    Span4Mux_v I__4102 (
            .O(N__25893),
            .I(N__25883));
    LocalMux I__4101 (
            .O(N__25890),
            .I(N__25878));
    LocalMux I__4100 (
            .O(N__25887),
            .I(N__25878));
    InMux I__4099 (
            .O(N__25886),
            .I(N__25875));
    Span4Mux_h I__4098 (
            .O(N__25883),
            .I(N__25872));
    Odrv12 I__4097 (
            .O(N__25878),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    LocalMux I__4096 (
            .O(N__25875),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    Odrv4 I__4095 (
            .O(N__25872),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    InMux I__4094 (
            .O(N__25865),
            .I(N__25862));
    LocalMux I__4093 (
            .O(N__25862),
            .I(N__25859));
    Odrv4 I__4092 (
            .O(N__25859),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ));
    InMux I__4091 (
            .O(N__25856),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ));
    CascadeMux I__4090 (
            .O(N__25853),
            .I(N__25849));
    CascadeMux I__4089 (
            .O(N__25852),
            .I(N__25844));
    InMux I__4088 (
            .O(N__25849),
            .I(N__25841));
    InMux I__4087 (
            .O(N__25848),
            .I(N__25838));
    InMux I__4086 (
            .O(N__25847),
            .I(N__25835));
    InMux I__4085 (
            .O(N__25844),
            .I(N__25832));
    LocalMux I__4084 (
            .O(N__25841),
            .I(N__25829));
    LocalMux I__4083 (
            .O(N__25838),
            .I(N__25826));
    LocalMux I__4082 (
            .O(N__25835),
            .I(N__25823));
    LocalMux I__4081 (
            .O(N__25832),
            .I(N__25820));
    Span4Mux_h I__4080 (
            .O(N__25829),
            .I(N__25817));
    Odrv4 I__4079 (
            .O(N__25826),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    Odrv4 I__4078 (
            .O(N__25823),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    Odrv4 I__4077 (
            .O(N__25820),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    Odrv4 I__4076 (
            .O(N__25817),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    InMux I__4075 (
            .O(N__25808),
            .I(N__25805));
    LocalMux I__4074 (
            .O(N__25805),
            .I(N__25802));
    Odrv4 I__4073 (
            .O(N__25802),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ));
    InMux I__4072 (
            .O(N__25799),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ));
    CascadeMux I__4071 (
            .O(N__25796),
            .I(N__25792));
    CascadeMux I__4070 (
            .O(N__25795),
            .I(N__25788));
    InMux I__4069 (
            .O(N__25792),
            .I(N__25784));
    CascadeMux I__4068 (
            .O(N__25791),
            .I(N__25781));
    InMux I__4067 (
            .O(N__25788),
            .I(N__25778));
    CascadeMux I__4066 (
            .O(N__25787),
            .I(N__25775));
    LocalMux I__4065 (
            .O(N__25784),
            .I(N__25772));
    InMux I__4064 (
            .O(N__25781),
            .I(N__25769));
    LocalMux I__4063 (
            .O(N__25778),
            .I(N__25766));
    InMux I__4062 (
            .O(N__25775),
            .I(N__25763));
    Span4Mux_h I__4061 (
            .O(N__25772),
            .I(N__25760));
    LocalMux I__4060 (
            .O(N__25769),
            .I(N__25755));
    Span4Mux_h I__4059 (
            .O(N__25766),
            .I(N__25755));
    LocalMux I__4058 (
            .O(N__25763),
            .I(N__25752));
    Odrv4 I__4057 (
            .O(N__25760),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    Odrv4 I__4056 (
            .O(N__25755),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    Odrv4 I__4055 (
            .O(N__25752),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    InMux I__4054 (
            .O(N__25745),
            .I(N__25742));
    LocalMux I__4053 (
            .O(N__25742),
            .I(N__25739));
    Odrv12 I__4052 (
            .O(N__25739),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ));
    InMux I__4051 (
            .O(N__25736),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ));
    CascadeMux I__4050 (
            .O(N__25733),
            .I(N__25725));
    CascadeMux I__4049 (
            .O(N__25732),
            .I(N__25721));
    CascadeMux I__4048 (
            .O(N__25731),
            .I(N__25717));
    InMux I__4047 (
            .O(N__25730),
            .I(N__25714));
    InMux I__4046 (
            .O(N__25729),
            .I(N__25699));
    InMux I__4045 (
            .O(N__25728),
            .I(N__25699));
    InMux I__4044 (
            .O(N__25725),
            .I(N__25699));
    InMux I__4043 (
            .O(N__25724),
            .I(N__25699));
    InMux I__4042 (
            .O(N__25721),
            .I(N__25699));
    InMux I__4041 (
            .O(N__25720),
            .I(N__25699));
    InMux I__4040 (
            .O(N__25717),
            .I(N__25699));
    LocalMux I__4039 (
            .O(N__25714),
            .I(N__25696));
    LocalMux I__4038 (
            .O(N__25699),
            .I(N__25693));
    Span4Mux_h I__4037 (
            .O(N__25696),
            .I(N__25690));
    Span4Mux_v I__4036 (
            .O(N__25693),
            .I(N__25687));
    Odrv4 I__4035 (
            .O(N__25690),
            .I(\current_shift_inst.control_inputZ0Z_25 ));
    Odrv4 I__4034 (
            .O(N__25687),
            .I(\current_shift_inst.control_inputZ0Z_25 ));
    CascadeMux I__4033 (
            .O(N__25682),
            .I(N__25679));
    InMux I__4032 (
            .O(N__25679),
            .I(N__25659));
    InMux I__4031 (
            .O(N__25678),
            .I(N__25659));
    CascadeMux I__4030 (
            .O(N__25677),
            .I(N__25655));
    CascadeMux I__4029 (
            .O(N__25676),
            .I(N__25650));
    CascadeMux I__4028 (
            .O(N__25675),
            .I(N__25646));
    CascadeMux I__4027 (
            .O(N__25674),
            .I(N__25642));
    CascadeMux I__4026 (
            .O(N__25673),
            .I(N__25639));
    CascadeMux I__4025 (
            .O(N__25672),
            .I(N__25636));
    CascadeMux I__4024 (
            .O(N__25671),
            .I(N__25629));
    CascadeMux I__4023 (
            .O(N__25670),
            .I(N__25626));
    CascadeMux I__4022 (
            .O(N__25669),
            .I(N__25623));
    CascadeMux I__4021 (
            .O(N__25668),
            .I(N__25620));
    CascadeMux I__4020 (
            .O(N__25667),
            .I(N__25615));
    CascadeMux I__4019 (
            .O(N__25666),
            .I(N__25610));
    CascadeMux I__4018 (
            .O(N__25665),
            .I(N__25607));
    CascadeMux I__4017 (
            .O(N__25664),
            .I(N__25604));
    LocalMux I__4016 (
            .O(N__25659),
            .I(N__25598));
    InMux I__4015 (
            .O(N__25658),
            .I(N__25595));
    InMux I__4014 (
            .O(N__25655),
            .I(N__25590));
    InMux I__4013 (
            .O(N__25654),
            .I(N__25590));
    InMux I__4012 (
            .O(N__25653),
            .I(N__25587));
    InMux I__4011 (
            .O(N__25650),
            .I(N__25582));
    InMux I__4010 (
            .O(N__25649),
            .I(N__25582));
    InMux I__4009 (
            .O(N__25646),
            .I(N__25579));
    InMux I__4008 (
            .O(N__25645),
            .I(N__25564));
    InMux I__4007 (
            .O(N__25642),
            .I(N__25564));
    InMux I__4006 (
            .O(N__25639),
            .I(N__25564));
    InMux I__4005 (
            .O(N__25636),
            .I(N__25564));
    InMux I__4004 (
            .O(N__25635),
            .I(N__25564));
    InMux I__4003 (
            .O(N__25634),
            .I(N__25564));
    InMux I__4002 (
            .O(N__25633),
            .I(N__25564));
    InMux I__4001 (
            .O(N__25632),
            .I(N__25561));
    InMux I__4000 (
            .O(N__25629),
            .I(N__25548));
    InMux I__3999 (
            .O(N__25626),
            .I(N__25548));
    InMux I__3998 (
            .O(N__25623),
            .I(N__25548));
    InMux I__3997 (
            .O(N__25620),
            .I(N__25548));
    InMux I__3996 (
            .O(N__25619),
            .I(N__25548));
    InMux I__3995 (
            .O(N__25618),
            .I(N__25548));
    InMux I__3994 (
            .O(N__25615),
            .I(N__25543));
    InMux I__3993 (
            .O(N__25614),
            .I(N__25543));
    InMux I__3992 (
            .O(N__25613),
            .I(N__25528));
    InMux I__3991 (
            .O(N__25610),
            .I(N__25528));
    InMux I__3990 (
            .O(N__25607),
            .I(N__25528));
    InMux I__3989 (
            .O(N__25604),
            .I(N__25528));
    InMux I__3988 (
            .O(N__25603),
            .I(N__25528));
    InMux I__3987 (
            .O(N__25602),
            .I(N__25528));
    InMux I__3986 (
            .O(N__25601),
            .I(N__25528));
    Span4Mux_v I__3985 (
            .O(N__25598),
            .I(N__25525));
    LocalMux I__3984 (
            .O(N__25595),
            .I(N__25518));
    LocalMux I__3983 (
            .O(N__25590),
            .I(N__25518));
    LocalMux I__3982 (
            .O(N__25587),
            .I(N__25518));
    LocalMux I__3981 (
            .O(N__25582),
            .I(N__25513));
    LocalMux I__3980 (
            .O(N__25579),
            .I(N__25513));
    LocalMux I__3979 (
            .O(N__25564),
            .I(N__25508));
    LocalMux I__3978 (
            .O(N__25561),
            .I(N__25508));
    LocalMux I__3977 (
            .O(N__25548),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__3976 (
            .O(N__25543),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__3975 (
            .O(N__25528),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__3974 (
            .O(N__25525),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv12 I__3973 (
            .O(N__25518),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv12 I__3972 (
            .O(N__25513),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__3971 (
            .O(N__25508),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    InMux I__3970 (
            .O(N__25493),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_30 ));
    InMux I__3969 (
            .O(N__25490),
            .I(N__25487));
    LocalMux I__3968 (
            .O(N__25487),
            .I(N__25484));
    Odrv4 I__3967 (
            .O(N__25484),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ));
    InMux I__3966 (
            .O(N__25481),
            .I(N__25478));
    LocalMux I__3965 (
            .O(N__25478),
            .I(\current_shift_inst.un38_control_input_0_cry_1_c_RNOZ0 ));
    InMux I__3964 (
            .O(N__25475),
            .I(N__25472));
    LocalMux I__3963 (
            .O(N__25472),
            .I(\current_shift_inst.N_1717_i ));
    CascadeMux I__3962 (
            .O(N__25469),
            .I(N__25466));
    InMux I__3961 (
            .O(N__25466),
            .I(N__25463));
    LocalMux I__3960 (
            .O(N__25463),
            .I(N__25457));
    InMux I__3959 (
            .O(N__25462),
            .I(N__25454));
    InMux I__3958 (
            .O(N__25461),
            .I(N__25449));
    InMux I__3957 (
            .O(N__25460),
            .I(N__25449));
    Odrv12 I__3956 (
            .O(N__25457),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    LocalMux I__3955 (
            .O(N__25454),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    LocalMux I__3954 (
            .O(N__25449),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    InMux I__3953 (
            .O(N__25442),
            .I(N__25438));
    CascadeMux I__3952 (
            .O(N__25441),
            .I(N__25435));
    LocalMux I__3951 (
            .O(N__25438),
            .I(N__25432));
    InMux I__3950 (
            .O(N__25435),
            .I(N__25429));
    Span4Mux_h I__3949 (
            .O(N__25432),
            .I(N__25426));
    LocalMux I__3948 (
            .O(N__25429),
            .I(N__25423));
    Span4Mux_v I__3947 (
            .O(N__25426),
            .I(N__25420));
    Span4Mux_h I__3946 (
            .O(N__25423),
            .I(N__25417));
    Odrv4 I__3945 (
            .O(N__25420),
            .I(\current_shift_inst.control_inputZ0Z_20 ));
    Odrv4 I__3944 (
            .O(N__25417),
            .I(\current_shift_inst.control_inputZ0Z_20 ));
    InMux I__3943 (
            .O(N__25412),
            .I(N__25409));
    LocalMux I__3942 (
            .O(N__25409),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ));
    InMux I__3941 (
            .O(N__25406),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ));
    CascadeMux I__3940 (
            .O(N__25403),
            .I(N__25400));
    InMux I__3939 (
            .O(N__25400),
            .I(N__25397));
    LocalMux I__3938 (
            .O(N__25397),
            .I(N__25393));
    InMux I__3937 (
            .O(N__25396),
            .I(N__25390));
    Span4Mux_v I__3936 (
            .O(N__25393),
            .I(N__25387));
    LocalMux I__3935 (
            .O(N__25390),
            .I(N__25382));
    Span4Mux_h I__3934 (
            .O(N__25387),
            .I(N__25379));
    InMux I__3933 (
            .O(N__25386),
            .I(N__25376));
    InMux I__3932 (
            .O(N__25385),
            .I(N__25373));
    Span4Mux_v I__3931 (
            .O(N__25382),
            .I(N__25370));
    Odrv4 I__3930 (
            .O(N__25379),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    LocalMux I__3929 (
            .O(N__25376),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    LocalMux I__3928 (
            .O(N__25373),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    Odrv4 I__3927 (
            .O(N__25370),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    InMux I__3926 (
            .O(N__25361),
            .I(N__25357));
    CascadeMux I__3925 (
            .O(N__25360),
            .I(N__25354));
    LocalMux I__3924 (
            .O(N__25357),
            .I(N__25351));
    InMux I__3923 (
            .O(N__25354),
            .I(N__25348));
    Span4Mux_v I__3922 (
            .O(N__25351),
            .I(N__25345));
    LocalMux I__3921 (
            .O(N__25348),
            .I(N__25342));
    Sp12to4 I__3920 (
            .O(N__25345),
            .I(N__25339));
    Span4Mux_h I__3919 (
            .O(N__25342),
            .I(N__25336));
    Odrv12 I__3918 (
            .O(N__25339),
            .I(\current_shift_inst.control_inputZ0Z_21 ));
    Odrv4 I__3917 (
            .O(N__25336),
            .I(\current_shift_inst.control_inputZ0Z_21 ));
    InMux I__3916 (
            .O(N__25331),
            .I(N__25328));
    LocalMux I__3915 (
            .O(N__25328),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ));
    InMux I__3914 (
            .O(N__25325),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ));
    InMux I__3913 (
            .O(N__25322),
            .I(N__25317));
    CascadeMux I__3912 (
            .O(N__25321),
            .I(N__25313));
    CascadeMux I__3911 (
            .O(N__25320),
            .I(N__25310));
    LocalMux I__3910 (
            .O(N__25317),
            .I(N__25307));
    InMux I__3909 (
            .O(N__25316),
            .I(N__25304));
    InMux I__3908 (
            .O(N__25313),
            .I(N__25299));
    InMux I__3907 (
            .O(N__25310),
            .I(N__25299));
    Odrv12 I__3906 (
            .O(N__25307),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    LocalMux I__3905 (
            .O(N__25304),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    LocalMux I__3904 (
            .O(N__25299),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    CascadeMux I__3903 (
            .O(N__25292),
            .I(N__25289));
    InMux I__3902 (
            .O(N__25289),
            .I(N__25285));
    InMux I__3901 (
            .O(N__25288),
            .I(N__25282));
    LocalMux I__3900 (
            .O(N__25285),
            .I(N__25279));
    LocalMux I__3899 (
            .O(N__25282),
            .I(N__25274));
    Span4Mux_h I__3898 (
            .O(N__25279),
            .I(N__25274));
    Span4Mux_v I__3897 (
            .O(N__25274),
            .I(N__25271));
    Odrv4 I__3896 (
            .O(N__25271),
            .I(\current_shift_inst.control_inputZ0Z_22 ));
    InMux I__3895 (
            .O(N__25268),
            .I(N__25265));
    LocalMux I__3894 (
            .O(N__25265),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ));
    InMux I__3893 (
            .O(N__25262),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ));
    InMux I__3892 (
            .O(N__25259),
            .I(N__25254));
    InMux I__3891 (
            .O(N__25258),
            .I(N__25251));
    InMux I__3890 (
            .O(N__25257),
            .I(N__25247));
    LocalMux I__3889 (
            .O(N__25254),
            .I(N__25244));
    LocalMux I__3888 (
            .O(N__25251),
            .I(N__25241));
    InMux I__3887 (
            .O(N__25250),
            .I(N__25238));
    LocalMux I__3886 (
            .O(N__25247),
            .I(N__25235));
    Odrv12 I__3885 (
            .O(N__25244),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    Odrv4 I__3884 (
            .O(N__25241),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    LocalMux I__3883 (
            .O(N__25238),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    Odrv4 I__3882 (
            .O(N__25235),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    CascadeMux I__3881 (
            .O(N__25226),
            .I(N__25223));
    InMux I__3880 (
            .O(N__25223),
            .I(N__25219));
    InMux I__3879 (
            .O(N__25222),
            .I(N__25216));
    LocalMux I__3878 (
            .O(N__25219),
            .I(N__25213));
    LocalMux I__3877 (
            .O(N__25216),
            .I(N__25208));
    Span4Mux_h I__3876 (
            .O(N__25213),
            .I(N__25208));
    Span4Mux_v I__3875 (
            .O(N__25208),
            .I(N__25205));
    Odrv4 I__3874 (
            .O(N__25205),
            .I(\current_shift_inst.control_inputZ0Z_23 ));
    CascadeMux I__3873 (
            .O(N__25202),
            .I(N__25199));
    InMux I__3872 (
            .O(N__25199),
            .I(N__25196));
    LocalMux I__3871 (
            .O(N__25196),
            .I(N__25193));
    Span4Mux_h I__3870 (
            .O(N__25193),
            .I(N__25190));
    Odrv4 I__3869 (
            .O(N__25190),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ));
    InMux I__3868 (
            .O(N__25187),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ));
    CascadeMux I__3867 (
            .O(N__25184),
            .I(N__25181));
    InMux I__3866 (
            .O(N__25181),
            .I(N__25177));
    InMux I__3865 (
            .O(N__25180),
            .I(N__25173));
    LocalMux I__3864 (
            .O(N__25177),
            .I(N__25170));
    InMux I__3863 (
            .O(N__25176),
            .I(N__25167));
    LocalMux I__3862 (
            .O(N__25173),
            .I(N__25163));
    Span4Mux_h I__3861 (
            .O(N__25170),
            .I(N__25158));
    LocalMux I__3860 (
            .O(N__25167),
            .I(N__25158));
    InMux I__3859 (
            .O(N__25166),
            .I(N__25155));
    Span4Mux_h I__3858 (
            .O(N__25163),
            .I(N__25152));
    Odrv4 I__3857 (
            .O(N__25158),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    LocalMux I__3856 (
            .O(N__25155),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv4 I__3855 (
            .O(N__25152),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    CascadeMux I__3854 (
            .O(N__25145),
            .I(N__25141));
    InMux I__3853 (
            .O(N__25144),
            .I(N__25138));
    InMux I__3852 (
            .O(N__25141),
            .I(N__25135));
    LocalMux I__3851 (
            .O(N__25138),
            .I(N__25132));
    LocalMux I__3850 (
            .O(N__25135),
            .I(N__25129));
    Span4Mux_h I__3849 (
            .O(N__25132),
            .I(N__25126));
    Span4Mux_h I__3848 (
            .O(N__25129),
            .I(N__25123));
    Odrv4 I__3847 (
            .O(N__25126),
            .I(\current_shift_inst.control_inputZ0Z_24 ));
    Odrv4 I__3846 (
            .O(N__25123),
            .I(\current_shift_inst.control_inputZ0Z_24 ));
    InMux I__3845 (
            .O(N__25118),
            .I(N__25115));
    LocalMux I__3844 (
            .O(N__25115),
            .I(N__25112));
    Odrv12 I__3843 (
            .O(N__25112),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ));
    InMux I__3842 (
            .O(N__25109),
            .I(bfn_9_16_0_));
    InMux I__3841 (
            .O(N__25106),
            .I(N__25102));
    InMux I__3840 (
            .O(N__25105),
            .I(N__25098));
    LocalMux I__3839 (
            .O(N__25102),
            .I(N__25095));
    InMux I__3838 (
            .O(N__25101),
            .I(N__25092));
    LocalMux I__3837 (
            .O(N__25098),
            .I(N__25088));
    Span4Mux_h I__3836 (
            .O(N__25095),
            .I(N__25083));
    LocalMux I__3835 (
            .O(N__25092),
            .I(N__25083));
    InMux I__3834 (
            .O(N__25091),
            .I(N__25080));
    Span4Mux_h I__3833 (
            .O(N__25088),
            .I(N__25077));
    Odrv4 I__3832 (
            .O(N__25083),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    LocalMux I__3831 (
            .O(N__25080),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    Odrv4 I__3830 (
            .O(N__25077),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    InMux I__3829 (
            .O(N__25070),
            .I(N__25067));
    LocalMux I__3828 (
            .O(N__25067),
            .I(N__25064));
    Span4Mux_h I__3827 (
            .O(N__25064),
            .I(N__25061));
    Odrv4 I__3826 (
            .O(N__25061),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ));
    InMux I__3825 (
            .O(N__25058),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ));
    CascadeMux I__3824 (
            .O(N__25055),
            .I(N__25051));
    CascadeMux I__3823 (
            .O(N__25054),
            .I(N__25047));
    InMux I__3822 (
            .O(N__25051),
            .I(N__25044));
    CascadeMux I__3821 (
            .O(N__25050),
            .I(N__25041));
    InMux I__3820 (
            .O(N__25047),
            .I(N__25037));
    LocalMux I__3819 (
            .O(N__25044),
            .I(N__25034));
    InMux I__3818 (
            .O(N__25041),
            .I(N__25031));
    CascadeMux I__3817 (
            .O(N__25040),
            .I(N__25028));
    LocalMux I__3816 (
            .O(N__25037),
            .I(N__25025));
    Span4Mux_h I__3815 (
            .O(N__25034),
            .I(N__25020));
    LocalMux I__3814 (
            .O(N__25031),
            .I(N__25020));
    InMux I__3813 (
            .O(N__25028),
            .I(N__25017));
    Span4Mux_h I__3812 (
            .O(N__25025),
            .I(N__25014));
    Odrv4 I__3811 (
            .O(N__25020),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    LocalMux I__3810 (
            .O(N__25017),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv4 I__3809 (
            .O(N__25014),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    InMux I__3808 (
            .O(N__25007),
            .I(N__25004));
    LocalMux I__3807 (
            .O(N__25004),
            .I(N__25001));
    Span4Mux_h I__3806 (
            .O(N__25001),
            .I(N__24998));
    Odrv4 I__3805 (
            .O(N__24998),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ));
    InMux I__3804 (
            .O(N__24995),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ));
    InMux I__3803 (
            .O(N__24992),
            .I(N__24989));
    LocalMux I__3802 (
            .O(N__24989),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ));
    InMux I__3801 (
            .O(N__24986),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ));
    CascadeMux I__3800 (
            .O(N__24983),
            .I(N__24979));
    InMux I__3799 (
            .O(N__24982),
            .I(N__24976));
    InMux I__3798 (
            .O(N__24979),
            .I(N__24973));
    LocalMux I__3797 (
            .O(N__24976),
            .I(N__24968));
    LocalMux I__3796 (
            .O(N__24973),
            .I(N__24965));
    InMux I__3795 (
            .O(N__24972),
            .I(N__24962));
    InMux I__3794 (
            .O(N__24971),
            .I(N__24959));
    Span4Mux_h I__3793 (
            .O(N__24968),
            .I(N__24956));
    Odrv12 I__3792 (
            .O(N__24965),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    LocalMux I__3791 (
            .O(N__24962),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    LocalMux I__3790 (
            .O(N__24959),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    Odrv4 I__3789 (
            .O(N__24956),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    CascadeMux I__3788 (
            .O(N__24947),
            .I(N__24943));
    InMux I__3787 (
            .O(N__24946),
            .I(N__24940));
    InMux I__3786 (
            .O(N__24943),
            .I(N__24937));
    LocalMux I__3785 (
            .O(N__24940),
            .I(N__24934));
    LocalMux I__3784 (
            .O(N__24937),
            .I(N__24931));
    Span4Mux_h I__3783 (
            .O(N__24934),
            .I(N__24926));
    Span4Mux_h I__3782 (
            .O(N__24931),
            .I(N__24926));
    Odrv4 I__3781 (
            .O(N__24926),
            .I(\current_shift_inst.control_inputZ0Z_13 ));
    InMux I__3780 (
            .O(N__24923),
            .I(N__24920));
    LocalMux I__3779 (
            .O(N__24920),
            .I(N__24917));
    Odrv4 I__3778 (
            .O(N__24917),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ));
    InMux I__3777 (
            .O(N__24914),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ));
    InMux I__3776 (
            .O(N__24911),
            .I(N__24907));
    InMux I__3775 (
            .O(N__24910),
            .I(N__24904));
    LocalMux I__3774 (
            .O(N__24907),
            .I(N__24901));
    LocalMux I__3773 (
            .O(N__24904),
            .I(N__24898));
    Span12Mux_v I__3772 (
            .O(N__24901),
            .I(N__24895));
    Span12Mux_v I__3771 (
            .O(N__24898),
            .I(N__24892));
    Odrv12 I__3770 (
            .O(N__24895),
            .I(\current_shift_inst.control_inputZ0Z_14 ));
    Odrv12 I__3769 (
            .O(N__24892),
            .I(\current_shift_inst.control_inputZ0Z_14 ));
    CascadeMux I__3768 (
            .O(N__24887),
            .I(N__24884));
    InMux I__3767 (
            .O(N__24884),
            .I(N__24881));
    LocalMux I__3766 (
            .O(N__24881),
            .I(N__24876));
    InMux I__3765 (
            .O(N__24880),
            .I(N__24872));
    CascadeMux I__3764 (
            .O(N__24879),
            .I(N__24869));
    Span4Mux_v I__3763 (
            .O(N__24876),
            .I(N__24866));
    InMux I__3762 (
            .O(N__24875),
            .I(N__24863));
    LocalMux I__3761 (
            .O(N__24872),
            .I(N__24860));
    InMux I__3760 (
            .O(N__24869),
            .I(N__24857));
    Span4Mux_h I__3759 (
            .O(N__24866),
            .I(N__24852));
    LocalMux I__3758 (
            .O(N__24863),
            .I(N__24852));
    Odrv4 I__3757 (
            .O(N__24860),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    LocalMux I__3756 (
            .O(N__24857),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    Odrv4 I__3755 (
            .O(N__24852),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    InMux I__3754 (
            .O(N__24845),
            .I(N__24842));
    LocalMux I__3753 (
            .O(N__24842),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ));
    InMux I__3752 (
            .O(N__24839),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ));
    CascadeMux I__3751 (
            .O(N__24836),
            .I(N__24833));
    InMux I__3750 (
            .O(N__24833),
            .I(N__24829));
    InMux I__3749 (
            .O(N__24832),
            .I(N__24826));
    LocalMux I__3748 (
            .O(N__24829),
            .I(N__24822));
    LocalMux I__3747 (
            .O(N__24826),
            .I(N__24818));
    InMux I__3746 (
            .O(N__24825),
            .I(N__24815));
    Span4Mux_h I__3745 (
            .O(N__24822),
            .I(N__24812));
    InMux I__3744 (
            .O(N__24821),
            .I(N__24809));
    Span4Mux_v I__3743 (
            .O(N__24818),
            .I(N__24804));
    LocalMux I__3742 (
            .O(N__24815),
            .I(N__24804));
    Odrv4 I__3741 (
            .O(N__24812),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    LocalMux I__3740 (
            .O(N__24809),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    Odrv4 I__3739 (
            .O(N__24804),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    InMux I__3738 (
            .O(N__24797),
            .I(N__24793));
    CascadeMux I__3737 (
            .O(N__24796),
            .I(N__24790));
    LocalMux I__3736 (
            .O(N__24793),
            .I(N__24787));
    InMux I__3735 (
            .O(N__24790),
            .I(N__24784));
    Span4Mux_h I__3734 (
            .O(N__24787),
            .I(N__24779));
    LocalMux I__3733 (
            .O(N__24784),
            .I(N__24779));
    Span4Mux_h I__3732 (
            .O(N__24779),
            .I(N__24776));
    Span4Mux_v I__3731 (
            .O(N__24776),
            .I(N__24773));
    Odrv4 I__3730 (
            .O(N__24773),
            .I(\current_shift_inst.control_inputZ0Z_15 ));
    InMux I__3729 (
            .O(N__24770),
            .I(N__24767));
    LocalMux I__3728 (
            .O(N__24767),
            .I(N__24764));
    Span4Mux_h I__3727 (
            .O(N__24764),
            .I(N__24761));
    Odrv4 I__3726 (
            .O(N__24761),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ));
    InMux I__3725 (
            .O(N__24758),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ));
    CascadeMux I__3724 (
            .O(N__24755),
            .I(N__24750));
    InMux I__3723 (
            .O(N__24754),
            .I(N__24747));
    CascadeMux I__3722 (
            .O(N__24753),
            .I(N__24743));
    InMux I__3721 (
            .O(N__24750),
            .I(N__24740));
    LocalMux I__3720 (
            .O(N__24747),
            .I(N__24737));
    InMux I__3719 (
            .O(N__24746),
            .I(N__24734));
    InMux I__3718 (
            .O(N__24743),
            .I(N__24731));
    LocalMux I__3717 (
            .O(N__24740),
            .I(N__24728));
    Odrv12 I__3716 (
            .O(N__24737),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    LocalMux I__3715 (
            .O(N__24734),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    LocalMux I__3714 (
            .O(N__24731),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    Odrv4 I__3713 (
            .O(N__24728),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    CascadeMux I__3712 (
            .O(N__24719),
            .I(N__24715));
    InMux I__3711 (
            .O(N__24718),
            .I(N__24712));
    InMux I__3710 (
            .O(N__24715),
            .I(N__24709));
    LocalMux I__3709 (
            .O(N__24712),
            .I(N__24706));
    LocalMux I__3708 (
            .O(N__24709),
            .I(N__24703));
    Span4Mux_h I__3707 (
            .O(N__24706),
            .I(N__24700));
    Span4Mux_h I__3706 (
            .O(N__24703),
            .I(N__24697));
    Odrv4 I__3705 (
            .O(N__24700),
            .I(\current_shift_inst.control_inputZ0Z_16 ));
    Odrv4 I__3704 (
            .O(N__24697),
            .I(\current_shift_inst.control_inputZ0Z_16 ));
    InMux I__3703 (
            .O(N__24692),
            .I(N__24689));
    LocalMux I__3702 (
            .O(N__24689),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ));
    InMux I__3701 (
            .O(N__24686),
            .I(bfn_9_15_0_));
    InMux I__3700 (
            .O(N__24683),
            .I(N__24680));
    LocalMux I__3699 (
            .O(N__24680),
            .I(N__24674));
    InMux I__3698 (
            .O(N__24679),
            .I(N__24671));
    InMux I__3697 (
            .O(N__24678),
            .I(N__24666));
    InMux I__3696 (
            .O(N__24677),
            .I(N__24666));
    Odrv12 I__3695 (
            .O(N__24674),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    LocalMux I__3694 (
            .O(N__24671),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    LocalMux I__3693 (
            .O(N__24666),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    InMux I__3692 (
            .O(N__24659),
            .I(N__24655));
    CascadeMux I__3691 (
            .O(N__24658),
            .I(N__24652));
    LocalMux I__3690 (
            .O(N__24655),
            .I(N__24649));
    InMux I__3689 (
            .O(N__24652),
            .I(N__24646));
    Span4Mux_h I__3688 (
            .O(N__24649),
            .I(N__24643));
    LocalMux I__3687 (
            .O(N__24646),
            .I(N__24640));
    Span4Mux_v I__3686 (
            .O(N__24643),
            .I(N__24637));
    Span4Mux_h I__3685 (
            .O(N__24640),
            .I(N__24634));
    Odrv4 I__3684 (
            .O(N__24637),
            .I(\current_shift_inst.control_inputZ0Z_17 ));
    Odrv4 I__3683 (
            .O(N__24634),
            .I(\current_shift_inst.control_inputZ0Z_17 ));
    InMux I__3682 (
            .O(N__24629),
            .I(N__24626));
    LocalMux I__3681 (
            .O(N__24626),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ));
    InMux I__3680 (
            .O(N__24623),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ));
    CascadeMux I__3679 (
            .O(N__24620),
            .I(N__24617));
    InMux I__3678 (
            .O(N__24617),
            .I(N__24614));
    LocalMux I__3677 (
            .O(N__24614),
            .I(N__24607));
    InMux I__3676 (
            .O(N__24613),
            .I(N__24600));
    InMux I__3675 (
            .O(N__24612),
            .I(N__24600));
    InMux I__3674 (
            .O(N__24611),
            .I(N__24600));
    InMux I__3673 (
            .O(N__24610),
            .I(N__24596));
    Span4Mux_h I__3672 (
            .O(N__24607),
            .I(N__24593));
    LocalMux I__3671 (
            .O(N__24600),
            .I(N__24590));
    InMux I__3670 (
            .O(N__24599),
            .I(N__24587));
    LocalMux I__3669 (
            .O(N__24596),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    Odrv4 I__3668 (
            .O(N__24593),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    Odrv4 I__3667 (
            .O(N__24590),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    LocalMux I__3666 (
            .O(N__24587),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    CascadeMux I__3665 (
            .O(N__24578),
            .I(N__24574));
    InMux I__3664 (
            .O(N__24577),
            .I(N__24571));
    InMux I__3663 (
            .O(N__24574),
            .I(N__24568));
    LocalMux I__3662 (
            .O(N__24571),
            .I(N__24565));
    LocalMux I__3661 (
            .O(N__24568),
            .I(N__24562));
    Span4Mux_h I__3660 (
            .O(N__24565),
            .I(N__24559));
    Span4Mux_h I__3659 (
            .O(N__24562),
            .I(N__24556));
    Odrv4 I__3658 (
            .O(N__24559),
            .I(\current_shift_inst.control_inputZ0Z_18 ));
    Odrv4 I__3657 (
            .O(N__24556),
            .I(\current_shift_inst.control_inputZ0Z_18 ));
    InMux I__3656 (
            .O(N__24551),
            .I(N__24548));
    LocalMux I__3655 (
            .O(N__24548),
            .I(N__24545));
    Odrv4 I__3654 (
            .O(N__24545),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ));
    InMux I__3653 (
            .O(N__24542),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ));
    InMux I__3652 (
            .O(N__24539),
            .I(N__24536));
    LocalMux I__3651 (
            .O(N__24536),
            .I(N__24530));
    InMux I__3650 (
            .O(N__24535),
            .I(N__24527));
    InMux I__3649 (
            .O(N__24534),
            .I(N__24522));
    InMux I__3648 (
            .O(N__24533),
            .I(N__24522));
    Odrv12 I__3647 (
            .O(N__24530),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    LocalMux I__3646 (
            .O(N__24527),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    LocalMux I__3645 (
            .O(N__24522),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    InMux I__3644 (
            .O(N__24515),
            .I(N__24511));
    CascadeMux I__3643 (
            .O(N__24514),
            .I(N__24508));
    LocalMux I__3642 (
            .O(N__24511),
            .I(N__24505));
    InMux I__3641 (
            .O(N__24508),
            .I(N__24502));
    Span4Mux_h I__3640 (
            .O(N__24505),
            .I(N__24499));
    LocalMux I__3639 (
            .O(N__24502),
            .I(N__24496));
    Span4Mux_v I__3638 (
            .O(N__24499),
            .I(N__24493));
    Span4Mux_h I__3637 (
            .O(N__24496),
            .I(N__24490));
    Odrv4 I__3636 (
            .O(N__24493),
            .I(\current_shift_inst.control_inputZ0Z_19 ));
    Odrv4 I__3635 (
            .O(N__24490),
            .I(\current_shift_inst.control_inputZ0Z_19 ));
    InMux I__3634 (
            .O(N__24485),
            .I(N__24482));
    LocalMux I__3633 (
            .O(N__24482),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ));
    InMux I__3632 (
            .O(N__24479),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ));
    InMux I__3631 (
            .O(N__24476),
            .I(N__24473));
    LocalMux I__3630 (
            .O(N__24473),
            .I(N__24469));
    InMux I__3629 (
            .O(N__24472),
            .I(N__24466));
    Span4Mux_h I__3628 (
            .O(N__24469),
            .I(N__24460));
    LocalMux I__3627 (
            .O(N__24466),
            .I(N__24460));
    CascadeMux I__3626 (
            .O(N__24465),
            .I(N__24456));
    Span4Mux_h I__3625 (
            .O(N__24460),
            .I(N__24453));
    InMux I__3624 (
            .O(N__24459),
            .I(N__24448));
    InMux I__3623 (
            .O(N__24456),
            .I(N__24448));
    Odrv4 I__3622 (
            .O(N__24453),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    LocalMux I__3621 (
            .O(N__24448),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    InMux I__3620 (
            .O(N__24443),
            .I(N__24439));
    CascadeMux I__3619 (
            .O(N__24442),
            .I(N__24436));
    LocalMux I__3618 (
            .O(N__24439),
            .I(N__24433));
    InMux I__3617 (
            .O(N__24436),
            .I(N__24430));
    Span4Mux_h I__3616 (
            .O(N__24433),
            .I(N__24427));
    LocalMux I__3615 (
            .O(N__24430),
            .I(N__24424));
    Span4Mux_v I__3614 (
            .O(N__24427),
            .I(N__24421));
    Span4Mux_h I__3613 (
            .O(N__24424),
            .I(N__24418));
    Odrv4 I__3612 (
            .O(N__24421),
            .I(\current_shift_inst.control_inputZ0Z_5 ));
    Odrv4 I__3611 (
            .O(N__24418),
            .I(\current_shift_inst.control_inputZ0Z_5 ));
    InMux I__3610 (
            .O(N__24413),
            .I(N__24410));
    LocalMux I__3609 (
            .O(N__24410),
            .I(N__24407));
    Span4Mux_h I__3608 (
            .O(N__24407),
            .I(N__24404));
    Odrv4 I__3607 (
            .O(N__24404),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ));
    InMux I__3606 (
            .O(N__24401),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ));
    InMux I__3605 (
            .O(N__24398),
            .I(N__24395));
    LocalMux I__3604 (
            .O(N__24395),
            .I(N__24391));
    InMux I__3603 (
            .O(N__24394),
            .I(N__24388));
    Span4Mux_h I__3602 (
            .O(N__24391),
            .I(N__24381));
    LocalMux I__3601 (
            .O(N__24388),
            .I(N__24381));
    InMux I__3600 (
            .O(N__24387),
            .I(N__24376));
    InMux I__3599 (
            .O(N__24386),
            .I(N__24376));
    Span4Mux_h I__3598 (
            .O(N__24381),
            .I(N__24373));
    LocalMux I__3597 (
            .O(N__24376),
            .I(N__24370));
    Odrv4 I__3596 (
            .O(N__24373),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    Odrv4 I__3595 (
            .O(N__24370),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    CascadeMux I__3594 (
            .O(N__24365),
            .I(N__24361));
    InMux I__3593 (
            .O(N__24364),
            .I(N__24358));
    InMux I__3592 (
            .O(N__24361),
            .I(N__24355));
    LocalMux I__3591 (
            .O(N__24358),
            .I(N__24352));
    LocalMux I__3590 (
            .O(N__24355),
            .I(N__24349));
    Span4Mux_h I__3589 (
            .O(N__24352),
            .I(N__24344));
    Span4Mux_h I__3588 (
            .O(N__24349),
            .I(N__24344));
    Span4Mux_v I__3587 (
            .O(N__24344),
            .I(N__24341));
    Odrv4 I__3586 (
            .O(N__24341),
            .I(\current_shift_inst.control_inputZ0Z_6 ));
    InMux I__3585 (
            .O(N__24338),
            .I(N__24335));
    LocalMux I__3584 (
            .O(N__24335),
            .I(N__24332));
    Span4Mux_h I__3583 (
            .O(N__24332),
            .I(N__24329));
    Odrv4 I__3582 (
            .O(N__24329),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ));
    InMux I__3581 (
            .O(N__24326),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ));
    InMux I__3580 (
            .O(N__24323),
            .I(N__24320));
    LocalMux I__3579 (
            .O(N__24320),
            .I(N__24317));
    Span4Mux_h I__3578 (
            .O(N__24317),
            .I(N__24313));
    InMux I__3577 (
            .O(N__24316),
            .I(N__24310));
    Span4Mux_v I__3576 (
            .O(N__24313),
            .I(N__24307));
    LocalMux I__3575 (
            .O(N__24310),
            .I(\current_shift_inst.control_inputZ0Z_7 ));
    Odrv4 I__3574 (
            .O(N__24307),
            .I(\current_shift_inst.control_inputZ0Z_7 ));
    InMux I__3573 (
            .O(N__24302),
            .I(N__24299));
    LocalMux I__3572 (
            .O(N__24299),
            .I(N__24295));
    CascadeMux I__3571 (
            .O(N__24298),
            .I(N__24292));
    Span4Mux_h I__3570 (
            .O(N__24295),
            .I(N__24287));
    InMux I__3569 (
            .O(N__24292),
            .I(N__24284));
    InMux I__3568 (
            .O(N__24291),
            .I(N__24279));
    InMux I__3567 (
            .O(N__24290),
            .I(N__24279));
    Odrv4 I__3566 (
            .O(N__24287),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    LocalMux I__3565 (
            .O(N__24284),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    LocalMux I__3564 (
            .O(N__24279),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    InMux I__3563 (
            .O(N__24272),
            .I(N__24269));
    LocalMux I__3562 (
            .O(N__24269),
            .I(N__24266));
    Odrv4 I__3561 (
            .O(N__24266),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ));
    InMux I__3560 (
            .O(N__24263),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ));
    InMux I__3559 (
            .O(N__24260),
            .I(N__24257));
    LocalMux I__3558 (
            .O(N__24257),
            .I(N__24251));
    InMux I__3557 (
            .O(N__24256),
            .I(N__24248));
    InMux I__3556 (
            .O(N__24255),
            .I(N__24243));
    InMux I__3555 (
            .O(N__24254),
            .I(N__24243));
    Odrv12 I__3554 (
            .O(N__24251),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    LocalMux I__3553 (
            .O(N__24248),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    LocalMux I__3552 (
            .O(N__24243),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    InMux I__3551 (
            .O(N__24236),
            .I(N__24232));
    CascadeMux I__3550 (
            .O(N__24235),
            .I(N__24229));
    LocalMux I__3549 (
            .O(N__24232),
            .I(N__24226));
    InMux I__3548 (
            .O(N__24229),
            .I(N__24223));
    Span4Mux_v I__3547 (
            .O(N__24226),
            .I(N__24220));
    LocalMux I__3546 (
            .O(N__24223),
            .I(N__24217));
    Span4Mux_v I__3545 (
            .O(N__24220),
            .I(N__24214));
    Span4Mux_h I__3544 (
            .O(N__24217),
            .I(N__24211));
    Odrv4 I__3543 (
            .O(N__24214),
            .I(\current_shift_inst.control_inputZ0Z_8 ));
    Odrv4 I__3542 (
            .O(N__24211),
            .I(\current_shift_inst.control_inputZ0Z_8 ));
    InMux I__3541 (
            .O(N__24206),
            .I(N__24203));
    LocalMux I__3540 (
            .O(N__24203),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ));
    InMux I__3539 (
            .O(N__24200),
            .I(bfn_9_14_0_));
    InMux I__3538 (
            .O(N__24197),
            .I(N__24194));
    LocalMux I__3537 (
            .O(N__24194),
            .I(N__24191));
    Span4Mux_h I__3536 (
            .O(N__24191),
            .I(N__24185));
    InMux I__3535 (
            .O(N__24190),
            .I(N__24180));
    InMux I__3534 (
            .O(N__24189),
            .I(N__24180));
    InMux I__3533 (
            .O(N__24188),
            .I(N__24177));
    Odrv4 I__3532 (
            .O(N__24185),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    LocalMux I__3531 (
            .O(N__24180),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    LocalMux I__3530 (
            .O(N__24177),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    InMux I__3529 (
            .O(N__24170),
            .I(N__24166));
    CascadeMux I__3528 (
            .O(N__24169),
            .I(N__24163));
    LocalMux I__3527 (
            .O(N__24166),
            .I(N__24160));
    InMux I__3526 (
            .O(N__24163),
            .I(N__24157));
    Span4Mux_h I__3525 (
            .O(N__24160),
            .I(N__24154));
    LocalMux I__3524 (
            .O(N__24157),
            .I(N__24151));
    Span4Mux_v I__3523 (
            .O(N__24154),
            .I(N__24148));
    Span4Mux_h I__3522 (
            .O(N__24151),
            .I(N__24145));
    Odrv4 I__3521 (
            .O(N__24148),
            .I(\current_shift_inst.control_inputZ0Z_9 ));
    Odrv4 I__3520 (
            .O(N__24145),
            .I(\current_shift_inst.control_inputZ0Z_9 ));
    InMux I__3519 (
            .O(N__24140),
            .I(N__24137));
    LocalMux I__3518 (
            .O(N__24137),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ));
    InMux I__3517 (
            .O(N__24134),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ));
    InMux I__3516 (
            .O(N__24131),
            .I(N__24128));
    LocalMux I__3515 (
            .O(N__24128),
            .I(N__24123));
    InMux I__3514 (
            .O(N__24127),
            .I(N__24120));
    InMux I__3513 (
            .O(N__24126),
            .I(N__24116));
    Span4Mux_h I__3512 (
            .O(N__24123),
            .I(N__24111));
    LocalMux I__3511 (
            .O(N__24120),
            .I(N__24111));
    InMux I__3510 (
            .O(N__24119),
            .I(N__24108));
    LocalMux I__3509 (
            .O(N__24116),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    Odrv4 I__3508 (
            .O(N__24111),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    LocalMux I__3507 (
            .O(N__24108),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    CascadeMux I__3506 (
            .O(N__24101),
            .I(N__24097));
    InMux I__3505 (
            .O(N__24100),
            .I(N__24094));
    InMux I__3504 (
            .O(N__24097),
            .I(N__24091));
    LocalMux I__3503 (
            .O(N__24094),
            .I(N__24088));
    LocalMux I__3502 (
            .O(N__24091),
            .I(N__24085));
    Span4Mux_h I__3501 (
            .O(N__24088),
            .I(N__24080));
    Span4Mux_h I__3500 (
            .O(N__24085),
            .I(N__24080));
    Odrv4 I__3499 (
            .O(N__24080),
            .I(\current_shift_inst.control_inputZ0Z_10 ));
    InMux I__3498 (
            .O(N__24077),
            .I(N__24074));
    LocalMux I__3497 (
            .O(N__24074),
            .I(N__24071));
    Odrv12 I__3496 (
            .O(N__24071),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ));
    InMux I__3495 (
            .O(N__24068),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ));
    InMux I__3494 (
            .O(N__24065),
            .I(N__24060));
    CascadeMux I__3493 (
            .O(N__24064),
            .I(N__24057));
    InMux I__3492 (
            .O(N__24063),
            .I(N__24054));
    LocalMux I__3491 (
            .O(N__24060),
            .I(N__24051));
    InMux I__3490 (
            .O(N__24057),
            .I(N__24047));
    LocalMux I__3489 (
            .O(N__24054),
            .I(N__24042));
    Span4Mux_h I__3488 (
            .O(N__24051),
            .I(N__24042));
    InMux I__3487 (
            .O(N__24050),
            .I(N__24039));
    LocalMux I__3486 (
            .O(N__24047),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv4 I__3485 (
            .O(N__24042),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    LocalMux I__3484 (
            .O(N__24039),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    InMux I__3483 (
            .O(N__24032),
            .I(N__24028));
    CascadeMux I__3482 (
            .O(N__24031),
            .I(N__24025));
    LocalMux I__3481 (
            .O(N__24028),
            .I(N__24022));
    InMux I__3480 (
            .O(N__24025),
            .I(N__24019));
    Span4Mux_v I__3479 (
            .O(N__24022),
            .I(N__24016));
    LocalMux I__3478 (
            .O(N__24019),
            .I(N__24013));
    Span4Mux_v I__3477 (
            .O(N__24016),
            .I(N__24010));
    Span4Mux_h I__3476 (
            .O(N__24013),
            .I(N__24007));
    Odrv4 I__3475 (
            .O(N__24010),
            .I(\current_shift_inst.control_inputZ0Z_11 ));
    Odrv4 I__3474 (
            .O(N__24007),
            .I(\current_shift_inst.control_inputZ0Z_11 ));
    InMux I__3473 (
            .O(N__24002),
            .I(N__23999));
    LocalMux I__3472 (
            .O(N__23999),
            .I(N__23996));
    Odrv12 I__3471 (
            .O(N__23996),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ));
    InMux I__3470 (
            .O(N__23993),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ));
    InMux I__3469 (
            .O(N__23990),
            .I(N__23985));
    InMux I__3468 (
            .O(N__23989),
            .I(N__23982));
    InMux I__3467 (
            .O(N__23988),
            .I(N__23978));
    LocalMux I__3466 (
            .O(N__23985),
            .I(N__23975));
    LocalMux I__3465 (
            .O(N__23982),
            .I(N__23972));
    InMux I__3464 (
            .O(N__23981),
            .I(N__23969));
    LocalMux I__3463 (
            .O(N__23978),
            .I(N__23964));
    Span4Mux_h I__3462 (
            .O(N__23975),
            .I(N__23964));
    Odrv12 I__3461 (
            .O(N__23972),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    LocalMux I__3460 (
            .O(N__23969),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    Odrv4 I__3459 (
            .O(N__23964),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    CascadeMux I__3458 (
            .O(N__23957),
            .I(N__23953));
    InMux I__3457 (
            .O(N__23956),
            .I(N__23950));
    InMux I__3456 (
            .O(N__23953),
            .I(N__23947));
    LocalMux I__3455 (
            .O(N__23950),
            .I(N__23944));
    LocalMux I__3454 (
            .O(N__23947),
            .I(N__23941));
    Span4Mux_h I__3453 (
            .O(N__23944),
            .I(N__23938));
    Span4Mux_h I__3452 (
            .O(N__23941),
            .I(N__23935));
    Odrv4 I__3451 (
            .O(N__23938),
            .I(\current_shift_inst.control_inputZ0Z_12 ));
    Odrv4 I__3450 (
            .O(N__23935),
            .I(\current_shift_inst.control_inputZ0Z_12 ));
    CascadeMux I__3449 (
            .O(N__23930),
            .I(N__23927));
    InMux I__3448 (
            .O(N__23927),
            .I(N__23924));
    LocalMux I__3447 (
            .O(N__23924),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ));
    InMux I__3446 (
            .O(N__23921),
            .I(N__23918));
    LocalMux I__3445 (
            .O(N__23918),
            .I(N__23915));
    Odrv4 I__3444 (
            .O(N__23915),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0 ));
    CascadeMux I__3443 (
            .O(N__23912),
            .I(N__23908));
    InMux I__3442 (
            .O(N__23911),
            .I(N__23905));
    InMux I__3441 (
            .O(N__23908),
            .I(N__23902));
    LocalMux I__3440 (
            .O(N__23905),
            .I(N__23899));
    LocalMux I__3439 (
            .O(N__23902),
            .I(N__23896));
    Span4Mux_h I__3438 (
            .O(N__23899),
            .I(N__23891));
    Span4Mux_h I__3437 (
            .O(N__23896),
            .I(N__23891));
    Odrv4 I__3436 (
            .O(N__23891),
            .I(\current_shift_inst.control_inputZ0Z_0 ));
    InMux I__3435 (
            .O(N__23888),
            .I(N__23885));
    LocalMux I__3434 (
            .O(N__23885),
            .I(N__23882));
    Span4Mux_h I__3433 (
            .O(N__23882),
            .I(N__23877));
    InMux I__3432 (
            .O(N__23881),
            .I(N__23874));
    InMux I__3431 (
            .O(N__23880),
            .I(N__23871));
    Odrv4 I__3430 (
            .O(N__23877),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ));
    LocalMux I__3429 (
            .O(N__23874),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ));
    LocalMux I__3428 (
            .O(N__23871),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ));
    InMux I__3427 (
            .O(N__23864),
            .I(N__23860));
    CascadeMux I__3426 (
            .O(N__23863),
            .I(N__23857));
    LocalMux I__3425 (
            .O(N__23860),
            .I(N__23854));
    InMux I__3424 (
            .O(N__23857),
            .I(N__23851));
    Span4Mux_h I__3423 (
            .O(N__23854),
            .I(N__23848));
    LocalMux I__3422 (
            .O(N__23851),
            .I(N__23845));
    Span4Mux_v I__3421 (
            .O(N__23848),
            .I(N__23842));
    Span4Mux_h I__3420 (
            .O(N__23845),
            .I(N__23839));
    Odrv4 I__3419 (
            .O(N__23842),
            .I(\current_shift_inst.control_inputZ0Z_1 ));
    Odrv4 I__3418 (
            .O(N__23839),
            .I(\current_shift_inst.control_inputZ0Z_1 ));
    InMux I__3417 (
            .O(N__23834),
            .I(N__23831));
    LocalMux I__3416 (
            .O(N__23831),
            .I(N__23826));
    InMux I__3415 (
            .O(N__23830),
            .I(N__23823));
    InMux I__3414 (
            .O(N__23829),
            .I(N__23820));
    Span4Mux_h I__3413 (
            .O(N__23826),
            .I(N__23815));
    LocalMux I__3412 (
            .O(N__23823),
            .I(N__23815));
    LocalMux I__3411 (
            .O(N__23820),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv4 I__3410 (
            .O(N__23815),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    InMux I__3409 (
            .O(N__23810),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_0 ));
    CascadeMux I__3408 (
            .O(N__23807),
            .I(N__23803));
    InMux I__3407 (
            .O(N__23806),
            .I(N__23800));
    InMux I__3406 (
            .O(N__23803),
            .I(N__23797));
    LocalMux I__3405 (
            .O(N__23800),
            .I(N__23794));
    LocalMux I__3404 (
            .O(N__23797),
            .I(N__23791));
    Span4Mux_h I__3403 (
            .O(N__23794),
            .I(N__23786));
    Span4Mux_h I__3402 (
            .O(N__23791),
            .I(N__23786));
    Odrv4 I__3401 (
            .O(N__23786),
            .I(\current_shift_inst.control_inputZ0Z_2 ));
    InMux I__3400 (
            .O(N__23783),
            .I(N__23780));
    LocalMux I__3399 (
            .O(N__23780),
            .I(N__23775));
    InMux I__3398 (
            .O(N__23779),
            .I(N__23772));
    InMux I__3397 (
            .O(N__23778),
            .I(N__23769));
    Span4Mux_h I__3396 (
            .O(N__23775),
            .I(N__23762));
    LocalMux I__3395 (
            .O(N__23772),
            .I(N__23762));
    LocalMux I__3394 (
            .O(N__23769),
            .I(N__23762));
    Odrv4 I__3393 (
            .O(N__23762),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    InMux I__3392 (
            .O(N__23759),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ));
    InMux I__3391 (
            .O(N__23756),
            .I(N__23750));
    InMux I__3390 (
            .O(N__23755),
            .I(N__23743));
    InMux I__3389 (
            .O(N__23754),
            .I(N__23743));
    InMux I__3388 (
            .O(N__23753),
            .I(N__23743));
    LocalMux I__3387 (
            .O(N__23750),
            .I(N__23738));
    LocalMux I__3386 (
            .O(N__23743),
            .I(N__23738));
    Odrv4 I__3385 (
            .O(N__23738),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    CascadeMux I__3384 (
            .O(N__23735),
            .I(N__23731));
    InMux I__3383 (
            .O(N__23734),
            .I(N__23728));
    InMux I__3382 (
            .O(N__23731),
            .I(N__23725));
    LocalMux I__3381 (
            .O(N__23728),
            .I(N__23722));
    LocalMux I__3380 (
            .O(N__23725),
            .I(N__23719));
    Span4Mux_h I__3379 (
            .O(N__23722),
            .I(N__23714));
    Span4Mux_h I__3378 (
            .O(N__23719),
            .I(N__23714));
    Odrv4 I__3377 (
            .O(N__23714),
            .I(\current_shift_inst.control_inputZ0Z_3 ));
    InMux I__3376 (
            .O(N__23711),
            .I(N__23705));
    InMux I__3375 (
            .O(N__23710),
            .I(N__23700));
    InMux I__3374 (
            .O(N__23709),
            .I(N__23700));
    InMux I__3373 (
            .O(N__23708),
            .I(N__23697));
    LocalMux I__3372 (
            .O(N__23705),
            .I(N__23692));
    LocalMux I__3371 (
            .O(N__23700),
            .I(N__23692));
    LocalMux I__3370 (
            .O(N__23697),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    Odrv12 I__3369 (
            .O(N__23692),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    InMux I__3368 (
            .O(N__23687),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ));
    CEMux I__3367 (
            .O(N__23684),
            .I(N__23680));
    CEMux I__3366 (
            .O(N__23683),
            .I(N__23668));
    LocalMux I__3365 (
            .O(N__23680),
            .I(N__23665));
    CEMux I__3364 (
            .O(N__23679),
            .I(N__23662));
    CEMux I__3363 (
            .O(N__23678),
            .I(N__23659));
    CEMux I__3362 (
            .O(N__23677),
            .I(N__23656));
    CEMux I__3361 (
            .O(N__23676),
            .I(N__23653));
    CEMux I__3360 (
            .O(N__23675),
            .I(N__23650));
    CEMux I__3359 (
            .O(N__23674),
            .I(N__23645));
    CEMux I__3358 (
            .O(N__23673),
            .I(N__23642));
    CEMux I__3357 (
            .O(N__23672),
            .I(N__23638));
    CEMux I__3356 (
            .O(N__23671),
            .I(N__23632));
    LocalMux I__3355 (
            .O(N__23668),
            .I(N__23628));
    Span4Mux_h I__3354 (
            .O(N__23665),
            .I(N__23623));
    LocalMux I__3353 (
            .O(N__23662),
            .I(N__23623));
    LocalMux I__3352 (
            .O(N__23659),
            .I(N__23616));
    LocalMux I__3351 (
            .O(N__23656),
            .I(N__23616));
    LocalMux I__3350 (
            .O(N__23653),
            .I(N__23616));
    LocalMux I__3349 (
            .O(N__23650),
            .I(N__23613));
    CEMux I__3348 (
            .O(N__23649),
            .I(N__23610));
    CEMux I__3347 (
            .O(N__23648),
            .I(N__23607));
    LocalMux I__3346 (
            .O(N__23645),
            .I(N__23604));
    LocalMux I__3345 (
            .O(N__23642),
            .I(N__23601));
    CEMux I__3344 (
            .O(N__23641),
            .I(N__23598));
    LocalMux I__3343 (
            .O(N__23638),
            .I(N__23595));
    CEMux I__3342 (
            .O(N__23637),
            .I(N__23592));
    CEMux I__3341 (
            .O(N__23636),
            .I(N__23589));
    CEMux I__3340 (
            .O(N__23635),
            .I(N__23586));
    LocalMux I__3339 (
            .O(N__23632),
            .I(N__23582));
    CEMux I__3338 (
            .O(N__23631),
            .I(N__23579));
    Span4Mux_v I__3337 (
            .O(N__23628),
            .I(N__23573));
    Span4Mux_v I__3336 (
            .O(N__23623),
            .I(N__23573));
    Span4Mux_v I__3335 (
            .O(N__23616),
            .I(N__23566));
    Span4Mux_v I__3334 (
            .O(N__23613),
            .I(N__23566));
    LocalMux I__3333 (
            .O(N__23610),
            .I(N__23566));
    LocalMux I__3332 (
            .O(N__23607),
            .I(N__23563));
    Span4Mux_v I__3331 (
            .O(N__23604),
            .I(N__23560));
    Span4Mux_v I__3330 (
            .O(N__23601),
            .I(N__23555));
    LocalMux I__3329 (
            .O(N__23598),
            .I(N__23555));
    Span4Mux_h I__3328 (
            .O(N__23595),
            .I(N__23552));
    LocalMux I__3327 (
            .O(N__23592),
            .I(N__23545));
    LocalMux I__3326 (
            .O(N__23589),
            .I(N__23545));
    LocalMux I__3325 (
            .O(N__23586),
            .I(N__23545));
    CEMux I__3324 (
            .O(N__23585),
            .I(N__23542));
    Sp12to4 I__3323 (
            .O(N__23582),
            .I(N__23537));
    LocalMux I__3322 (
            .O(N__23579),
            .I(N__23537));
    CEMux I__3321 (
            .O(N__23578),
            .I(N__23534));
    Span4Mux_v I__3320 (
            .O(N__23573),
            .I(N__23531));
    Span4Mux_v I__3319 (
            .O(N__23566),
            .I(N__23526));
    Span4Mux_h I__3318 (
            .O(N__23563),
            .I(N__23526));
    Span4Mux_h I__3317 (
            .O(N__23560),
            .I(N__23517));
    Span4Mux_v I__3316 (
            .O(N__23555),
            .I(N__23517));
    Span4Mux_h I__3315 (
            .O(N__23552),
            .I(N__23517));
    Span4Mux_v I__3314 (
            .O(N__23545),
            .I(N__23517));
    LocalMux I__3313 (
            .O(N__23542),
            .I(N__23514));
    Span12Mux_v I__3312 (
            .O(N__23537),
            .I(N__23509));
    LocalMux I__3311 (
            .O(N__23534),
            .I(N__23509));
    Odrv4 I__3310 (
            .O(N__23531),
            .I(N_702_g));
    Odrv4 I__3309 (
            .O(N__23526),
            .I(N_702_g));
    Odrv4 I__3308 (
            .O(N__23517),
            .I(N_702_g));
    Odrv12 I__3307 (
            .O(N__23514),
            .I(N_702_g));
    Odrv12 I__3306 (
            .O(N__23509),
            .I(N_702_g));
    CascadeMux I__3305 (
            .O(N__23498),
            .I(N__23494));
    InMux I__3304 (
            .O(N__23497),
            .I(N__23490));
    InMux I__3303 (
            .O(N__23494),
            .I(N__23486));
    InMux I__3302 (
            .O(N__23493),
            .I(N__23483));
    LocalMux I__3301 (
            .O(N__23490),
            .I(N__23480));
    InMux I__3300 (
            .O(N__23489),
            .I(N__23477));
    LocalMux I__3299 (
            .O(N__23486),
            .I(N__23468));
    LocalMux I__3298 (
            .O(N__23483),
            .I(N__23468));
    Span4Mux_h I__3297 (
            .O(N__23480),
            .I(N__23468));
    LocalMux I__3296 (
            .O(N__23477),
            .I(N__23468));
    Span4Mux_h I__3295 (
            .O(N__23468),
            .I(N__23465));
    Odrv4 I__3294 (
            .O(N__23465),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    CascadeMux I__3293 (
            .O(N__23462),
            .I(N__23458));
    InMux I__3292 (
            .O(N__23461),
            .I(N__23455));
    InMux I__3291 (
            .O(N__23458),
            .I(N__23452));
    LocalMux I__3290 (
            .O(N__23455),
            .I(N__23449));
    LocalMux I__3289 (
            .O(N__23452),
            .I(N__23446));
    Span4Mux_h I__3288 (
            .O(N__23449),
            .I(N__23441));
    Span4Mux_h I__3287 (
            .O(N__23446),
            .I(N__23441));
    Odrv4 I__3286 (
            .O(N__23441),
            .I(\current_shift_inst.control_inputZ0Z_4 ));
    CascadeMux I__3285 (
            .O(N__23438),
            .I(N__23435));
    InMux I__3284 (
            .O(N__23435),
            .I(N__23432));
    LocalMux I__3283 (
            .O(N__23432),
            .I(N__23429));
    Span4Mux_h I__3282 (
            .O(N__23429),
            .I(N__23426));
    Odrv4 I__3281 (
            .O(N__23426),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ));
    InMux I__3280 (
            .O(N__23423),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ));
    CascadeMux I__3279 (
            .O(N__23420),
            .I(N__23417));
    InMux I__3278 (
            .O(N__23417),
            .I(N__23414));
    LocalMux I__3277 (
            .O(N__23414),
            .I(N__23411));
    Odrv4 I__3276 (
            .O(N__23411),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ));
    CascadeMux I__3275 (
            .O(N__23408),
            .I(N__23405));
    InMux I__3274 (
            .O(N__23405),
            .I(N__23402));
    LocalMux I__3273 (
            .O(N__23402),
            .I(N__23399));
    Odrv4 I__3272 (
            .O(N__23399),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ));
    CascadeMux I__3271 (
            .O(N__23396),
            .I(N__23393));
    InMux I__3270 (
            .O(N__23393),
            .I(N__23390));
    LocalMux I__3269 (
            .O(N__23390),
            .I(N__23387));
    Span4Mux_h I__3268 (
            .O(N__23387),
            .I(N__23384));
    Odrv4 I__3267 (
            .O(N__23384),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ));
    CascadeMux I__3266 (
            .O(N__23381),
            .I(N__23378));
    InMux I__3265 (
            .O(N__23378),
            .I(N__23375));
    LocalMux I__3264 (
            .O(N__23375),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_0 ));
    CascadeMux I__3263 (
            .O(N__23372),
            .I(N__23369));
    InMux I__3262 (
            .O(N__23369),
            .I(N__23366));
    LocalMux I__3261 (
            .O(N__23366),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ));
    CascadeMux I__3260 (
            .O(N__23363),
            .I(N__23360));
    InMux I__3259 (
            .O(N__23360),
            .I(N__23357));
    LocalMux I__3258 (
            .O(N__23357),
            .I(N__23354));
    Odrv4 I__3257 (
            .O(N__23354),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ));
    CascadeMux I__3256 (
            .O(N__23351),
            .I(N__23348));
    InMux I__3255 (
            .O(N__23348),
            .I(N__23345));
    LocalMux I__3254 (
            .O(N__23345),
            .I(N__23342));
    Odrv4 I__3253 (
            .O(N__23342),
            .I(\pwm_generator_inst.thresholdZ0Z_6 ));
    InMux I__3252 (
            .O(N__23339),
            .I(N__23336));
    LocalMux I__3251 (
            .O(N__23336),
            .I(\pwm_generator_inst.counter_i_6 ));
    InMux I__3250 (
            .O(N__23333),
            .I(N__23330));
    LocalMux I__3249 (
            .O(N__23330),
            .I(N__23327));
    Odrv12 I__3248 (
            .O(N__23327),
            .I(\pwm_generator_inst.thresholdZ0Z_7 ));
    CascadeMux I__3247 (
            .O(N__23324),
            .I(N__23321));
    InMux I__3246 (
            .O(N__23321),
            .I(N__23318));
    LocalMux I__3245 (
            .O(N__23318),
            .I(\pwm_generator_inst.counter_i_7 ));
    CascadeMux I__3244 (
            .O(N__23315),
            .I(N__23312));
    InMux I__3243 (
            .O(N__23312),
            .I(N__23309));
    LocalMux I__3242 (
            .O(N__23309),
            .I(N__23306));
    Span4Mux_h I__3241 (
            .O(N__23306),
            .I(N__23303));
    Odrv4 I__3240 (
            .O(N__23303),
            .I(\pwm_generator_inst.thresholdZ0Z_8 ));
    InMux I__3239 (
            .O(N__23300),
            .I(N__23297));
    LocalMux I__3238 (
            .O(N__23297),
            .I(\pwm_generator_inst.counter_i_8 ));
    CascadeMux I__3237 (
            .O(N__23294),
            .I(N__23291));
    InMux I__3236 (
            .O(N__23291),
            .I(N__23288));
    LocalMux I__3235 (
            .O(N__23288),
            .I(N__23285));
    Span4Mux_h I__3234 (
            .O(N__23285),
            .I(N__23282));
    Odrv4 I__3233 (
            .O(N__23282),
            .I(\pwm_generator_inst.thresholdZ0Z_9 ));
    InMux I__3232 (
            .O(N__23279),
            .I(N__23276));
    LocalMux I__3231 (
            .O(N__23276),
            .I(\pwm_generator_inst.counter_i_9 ));
    InMux I__3230 (
            .O(N__23273),
            .I(\pwm_generator_inst.un14_counter_cry_9 ));
    IoInMux I__3229 (
            .O(N__23270),
            .I(N__23267));
    LocalMux I__3228 (
            .O(N__23267),
            .I(N__23264));
    Span4Mux_s3_v I__3227 (
            .O(N__23264),
            .I(N__23261));
    Span4Mux_v I__3226 (
            .O(N__23261),
            .I(N__23258));
    Span4Mux_h I__3225 (
            .O(N__23258),
            .I(N__23255));
    Span4Mux_h I__3224 (
            .O(N__23255),
            .I(N__23252));
    Span4Mux_h I__3223 (
            .O(N__23252),
            .I(N__23249));
    Odrv4 I__3222 (
            .O(N__23249),
            .I(pwm_output_c));
    InMux I__3221 (
            .O(N__23246),
            .I(N__23243));
    LocalMux I__3220 (
            .O(N__23243),
            .I(il_min_comp2_D1));
    InMux I__3219 (
            .O(N__23240),
            .I(N__23237));
    LocalMux I__3218 (
            .O(N__23237),
            .I(N__23234));
    Span4Mux_h I__3217 (
            .O(N__23234),
            .I(N__23231));
    Span4Mux_v I__3216 (
            .O(N__23231),
            .I(N__23228));
    Odrv4 I__3215 (
            .O(N__23228),
            .I(il_max_comp1_c));
    CascadeMux I__3214 (
            .O(N__23225),
            .I(N__23222));
    InMux I__3213 (
            .O(N__23222),
            .I(N__23219));
    LocalMux I__3212 (
            .O(N__23219),
            .I(\pwm_generator_inst.thresholdZ0Z_0 ));
    InMux I__3211 (
            .O(N__23216),
            .I(N__23213));
    LocalMux I__3210 (
            .O(N__23213),
            .I(\pwm_generator_inst.counter_i_0 ));
    InMux I__3209 (
            .O(N__23210),
            .I(N__23207));
    LocalMux I__3208 (
            .O(N__23207),
            .I(N__23204));
    Odrv4 I__3207 (
            .O(N__23204),
            .I(\pwm_generator_inst.thresholdZ0Z_1 ));
    CascadeMux I__3206 (
            .O(N__23201),
            .I(N__23198));
    InMux I__3205 (
            .O(N__23198),
            .I(N__23195));
    LocalMux I__3204 (
            .O(N__23195),
            .I(\pwm_generator_inst.counter_i_1 ));
    CascadeMux I__3203 (
            .O(N__23192),
            .I(N__23189));
    InMux I__3202 (
            .O(N__23189),
            .I(N__23186));
    LocalMux I__3201 (
            .O(N__23186),
            .I(N__23183));
    Odrv12 I__3200 (
            .O(N__23183),
            .I(\pwm_generator_inst.thresholdZ0Z_2 ));
    InMux I__3199 (
            .O(N__23180),
            .I(N__23177));
    LocalMux I__3198 (
            .O(N__23177),
            .I(\pwm_generator_inst.counter_i_2 ));
    InMux I__3197 (
            .O(N__23174),
            .I(N__23171));
    LocalMux I__3196 (
            .O(N__23171),
            .I(\pwm_generator_inst.thresholdZ0Z_3 ));
    CascadeMux I__3195 (
            .O(N__23168),
            .I(N__23165));
    InMux I__3194 (
            .O(N__23165),
            .I(N__23162));
    LocalMux I__3193 (
            .O(N__23162),
            .I(\pwm_generator_inst.counter_i_3 ));
    InMux I__3192 (
            .O(N__23159),
            .I(N__23156));
    LocalMux I__3191 (
            .O(N__23156),
            .I(N__23153));
    Span4Mux_h I__3190 (
            .O(N__23153),
            .I(N__23150));
    Odrv4 I__3189 (
            .O(N__23150),
            .I(\pwm_generator_inst.thresholdZ0Z_4 ));
    CascadeMux I__3188 (
            .O(N__23147),
            .I(N__23144));
    InMux I__3187 (
            .O(N__23144),
            .I(N__23141));
    LocalMux I__3186 (
            .O(N__23141),
            .I(N__23138));
    Odrv4 I__3185 (
            .O(N__23138),
            .I(\pwm_generator_inst.counter_i_4 ));
    CascadeMux I__3184 (
            .O(N__23135),
            .I(N__23132));
    InMux I__3183 (
            .O(N__23132),
            .I(N__23129));
    LocalMux I__3182 (
            .O(N__23129),
            .I(N__23126));
    Odrv4 I__3181 (
            .O(N__23126),
            .I(\pwm_generator_inst.thresholdZ0Z_5 ));
    InMux I__3180 (
            .O(N__23123),
            .I(N__23120));
    LocalMux I__3179 (
            .O(N__23120),
            .I(\pwm_generator_inst.counter_i_5 ));
    InMux I__3178 (
            .O(N__23117),
            .I(N__23114));
    LocalMux I__3177 (
            .O(N__23114),
            .I(\current_shift_inst.control_input_1_axb_18 ));
    InMux I__3176 (
            .O(N__23111),
            .I(\current_shift_inst.un38_control_input_0_cry_23 ));
    InMux I__3175 (
            .O(N__23108),
            .I(N__23105));
    LocalMux I__3174 (
            .O(N__23105),
            .I(\current_shift_inst.control_input_1_axb_19 ));
    InMux I__3173 (
            .O(N__23102),
            .I(\current_shift_inst.un38_control_input_0_cry_24 ));
    InMux I__3172 (
            .O(N__23099),
            .I(N__23096));
    LocalMux I__3171 (
            .O(N__23096),
            .I(\current_shift_inst.control_input_1_axb_20 ));
    InMux I__3170 (
            .O(N__23093),
            .I(\current_shift_inst.un38_control_input_0_cry_25 ));
    InMux I__3169 (
            .O(N__23090),
            .I(N__23087));
    LocalMux I__3168 (
            .O(N__23087),
            .I(\current_shift_inst.control_input_1_axb_21 ));
    InMux I__3167 (
            .O(N__23084),
            .I(\current_shift_inst.un38_control_input_0_cry_26 ));
    InMux I__3166 (
            .O(N__23081),
            .I(N__23078));
    LocalMux I__3165 (
            .O(N__23078),
            .I(\current_shift_inst.control_input_1_axb_22 ));
    InMux I__3164 (
            .O(N__23075),
            .I(\current_shift_inst.un38_control_input_0_cry_27 ));
    InMux I__3163 (
            .O(N__23072),
            .I(N__23069));
    LocalMux I__3162 (
            .O(N__23069),
            .I(\current_shift_inst.control_input_1_axb_23 ));
    InMux I__3161 (
            .O(N__23066),
            .I(\current_shift_inst.un38_control_input_0_cry_28 ));
    InMux I__3160 (
            .O(N__23063),
            .I(N__23060));
    LocalMux I__3159 (
            .O(N__23060),
            .I(\current_shift_inst.control_input_1_axb_24 ));
    InMux I__3158 (
            .O(N__23057),
            .I(\current_shift_inst.un38_control_input_0_cry_29 ));
    CascadeMux I__3157 (
            .O(N__23054),
            .I(N__23051));
    InMux I__3156 (
            .O(N__23051),
            .I(N__23048));
    LocalMux I__3155 (
            .O(N__23048),
            .I(\current_shift_inst.control_input_1_cry_24_THRU_CO ));
    InMux I__3154 (
            .O(N__23045),
            .I(bfn_8_21_0_));
    CEMux I__3153 (
            .O(N__23042),
            .I(N__23039));
    LocalMux I__3152 (
            .O(N__23039),
            .I(N__23034));
    CEMux I__3151 (
            .O(N__23038),
            .I(N__23031));
    CEMux I__3150 (
            .O(N__23037),
            .I(N__23028));
    Span4Mux_h I__3149 (
            .O(N__23034),
            .I(N__23021));
    LocalMux I__3148 (
            .O(N__23031),
            .I(N__23021));
    LocalMux I__3147 (
            .O(N__23028),
            .I(N__23018));
    CEMux I__3146 (
            .O(N__23027),
            .I(N__23015));
    CEMux I__3145 (
            .O(N__23026),
            .I(N__23012));
    Span4Mux_v I__3144 (
            .O(N__23021),
            .I(N__23005));
    Span4Mux_v I__3143 (
            .O(N__23018),
            .I(N__23005));
    LocalMux I__3142 (
            .O(N__23015),
            .I(N__23005));
    LocalMux I__3141 (
            .O(N__23012),
            .I(N__23002));
    Span4Mux_v I__3140 (
            .O(N__23005),
            .I(N__22999));
    Span12Mux_v I__3139 (
            .O(N__23002),
            .I(N__22996));
    Span4Mux_v I__3138 (
            .O(N__22999),
            .I(N__22993));
    Odrv12 I__3137 (
            .O(N__22996),
            .I(\current_shift_inst.phase_valid_RNISLORZ0Z2 ));
    Odrv4 I__3136 (
            .O(N__22993),
            .I(\current_shift_inst.phase_valid_RNISLORZ0Z2 ));
    InMux I__3135 (
            .O(N__22988),
            .I(N__22985));
    LocalMux I__3134 (
            .O(N__22985),
            .I(\current_shift_inst.control_input_1_axb_9 ));
    InMux I__3133 (
            .O(N__22982),
            .I(bfn_8_19_0_));
    InMux I__3132 (
            .O(N__22979),
            .I(N__22976));
    LocalMux I__3131 (
            .O(N__22976),
            .I(\current_shift_inst.control_input_1_axb_10 ));
    InMux I__3130 (
            .O(N__22973),
            .I(\current_shift_inst.un38_control_input_0_cry_15 ));
    InMux I__3129 (
            .O(N__22970),
            .I(N__22967));
    LocalMux I__3128 (
            .O(N__22967),
            .I(\current_shift_inst.control_input_1_axb_11 ));
    InMux I__3127 (
            .O(N__22964),
            .I(\current_shift_inst.un38_control_input_0_cry_16 ));
    CascadeMux I__3126 (
            .O(N__22961),
            .I(N__22958));
    InMux I__3125 (
            .O(N__22958),
            .I(N__22955));
    LocalMux I__3124 (
            .O(N__22955),
            .I(N__22952));
    Odrv4 I__3123 (
            .O(N__22952),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIH6661_17 ));
    InMux I__3122 (
            .O(N__22949),
            .I(N__22946));
    LocalMux I__3121 (
            .O(N__22946),
            .I(\current_shift_inst.control_input_1_axb_12 ));
    InMux I__3120 (
            .O(N__22943),
            .I(\current_shift_inst.un38_control_input_0_cry_17 ));
    CascadeMux I__3119 (
            .O(N__22940),
            .I(N__22937));
    InMux I__3118 (
            .O(N__22937),
            .I(N__22934));
    LocalMux I__3117 (
            .O(N__22934),
            .I(N__22931));
    Odrv12 I__3116 (
            .O(N__22931),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIAL3J_18 ));
    InMux I__3115 (
            .O(N__22928),
            .I(N__22925));
    LocalMux I__3114 (
            .O(N__22925),
            .I(\current_shift_inst.control_input_1_axb_13 ));
    InMux I__3113 (
            .O(N__22922),
            .I(\current_shift_inst.un38_control_input_0_cry_18 ));
    CascadeMux I__3112 (
            .O(N__22919),
            .I(N__22916));
    InMux I__3111 (
            .O(N__22916),
            .I(N__22913));
    LocalMux I__3110 (
            .O(N__22913),
            .I(N__22910));
    Odrv4 I__3109 (
            .O(N__22910),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI4H5J_19 ));
    InMux I__3108 (
            .O(N__22907),
            .I(N__22904));
    LocalMux I__3107 (
            .O(N__22904),
            .I(\current_shift_inst.control_input_1_axb_14 ));
    InMux I__3106 (
            .O(N__22901),
            .I(\current_shift_inst.un38_control_input_0_cry_19 ));
    InMux I__3105 (
            .O(N__22898),
            .I(N__22895));
    LocalMux I__3104 (
            .O(N__22895),
            .I(\current_shift_inst.control_input_1_axb_15 ));
    InMux I__3103 (
            .O(N__22892),
            .I(\current_shift_inst.un38_control_input_0_cry_20 ));
    InMux I__3102 (
            .O(N__22889),
            .I(N__22886));
    LocalMux I__3101 (
            .O(N__22886),
            .I(\current_shift_inst.control_input_1_axb_16 ));
    InMux I__3100 (
            .O(N__22883),
            .I(\current_shift_inst.un38_control_input_0_cry_21 ));
    InMux I__3099 (
            .O(N__22880),
            .I(N__22877));
    LocalMux I__3098 (
            .O(N__22877),
            .I(\current_shift_inst.control_input_1_axb_17 ));
    InMux I__3097 (
            .O(N__22874),
            .I(bfn_8_20_0_));
    InMux I__3096 (
            .O(N__22871),
            .I(N__22868));
    LocalMux I__3095 (
            .O(N__22868),
            .I(\current_shift_inst.control_input_1_axb_1 ));
    InMux I__3094 (
            .O(N__22865),
            .I(bfn_8_18_0_));
    InMux I__3093 (
            .O(N__22862),
            .I(N__22859));
    LocalMux I__3092 (
            .O(N__22859),
            .I(\current_shift_inst.control_input_1_axb_2 ));
    InMux I__3091 (
            .O(N__22856),
            .I(\current_shift_inst.un38_control_input_0_cry_7 ));
    InMux I__3090 (
            .O(N__22853),
            .I(N__22850));
    LocalMux I__3089 (
            .O(N__22850),
            .I(\current_shift_inst.control_input_1_axb_3 ));
    InMux I__3088 (
            .O(N__22847),
            .I(\current_shift_inst.un38_control_input_0_cry_8 ));
    InMux I__3087 (
            .O(N__22844),
            .I(N__22841));
    LocalMux I__3086 (
            .O(N__22841),
            .I(\current_shift_inst.control_input_1_axb_4 ));
    InMux I__3085 (
            .O(N__22838),
            .I(\current_shift_inst.un38_control_input_0_cry_9 ));
    InMux I__3084 (
            .O(N__22835),
            .I(N__22832));
    LocalMux I__3083 (
            .O(N__22832),
            .I(\current_shift_inst.control_input_1_axb_5 ));
    InMux I__3082 (
            .O(N__22829),
            .I(\current_shift_inst.un38_control_input_0_cry_10 ));
    InMux I__3081 (
            .O(N__22826),
            .I(N__22823));
    LocalMux I__3080 (
            .O(N__22823),
            .I(\current_shift_inst.control_input_1_axb_6 ));
    InMux I__3079 (
            .O(N__22820),
            .I(\current_shift_inst.un38_control_input_0_cry_11 ));
    InMux I__3078 (
            .O(N__22817),
            .I(N__22814));
    LocalMux I__3077 (
            .O(N__22814),
            .I(\current_shift_inst.control_input_1_axb_7 ));
    InMux I__3076 (
            .O(N__22811),
            .I(\current_shift_inst.un38_control_input_0_cry_12 ));
    CascadeMux I__3075 (
            .O(N__22808),
            .I(N__22805));
    InMux I__3074 (
            .O(N__22805),
            .I(N__22802));
    LocalMux I__3073 (
            .O(N__22802),
            .I(N__22799));
    Odrv4 I__3072 (
            .O(N__22799),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIR0UI_13 ));
    InMux I__3071 (
            .O(N__22796),
            .I(N__22793));
    LocalMux I__3070 (
            .O(N__22793),
            .I(\current_shift_inst.control_input_1_axb_8 ));
    InMux I__3069 (
            .O(N__22790),
            .I(\current_shift_inst.un38_control_input_0_cry_13 ));
    InMux I__3068 (
            .O(N__22787),
            .I(N__22784));
    LocalMux I__3067 (
            .O(N__22784),
            .I(\current_shift_inst.z_i_0_31 ));
    CascadeMux I__3066 (
            .O(N__22781),
            .I(N__22778));
    InMux I__3065 (
            .O(N__22778),
            .I(N__22775));
    LocalMux I__3064 (
            .O(N__22775),
            .I(\current_shift_inst.un38_control_input_0_cry_3_c_invZ0 ));
    InMux I__3063 (
            .O(N__22772),
            .I(N__22769));
    LocalMux I__3062 (
            .O(N__22769),
            .I(\current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0 ));
    CascadeMux I__3061 (
            .O(N__22766),
            .I(N__22763));
    InMux I__3060 (
            .O(N__22763),
            .I(N__22760));
    LocalMux I__3059 (
            .O(N__22760),
            .I(\current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0Z_0 ));
    InMux I__3058 (
            .O(N__22757),
            .I(N__22754));
    LocalMux I__3057 (
            .O(N__22754),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIVQKU1_5 ));
    InMux I__3056 (
            .O(N__22751),
            .I(N__22748));
    LocalMux I__3055 (
            .O(N__22748),
            .I(\current_shift_inst.control_input_1_axb_0 ));
    InMux I__3054 (
            .O(N__22745),
            .I(\current_shift_inst.un38_control_input_0_cry_5 ));
    InMux I__3053 (
            .O(N__22742),
            .I(N__22727));
    InMux I__3052 (
            .O(N__22741),
            .I(N__22727));
    InMux I__3051 (
            .O(N__22740),
            .I(N__22714));
    InMux I__3050 (
            .O(N__22739),
            .I(N__22714));
    InMux I__3049 (
            .O(N__22738),
            .I(N__22699));
    InMux I__3048 (
            .O(N__22737),
            .I(N__22699));
    InMux I__3047 (
            .O(N__22736),
            .I(N__22699));
    InMux I__3046 (
            .O(N__22735),
            .I(N__22699));
    InMux I__3045 (
            .O(N__22734),
            .I(N__22699));
    InMux I__3044 (
            .O(N__22733),
            .I(N__22699));
    InMux I__3043 (
            .O(N__22732),
            .I(N__22699));
    LocalMux I__3042 (
            .O(N__22727),
            .I(N__22696));
    InMux I__3041 (
            .O(N__22726),
            .I(N__22691));
    InMux I__3040 (
            .O(N__22725),
            .I(N__22691));
    InMux I__3039 (
            .O(N__22724),
            .I(N__22669));
    InMux I__3038 (
            .O(N__22723),
            .I(N__22669));
    InMux I__3037 (
            .O(N__22722),
            .I(N__22669));
    InMux I__3036 (
            .O(N__22721),
            .I(N__22669));
    InMux I__3035 (
            .O(N__22720),
            .I(N__22669));
    InMux I__3034 (
            .O(N__22719),
            .I(N__22669));
    LocalMux I__3033 (
            .O(N__22714),
            .I(N__22666));
    LocalMux I__3032 (
            .O(N__22699),
            .I(N__22663));
    Span4Mux_v I__3031 (
            .O(N__22696),
            .I(N__22658));
    LocalMux I__3030 (
            .O(N__22691),
            .I(N__22658));
    InMux I__3029 (
            .O(N__22690),
            .I(N__22653));
    InMux I__3028 (
            .O(N__22689),
            .I(N__22653));
    InMux I__3027 (
            .O(N__22688),
            .I(N__22638));
    InMux I__3026 (
            .O(N__22687),
            .I(N__22638));
    InMux I__3025 (
            .O(N__22686),
            .I(N__22638));
    InMux I__3024 (
            .O(N__22685),
            .I(N__22638));
    InMux I__3023 (
            .O(N__22684),
            .I(N__22638));
    InMux I__3022 (
            .O(N__22683),
            .I(N__22638));
    InMux I__3021 (
            .O(N__22682),
            .I(N__22638));
    LocalMux I__3020 (
            .O(N__22669),
            .I(\current_shift_inst.PI_CTRL.N_76 ));
    Odrv4 I__3019 (
            .O(N__22666),
            .I(\current_shift_inst.PI_CTRL.N_76 ));
    Odrv4 I__3018 (
            .O(N__22663),
            .I(\current_shift_inst.PI_CTRL.N_76 ));
    Odrv4 I__3017 (
            .O(N__22658),
            .I(\current_shift_inst.PI_CTRL.N_76 ));
    LocalMux I__3016 (
            .O(N__22653),
            .I(\current_shift_inst.PI_CTRL.N_76 ));
    LocalMux I__3015 (
            .O(N__22638),
            .I(\current_shift_inst.PI_CTRL.N_76 ));
    CascadeMux I__3014 (
            .O(N__22625),
            .I(N__22616));
    CascadeMux I__3013 (
            .O(N__22624),
            .I(N__22605));
    CascadeMux I__3012 (
            .O(N__22623),
            .I(N__22601));
    CascadeMux I__3011 (
            .O(N__22622),
            .I(N__22598));
    CascadeMux I__3010 (
            .O(N__22621),
            .I(N__22595));
    CascadeMux I__3009 (
            .O(N__22620),
            .I(N__22592));
    InMux I__3008 (
            .O(N__22619),
            .I(N__22584));
    InMux I__3007 (
            .O(N__22616),
            .I(N__22584));
    InMux I__3006 (
            .O(N__22615),
            .I(N__22581));
    InMux I__3005 (
            .O(N__22614),
            .I(N__22578));
    CascadeMux I__3004 (
            .O(N__22613),
            .I(N__22571));
    CascadeMux I__3003 (
            .O(N__22612),
            .I(N__22568));
    CascadeMux I__3002 (
            .O(N__22611),
            .I(N__22565));
    CascadeMux I__3001 (
            .O(N__22610),
            .I(N__22562));
    CascadeMux I__3000 (
            .O(N__22609),
            .I(N__22559));
    CascadeMux I__2999 (
            .O(N__22608),
            .I(N__22556));
    InMux I__2998 (
            .O(N__22605),
            .I(N__22546));
    InMux I__2997 (
            .O(N__22604),
            .I(N__22546));
    InMux I__2996 (
            .O(N__22601),
            .I(N__22531));
    InMux I__2995 (
            .O(N__22598),
            .I(N__22531));
    InMux I__2994 (
            .O(N__22595),
            .I(N__22531));
    InMux I__2993 (
            .O(N__22592),
            .I(N__22531));
    InMux I__2992 (
            .O(N__22591),
            .I(N__22531));
    InMux I__2991 (
            .O(N__22590),
            .I(N__22531));
    InMux I__2990 (
            .O(N__22589),
            .I(N__22531));
    LocalMux I__2989 (
            .O(N__22584),
            .I(N__22528));
    LocalMux I__2988 (
            .O(N__22581),
            .I(N__22523));
    LocalMux I__2987 (
            .O(N__22578),
            .I(N__22523));
    InMux I__2986 (
            .O(N__22577),
            .I(N__22510));
    InMux I__2985 (
            .O(N__22576),
            .I(N__22510));
    InMux I__2984 (
            .O(N__22575),
            .I(N__22510));
    InMux I__2983 (
            .O(N__22574),
            .I(N__22510));
    InMux I__2982 (
            .O(N__22571),
            .I(N__22510));
    InMux I__2981 (
            .O(N__22568),
            .I(N__22510));
    InMux I__2980 (
            .O(N__22565),
            .I(N__22495));
    InMux I__2979 (
            .O(N__22562),
            .I(N__22495));
    InMux I__2978 (
            .O(N__22559),
            .I(N__22495));
    InMux I__2977 (
            .O(N__22556),
            .I(N__22495));
    InMux I__2976 (
            .O(N__22555),
            .I(N__22495));
    InMux I__2975 (
            .O(N__22554),
            .I(N__22495));
    InMux I__2974 (
            .O(N__22553),
            .I(N__22495));
    InMux I__2973 (
            .O(N__22552),
            .I(N__22490));
    InMux I__2972 (
            .O(N__22551),
            .I(N__22490));
    LocalMux I__2971 (
            .O(N__22546),
            .I(N__22487));
    LocalMux I__2970 (
            .O(N__22531),
            .I(N__22484));
    Span4Mux_h I__2969 (
            .O(N__22528),
            .I(N__22479));
    Span4Mux_v I__2968 (
            .O(N__22523),
            .I(N__22479));
    LocalMux I__2967 (
            .O(N__22510),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    LocalMux I__2966 (
            .O(N__22495),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    LocalMux I__2965 (
            .O(N__22490),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    Odrv4 I__2964 (
            .O(N__22487),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    Odrv4 I__2963 (
            .O(N__22484),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    Odrv4 I__2962 (
            .O(N__22479),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    CascadeMux I__2961 (
            .O(N__22466),
            .I(N__22462));
    CascadeMux I__2960 (
            .O(N__22465),
            .I(N__22459));
    InMux I__2959 (
            .O(N__22462),
            .I(N__22456));
    InMux I__2958 (
            .O(N__22459),
            .I(N__22453));
    LocalMux I__2957 (
            .O(N__22456),
            .I(\current_shift_inst.PI_CTRL.N_47_16 ));
    LocalMux I__2956 (
            .O(N__22453),
            .I(\current_shift_inst.PI_CTRL.N_47_16 ));
    InMux I__2955 (
            .O(N__22448),
            .I(N__22444));
    InMux I__2954 (
            .O(N__22447),
            .I(N__22441));
    LocalMux I__2953 (
            .O(N__22444),
            .I(N__22436));
    LocalMux I__2952 (
            .O(N__22441),
            .I(N__22436));
    Odrv4 I__2951 (
            .O(N__22436),
            .I(\current_shift_inst.PI_CTRL.N_46_16 ));
    InMux I__2950 (
            .O(N__22433),
            .I(N__22430));
    LocalMux I__2949 (
            .O(N__22430),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_16 ));
    InMux I__2948 (
            .O(N__22427),
            .I(N__22424));
    LocalMux I__2947 (
            .O(N__22424),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_17 ));
    InMux I__2946 (
            .O(N__22421),
            .I(N__22418));
    LocalMux I__2945 (
            .O(N__22418),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_18 ));
    InMux I__2944 (
            .O(N__22415),
            .I(N__22412));
    LocalMux I__2943 (
            .O(N__22412),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_19 ));
    InMux I__2942 (
            .O(N__22409),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ));
    InMux I__2941 (
            .O(N__22406),
            .I(N__22403));
    LocalMux I__2940 (
            .O(N__22403),
            .I(\current_shift_inst.PI_CTRL.un1_enablelt3_0 ));
    CascadeMux I__2939 (
            .O(N__22400),
            .I(N__22397));
    InMux I__2938 (
            .O(N__22397),
            .I(N__22394));
    LocalMux I__2937 (
            .O(N__22394),
            .I(N__22391));
    Odrv4 I__2936 (
            .O(N__22391),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ));
    InMux I__2935 (
            .O(N__22388),
            .I(N__22385));
    LocalMux I__2934 (
            .O(N__22385),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ));
    InMux I__2933 (
            .O(N__22382),
            .I(N__22379));
    LocalMux I__2932 (
            .O(N__22379),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ));
    InMux I__2931 (
            .O(N__22376),
            .I(N__22373));
    LocalMux I__2930 (
            .O(N__22373),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ));
    InMux I__2929 (
            .O(N__22370),
            .I(N__22367));
    LocalMux I__2928 (
            .O(N__22367),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ));
    InMux I__2927 (
            .O(N__22364),
            .I(N__22361));
    LocalMux I__2926 (
            .O(N__22361),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ));
    InMux I__2925 (
            .O(N__22358),
            .I(N__22355));
    LocalMux I__2924 (
            .O(N__22355),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ));
    InMux I__2923 (
            .O(N__22352),
            .I(N__22349));
    LocalMux I__2922 (
            .O(N__22349),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ));
    InMux I__2921 (
            .O(N__22346),
            .I(N__22343));
    LocalMux I__2920 (
            .O(N__22343),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ));
    CascadeMux I__2919 (
            .O(N__22340),
            .I(N__22337));
    InMux I__2918 (
            .O(N__22337),
            .I(N__22334));
    LocalMux I__2917 (
            .O(N__22334),
            .I(N__22331));
    Span4Mux_h I__2916 (
            .O(N__22331),
            .I(N__22328));
    Span4Mux_h I__2915 (
            .O(N__22328),
            .I(N__22325));
    Odrv4 I__2914 (
            .O(N__22325),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ));
    InMux I__2913 (
            .O(N__22322),
            .I(N__22319));
    LocalMux I__2912 (
            .O(N__22319),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ));
    CascadeMux I__2911 (
            .O(N__22316),
            .I(N__22313));
    InMux I__2910 (
            .O(N__22313),
            .I(N__22310));
    LocalMux I__2909 (
            .O(N__22310),
            .I(N__22307));
    Span4Mux_v I__2908 (
            .O(N__22307),
            .I(N__22304));
    Span4Mux_h I__2907 (
            .O(N__22304),
            .I(N__22301));
    Odrv4 I__2906 (
            .O(N__22301),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ));
    InMux I__2905 (
            .O(N__22298),
            .I(N__22295));
    LocalMux I__2904 (
            .O(N__22295),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ));
    CascadeMux I__2903 (
            .O(N__22292),
            .I(N__22289));
    InMux I__2902 (
            .O(N__22289),
            .I(N__22286));
    LocalMux I__2901 (
            .O(N__22286),
            .I(N__22283));
    Span4Mux_h I__2900 (
            .O(N__22283),
            .I(N__22280));
    Span4Mux_h I__2899 (
            .O(N__22280),
            .I(N__22277));
    Odrv4 I__2898 (
            .O(N__22277),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ));
    InMux I__2897 (
            .O(N__22274),
            .I(N__22271));
    LocalMux I__2896 (
            .O(N__22271),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ));
    InMux I__2895 (
            .O(N__22268),
            .I(N__22265));
    LocalMux I__2894 (
            .O(N__22265),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ));
    InMux I__2893 (
            .O(N__22262),
            .I(N__22259));
    LocalMux I__2892 (
            .O(N__22259),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ));
    CascadeMux I__2891 (
            .O(N__22256),
            .I(N__22253));
    InMux I__2890 (
            .O(N__22253),
            .I(N__22250));
    LocalMux I__2889 (
            .O(N__22250),
            .I(N__22247));
    Span4Mux_h I__2888 (
            .O(N__22247),
            .I(N__22244));
    Span4Mux_h I__2887 (
            .O(N__22244),
            .I(N__22241));
    Odrv4 I__2886 (
            .O(N__22241),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ1Z_6 ));
    InMux I__2885 (
            .O(N__22238),
            .I(N__22235));
    LocalMux I__2884 (
            .O(N__22235),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ));
    InMux I__2883 (
            .O(N__22232),
            .I(N__22229));
    LocalMux I__2882 (
            .O(N__22229),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ));
    InMux I__2881 (
            .O(N__22226),
            .I(\current_shift_inst.control_input_1_cry_24 ));
    InMux I__2880 (
            .O(N__22223),
            .I(N__22220));
    LocalMux I__2879 (
            .O(N__22220),
            .I(N__22217));
    Span12Mux_h I__2878 (
            .O(N__22217),
            .I(N__22214));
    Odrv12 I__2877 (
            .O(N__22214),
            .I(il_min_comp2_c));
    InMux I__2876 (
            .O(N__22211),
            .I(N__22208));
    LocalMux I__2875 (
            .O(N__22208),
            .I(N__22205));
    Span4Mux_v I__2874 (
            .O(N__22205),
            .I(N__22202));
    Span4Mux_h I__2873 (
            .O(N__22202),
            .I(N__22199));
    Odrv4 I__2872 (
            .O(N__22199),
            .I(il_max_comp2_c));
    InMux I__2871 (
            .O(N__22196),
            .I(N__22193));
    LocalMux I__2870 (
            .O(N__22193),
            .I(N__22190));
    Span4Mux_v I__2869 (
            .O(N__22190),
            .I(N__22187));
    Odrv4 I__2868 (
            .O(N__22187),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_0 ));
    InMux I__2867 (
            .O(N__22184),
            .I(N__22181));
    LocalMux I__2866 (
            .O(N__22181),
            .I(N__22178));
    Span4Mux_h I__2865 (
            .O(N__22178),
            .I(N__22175));
    Odrv4 I__2864 (
            .O(N__22175),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_6 ));
    InMux I__2863 (
            .O(N__22172),
            .I(N__22169));
    LocalMux I__2862 (
            .O(N__22169),
            .I(N__22166));
    Odrv12 I__2861 (
            .O(N__22166),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_3 ));
    InMux I__2860 (
            .O(N__22163),
            .I(N__22160));
    LocalMux I__2859 (
            .O(N__22160),
            .I(N__22157));
    Odrv12 I__2858 (
            .O(N__22157),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_5 ));
    InMux I__2857 (
            .O(N__22154),
            .I(bfn_7_19_0_));
    InMux I__2856 (
            .O(N__22151),
            .I(\current_shift_inst.control_input_1_cry_16 ));
    InMux I__2855 (
            .O(N__22148),
            .I(\current_shift_inst.control_input_1_cry_17 ));
    InMux I__2854 (
            .O(N__22145),
            .I(\current_shift_inst.control_input_1_cry_18 ));
    InMux I__2853 (
            .O(N__22142),
            .I(\current_shift_inst.control_input_1_cry_19 ));
    InMux I__2852 (
            .O(N__22139),
            .I(\current_shift_inst.control_input_1_cry_20 ));
    InMux I__2851 (
            .O(N__22136),
            .I(\current_shift_inst.control_input_1_cry_21 ));
    InMux I__2850 (
            .O(N__22133),
            .I(\current_shift_inst.control_input_1_cry_22 ));
    InMux I__2849 (
            .O(N__22130),
            .I(bfn_7_20_0_));
    InMux I__2848 (
            .O(N__22127),
            .I(\current_shift_inst.control_input_1_cry_6 ));
    InMux I__2847 (
            .O(N__22124),
            .I(bfn_7_18_0_));
    InMux I__2846 (
            .O(N__22121),
            .I(\current_shift_inst.control_input_1_cry_8 ));
    InMux I__2845 (
            .O(N__22118),
            .I(\current_shift_inst.control_input_1_cry_9 ));
    InMux I__2844 (
            .O(N__22115),
            .I(\current_shift_inst.control_input_1_cry_10 ));
    InMux I__2843 (
            .O(N__22112),
            .I(\current_shift_inst.control_input_1_cry_11 ));
    InMux I__2842 (
            .O(N__22109),
            .I(\current_shift_inst.control_input_1_cry_12 ));
    InMux I__2841 (
            .O(N__22106),
            .I(\current_shift_inst.control_input_1_cry_13 ));
    InMux I__2840 (
            .O(N__22103),
            .I(\current_shift_inst.control_input_1_cry_14 ));
    InMux I__2839 (
            .O(N__22100),
            .I(\current_shift_inst.control_input_1_cry_0 ));
    InMux I__2838 (
            .O(N__22097),
            .I(\current_shift_inst.control_input_1_cry_1 ));
    InMux I__2837 (
            .O(N__22094),
            .I(\current_shift_inst.control_input_1_cry_2 ));
    InMux I__2836 (
            .O(N__22091),
            .I(\current_shift_inst.control_input_1_cry_3 ));
    InMux I__2835 (
            .O(N__22088),
            .I(\current_shift_inst.control_input_1_cry_4 ));
    InMux I__2834 (
            .O(N__22085),
            .I(\current_shift_inst.control_input_1_cry_5 ));
    InMux I__2833 (
            .O(N__22082),
            .I(N__22079));
    LocalMux I__2832 (
            .O(N__22079),
            .I(N__22076));
    Odrv4 I__2831 (
            .O(N__22076),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31 ));
    InMux I__2830 (
            .O(N__22073),
            .I(N__22070));
    LocalMux I__2829 (
            .O(N__22070),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31 ));
    CascadeMux I__2828 (
            .O(N__22067),
            .I(N__22064));
    InMux I__2827 (
            .O(N__22064),
            .I(N__22061));
    LocalMux I__2826 (
            .O(N__22061),
            .I(N__22058));
    Span4Mux_v I__2825 (
            .O(N__22058),
            .I(N__22055));
    Odrv4 I__2824 (
            .O(N__22055),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ));
    CascadeMux I__2823 (
            .O(N__22052),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_ ));
    InMux I__2822 (
            .O(N__22049),
            .I(N__22046));
    LocalMux I__2821 (
            .O(N__22046),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_3 ));
    CascadeMux I__2820 (
            .O(N__22043),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_2_cascade_ ));
    InMux I__2819 (
            .O(N__22040),
            .I(N__22037));
    LocalMux I__2818 (
            .O(N__22037),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_2 ));
    InMux I__2817 (
            .O(N__22034),
            .I(N__22028));
    InMux I__2816 (
            .O(N__22033),
            .I(N__22028));
    LocalMux I__2815 (
            .O(N__22028),
            .I(N__22025));
    Span4Mux_v I__2814 (
            .O(N__22025),
            .I(N__22022));
    Odrv4 I__2813 (
            .O(N__22022),
            .I(\current_shift_inst.PI_CTRL.N_47_21 ));
    InMux I__2812 (
            .O(N__22019),
            .I(N__22015));
    InMux I__2811 (
            .O(N__22018),
            .I(N__22012));
    LocalMux I__2810 (
            .O(N__22015),
            .I(\current_shift_inst.PI_CTRL.N_43 ));
    LocalMux I__2809 (
            .O(N__22012),
            .I(\current_shift_inst.PI_CTRL.N_43 ));
    CascadeMux I__2808 (
            .O(N__22007),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31_cascade_ ));
    InMux I__2807 (
            .O(N__22004),
            .I(N__22001));
    LocalMux I__2806 (
            .O(N__22001),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31 ));
    InMux I__2805 (
            .O(N__21998),
            .I(N__21995));
    LocalMux I__2804 (
            .O(N__21995),
            .I(\current_shift_inst.PI_CTRL.N_46_21 ));
    CascadeMux I__2803 (
            .O(N__21992),
            .I(\current_shift_inst.PI_CTRL.N_46_21_cascade_ ));
    InMux I__2802 (
            .O(N__21989),
            .I(N__21985));
    InMux I__2801 (
            .O(N__21988),
            .I(N__21982));
    LocalMux I__2800 (
            .O(N__21985),
            .I(\current_shift_inst.PI_CTRL.N_44 ));
    LocalMux I__2799 (
            .O(N__21982),
            .I(\current_shift_inst.PI_CTRL.N_44 ));
    InMux I__2798 (
            .O(N__21977),
            .I(N__21974));
    LocalMux I__2797 (
            .O(N__21974),
            .I(N__21971));
    Span4Mux_h I__2796 (
            .O(N__21971),
            .I(N__21968));
    Odrv4 I__2795 (
            .O(N__21968),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_1 ));
    InMux I__2794 (
            .O(N__21965),
            .I(N__21962));
    LocalMux I__2793 (
            .O(N__21962),
            .I(N__21959));
    Odrv4 I__2792 (
            .O(N__21959),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_4 ));
    InMux I__2791 (
            .O(N__21956),
            .I(N__21953));
    LocalMux I__2790 (
            .O(N__21953),
            .I(N__21950));
    Span4Mux_v I__2789 (
            .O(N__21950),
            .I(N__21947));
    Span4Mux_h I__2788 (
            .O(N__21947),
            .I(N__21944));
    Odrv4 I__2787 (
            .O(N__21944),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_9 ));
    CascadeMux I__2786 (
            .O(N__21941),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ));
    InMux I__2785 (
            .O(N__21938),
            .I(N__21935));
    LocalMux I__2784 (
            .O(N__21935),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_18 ));
    CascadeMux I__2783 (
            .O(N__21932),
            .I(N__21929));
    InMux I__2782 (
            .O(N__21929),
            .I(N__21926));
    LocalMux I__2781 (
            .O(N__21926),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_23 ));
    CascadeMux I__2780 (
            .O(N__21923),
            .I(N__21920));
    InMux I__2779 (
            .O(N__21920),
            .I(N__21917));
    LocalMux I__2778 (
            .O(N__21917),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_22 ));
    InMux I__2777 (
            .O(N__21914),
            .I(N__21911));
    LocalMux I__2776 (
            .O(N__21911),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_24 ));
    CascadeMux I__2775 (
            .O(N__21908),
            .I(N__21901));
    CascadeMux I__2774 (
            .O(N__21907),
            .I(N__21897));
    CascadeMux I__2773 (
            .O(N__21906),
            .I(N__21893));
    InMux I__2772 (
            .O(N__21905),
            .I(N__21878));
    InMux I__2771 (
            .O(N__21904),
            .I(N__21878));
    InMux I__2770 (
            .O(N__21901),
            .I(N__21878));
    InMux I__2769 (
            .O(N__21900),
            .I(N__21878));
    InMux I__2768 (
            .O(N__21897),
            .I(N__21878));
    InMux I__2767 (
            .O(N__21896),
            .I(N__21878));
    InMux I__2766 (
            .O(N__21893),
            .I(N__21878));
    LocalMux I__2765 (
            .O(N__21878),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_25 ));
    InMux I__2764 (
            .O(N__21875),
            .I(N__21872));
    LocalMux I__2763 (
            .O(N__21872),
            .I(N__21866));
    InMux I__2762 (
            .O(N__21871),
            .I(N__21859));
    InMux I__2761 (
            .O(N__21870),
            .I(N__21859));
    InMux I__2760 (
            .O(N__21869),
            .I(N__21859));
    Odrv4 I__2759 (
            .O(N__21866),
            .I(clk_10khz_i));
    LocalMux I__2758 (
            .O(N__21859),
            .I(clk_10khz_i));
    InMux I__2757 (
            .O(N__21854),
            .I(N__21851));
    LocalMux I__2756 (
            .O(N__21851),
            .I(N__21848));
    Odrv4 I__2755 (
            .O(N__21848),
            .I(clk_10khz_RNIIENAZ0Z2));
    InMux I__2754 (
            .O(N__21845),
            .I(N__21842));
    LocalMux I__2753 (
            .O(N__21842),
            .I(N__21839));
    Odrv12 I__2752 (
            .O(N__21839),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_7 ));
    InMux I__2751 (
            .O(N__21836),
            .I(N__21833));
    LocalMux I__2750 (
            .O(N__21833),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ));
    InMux I__2749 (
            .O(N__21830),
            .I(N__21827));
    LocalMux I__2748 (
            .O(N__21827),
            .I(N__21824));
    Odrv4 I__2747 (
            .O(N__21824),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_20 ));
    CascadeMux I__2746 (
            .O(N__21821),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_10_31_cascade_ ));
    InMux I__2745 (
            .O(N__21818),
            .I(N__21815));
    LocalMux I__2744 (
            .O(N__21815),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_11_31 ));
    InMux I__2743 (
            .O(N__21812),
            .I(N__21809));
    LocalMux I__2742 (
            .O(N__21809),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_9_31 ));
    InMux I__2741 (
            .O(N__21806),
            .I(N__21803));
    LocalMux I__2740 (
            .O(N__21803),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_8_31 ));
    CascadeMux I__2739 (
            .O(N__21800),
            .I(N__21797));
    InMux I__2738 (
            .O(N__21797),
            .I(N__21794));
    LocalMux I__2737 (
            .O(N__21794),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_16 ));
    InMux I__2736 (
            .O(N__21791),
            .I(N__21788));
    LocalMux I__2735 (
            .O(N__21788),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_21 ));
    CascadeMux I__2734 (
            .O(N__21785),
            .I(N__21782));
    InMux I__2733 (
            .O(N__21782),
            .I(N__21779));
    LocalMux I__2732 (
            .O(N__21779),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ));
    CascadeMux I__2731 (
            .O(N__21776),
            .I(N__21773));
    InMux I__2730 (
            .O(N__21773),
            .I(N__21770));
    LocalMux I__2729 (
            .O(N__21770),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ));
    CascadeMux I__2728 (
            .O(N__21767),
            .I(N__21764));
    InMux I__2727 (
            .O(N__21764),
            .I(N__21761));
    LocalMux I__2726 (
            .O(N__21761),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ));
    CascadeMux I__2725 (
            .O(N__21758),
            .I(N__21755));
    InMux I__2724 (
            .O(N__21755),
            .I(N__21752));
    LocalMux I__2723 (
            .O(N__21752),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ));
    InMux I__2722 (
            .O(N__21749),
            .I(N__21746));
    LocalMux I__2721 (
            .O(N__21746),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_15 ));
    CascadeMux I__2720 (
            .O(N__21743),
            .I(N__21740));
    InMux I__2719 (
            .O(N__21740),
            .I(N__21737));
    LocalMux I__2718 (
            .O(N__21737),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_19 ));
    CascadeMux I__2717 (
            .O(N__21734),
            .I(N__21731));
    InMux I__2716 (
            .O(N__21731),
            .I(N__21728));
    LocalMux I__2715 (
            .O(N__21728),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ));
    InMux I__2714 (
            .O(N__21725),
            .I(N__21722));
    LocalMux I__2713 (
            .O(N__21722),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ));
    InMux I__2712 (
            .O(N__21719),
            .I(N__21716));
    LocalMux I__2711 (
            .O(N__21716),
            .I(N__21708));
    InMux I__2710 (
            .O(N__21715),
            .I(N__21705));
    InMux I__2709 (
            .O(N__21714),
            .I(N__21702));
    InMux I__2708 (
            .O(N__21713),
            .I(N__21697));
    InMux I__2707 (
            .O(N__21712),
            .I(N__21697));
    InMux I__2706 (
            .O(N__21711),
            .I(N__21694));
    Span4Mux_v I__2705 (
            .O(N__21708),
            .I(N__21685));
    LocalMux I__2704 (
            .O(N__21705),
            .I(N__21685));
    LocalMux I__2703 (
            .O(N__21702),
            .I(N__21685));
    LocalMux I__2702 (
            .O(N__21697),
            .I(N__21685));
    LocalMux I__2701 (
            .O(N__21694),
            .I(un2_counter_8));
    Odrv4 I__2700 (
            .O(N__21685),
            .I(un2_counter_8));
    InMux I__2699 (
            .O(N__21680),
            .I(N__21677));
    LocalMux I__2698 (
            .O(N__21677),
            .I(counter_RNO_0Z0Z_10));
    CascadeMux I__2697 (
            .O(N__21674),
            .I(N__21671));
    InMux I__2696 (
            .O(N__21671),
            .I(N__21668));
    LocalMux I__2695 (
            .O(N__21668),
            .I(N__21662));
    InMux I__2694 (
            .O(N__21667),
            .I(N__21659));
    CascadeMux I__2693 (
            .O(N__21666),
            .I(N__21656));
    CascadeMux I__2692 (
            .O(N__21665),
            .I(N__21652));
    Span4Mux_h I__2691 (
            .O(N__21662),
            .I(N__21649));
    LocalMux I__2690 (
            .O(N__21659),
            .I(N__21646));
    InMux I__2689 (
            .O(N__21656),
            .I(N__21643));
    InMux I__2688 (
            .O(N__21655),
            .I(N__21638));
    InMux I__2687 (
            .O(N__21652),
            .I(N__21638));
    Odrv4 I__2686 (
            .O(N__21649),
            .I(un2_counter_9));
    Odrv4 I__2685 (
            .O(N__21646),
            .I(un2_counter_9));
    LocalMux I__2684 (
            .O(N__21643),
            .I(un2_counter_9));
    LocalMux I__2683 (
            .O(N__21638),
            .I(un2_counter_9));
    CascadeMux I__2682 (
            .O(N__21629),
            .I(N__21625));
    InMux I__2681 (
            .O(N__21628),
            .I(N__21622));
    InMux I__2680 (
            .O(N__21625),
            .I(N__21616));
    LocalMux I__2679 (
            .O(N__21622),
            .I(N__21613));
    InMux I__2678 (
            .O(N__21621),
            .I(N__21608));
    InMux I__2677 (
            .O(N__21620),
            .I(N__21608));
    InMux I__2676 (
            .O(N__21619),
            .I(N__21605));
    LocalMux I__2675 (
            .O(N__21616),
            .I(N__21598));
    Span4Mux_v I__2674 (
            .O(N__21613),
            .I(N__21598));
    LocalMux I__2673 (
            .O(N__21608),
            .I(N__21598));
    LocalMux I__2672 (
            .O(N__21605),
            .I(un2_counter_7));
    Odrv4 I__2671 (
            .O(N__21598),
            .I(un2_counter_7));
    InMux I__2670 (
            .O(N__21593),
            .I(N__21589));
    InMux I__2669 (
            .O(N__21592),
            .I(N__21586));
    LocalMux I__2668 (
            .O(N__21589),
            .I(counterZ0Z_10));
    LocalMux I__2667 (
            .O(N__21586),
            .I(counterZ0Z_10));
    InMux I__2666 (
            .O(N__21581),
            .I(N__21578));
    LocalMux I__2665 (
            .O(N__21578),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_8 ));
    CascadeMux I__2664 (
            .O(N__21575),
            .I(N__21572));
    InMux I__2663 (
            .O(N__21572),
            .I(N__21569));
    LocalMux I__2662 (
            .O(N__21569),
            .I(N__21566));
    Span4Mux_v I__2661 (
            .O(N__21566),
            .I(N__21563));
    Odrv4 I__2660 (
            .O(N__21563),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ));
    InMux I__2659 (
            .O(N__21560),
            .I(N__21557));
    LocalMux I__2658 (
            .O(N__21557),
            .I(N__21554));
    Odrv4 I__2657 (
            .O(N__21554),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ));
    CascadeMux I__2656 (
            .O(N__21551),
            .I(N__21548));
    InMux I__2655 (
            .O(N__21548),
            .I(N__21545));
    LocalMux I__2654 (
            .O(N__21545),
            .I(N__21542));
    Odrv4 I__2653 (
            .O(N__21542),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ));
    CascadeMux I__2652 (
            .O(N__21539),
            .I(N__21536));
    InMux I__2651 (
            .O(N__21536),
            .I(N__21533));
    LocalMux I__2650 (
            .O(N__21533),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ));
    CascadeMux I__2649 (
            .O(N__21530),
            .I(N__21527));
    InMux I__2648 (
            .O(N__21527),
            .I(N__21524));
    LocalMux I__2647 (
            .O(N__21524),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ));
    CascadeMux I__2646 (
            .O(N__21521),
            .I(N__21518));
    InMux I__2645 (
            .O(N__21518),
            .I(N__21515));
    LocalMux I__2644 (
            .O(N__21515),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ));
    CascadeMux I__2643 (
            .O(N__21512),
            .I(N__21509));
    InMux I__2642 (
            .O(N__21509),
            .I(N__21506));
    LocalMux I__2641 (
            .O(N__21506),
            .I(N__21503));
    Span4Mux_v I__2640 (
            .O(N__21503),
            .I(N__21500));
    Odrv4 I__2639 (
            .O(N__21500),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_17 ));
    CascadeMux I__2638 (
            .O(N__21497),
            .I(N__21494));
    InMux I__2637 (
            .O(N__21494),
            .I(N__21491));
    LocalMux I__2636 (
            .O(N__21491),
            .I(N__21488));
    Odrv12 I__2635 (
            .O(N__21488),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ));
    InMux I__2634 (
            .O(N__21485),
            .I(N__21482));
    LocalMux I__2633 (
            .O(N__21482),
            .I(counter_RNO_0Z0Z_7));
    InMux I__2632 (
            .O(N__21479),
            .I(N__21475));
    InMux I__2631 (
            .O(N__21478),
            .I(N__21472));
    LocalMux I__2630 (
            .O(N__21475),
            .I(counterZ0Z_7));
    LocalMux I__2629 (
            .O(N__21472),
            .I(counterZ0Z_7));
    CascadeMux I__2628 (
            .O(N__21467),
            .I(N__21462));
    InMux I__2627 (
            .O(N__21466),
            .I(N__21459));
    InMux I__2626 (
            .O(N__21465),
            .I(N__21456));
    InMux I__2625 (
            .O(N__21462),
            .I(N__21453));
    LocalMux I__2624 (
            .O(N__21459),
            .I(N__21448));
    LocalMux I__2623 (
            .O(N__21456),
            .I(N__21448));
    LocalMux I__2622 (
            .O(N__21453),
            .I(counterZ0Z_1));
    Odrv4 I__2621 (
            .O(N__21448),
            .I(counterZ0Z_1));
    InMux I__2620 (
            .O(N__21443),
            .I(N__21439));
    InMux I__2619 (
            .O(N__21442),
            .I(N__21436));
    LocalMux I__2618 (
            .O(N__21439),
            .I(counterZ0Z_2));
    LocalMux I__2617 (
            .O(N__21436),
            .I(counterZ0Z_2));
    CascadeMux I__2616 (
            .O(N__21431),
            .I(un2_counter_5_cascade_));
    InMux I__2615 (
            .O(N__21428),
            .I(N__21422));
    InMux I__2614 (
            .O(N__21427),
            .I(N__21417));
    InMux I__2613 (
            .O(N__21426),
            .I(N__21417));
    InMux I__2612 (
            .O(N__21425),
            .I(N__21414));
    LocalMux I__2611 (
            .O(N__21422),
            .I(N__21411));
    LocalMux I__2610 (
            .O(N__21417),
            .I(counterZ0Z_0));
    LocalMux I__2609 (
            .O(N__21414),
            .I(counterZ0Z_0));
    Odrv4 I__2608 (
            .O(N__21411),
            .I(counterZ0Z_0));
    CascadeMux I__2607 (
            .O(N__21404),
            .I(un2_counter_9_cascade_));
    CascadeMux I__2606 (
            .O(N__21401),
            .I(clk_10khz_RNIIENAZ0Z2_cascade_));
    InMux I__2605 (
            .O(N__21398),
            .I(N__21395));
    LocalMux I__2604 (
            .O(N__21395),
            .I(N__21392));
    Odrv4 I__2603 (
            .O(N__21392),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_2 ));
    InMux I__2602 (
            .O(N__21389),
            .I(N__21385));
    InMux I__2601 (
            .O(N__21388),
            .I(N__21382));
    LocalMux I__2600 (
            .O(N__21385),
            .I(N__21377));
    LocalMux I__2599 (
            .O(N__21382),
            .I(N__21377));
    Odrv4 I__2598 (
            .O(N__21377),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ));
    InMux I__2597 (
            .O(N__21374),
            .I(bfn_4_16_0_));
    InMux I__2596 (
            .O(N__21371),
            .I(N__21365));
    InMux I__2595 (
            .O(N__21370),
            .I(N__21365));
    LocalMux I__2594 (
            .O(N__21365),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ));
    InMux I__2593 (
            .O(N__21362),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ));
    InMux I__2592 (
            .O(N__21359),
            .I(N__21355));
    CascadeMux I__2591 (
            .O(N__21358),
            .I(N__21352));
    LocalMux I__2590 (
            .O(N__21355),
            .I(N__21349));
    InMux I__2589 (
            .O(N__21352),
            .I(N__21346));
    Span4Mux_v I__2588 (
            .O(N__21349),
            .I(N__21343));
    LocalMux I__2587 (
            .O(N__21346),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ));
    Odrv4 I__2586 (
            .O(N__21343),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ));
    InMux I__2585 (
            .O(N__21338),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ));
    InMux I__2584 (
            .O(N__21335),
            .I(N__21331));
    InMux I__2583 (
            .O(N__21334),
            .I(N__21328));
    LocalMux I__2582 (
            .O(N__21331),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    LocalMux I__2581 (
            .O(N__21328),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    InMux I__2580 (
            .O(N__21323),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ));
    InMux I__2579 (
            .O(N__21320),
            .I(N__21316));
    InMux I__2578 (
            .O(N__21319),
            .I(N__21313));
    LocalMux I__2577 (
            .O(N__21316),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    LocalMux I__2576 (
            .O(N__21313),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    InMux I__2575 (
            .O(N__21308),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ));
    InMux I__2574 (
            .O(N__21305),
            .I(N__21301));
    InMux I__2573 (
            .O(N__21304),
            .I(N__21298));
    LocalMux I__2572 (
            .O(N__21301),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    LocalMux I__2571 (
            .O(N__21298),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    InMux I__2570 (
            .O(N__21293),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ));
    CascadeMux I__2569 (
            .O(N__21290),
            .I(N__21286));
    InMux I__2568 (
            .O(N__21289),
            .I(N__21283));
    InMux I__2567 (
            .O(N__21286),
            .I(N__21280));
    LocalMux I__2566 (
            .O(N__21283),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    LocalMux I__2565 (
            .O(N__21280),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    InMux I__2564 (
            .O(N__21275),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ));
    InMux I__2563 (
            .O(N__21272),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ));
    InMux I__2562 (
            .O(N__21269),
            .I(N__21262));
    CascadeMux I__2561 (
            .O(N__21268),
            .I(N__21259));
    CascadeMux I__2560 (
            .O(N__21267),
            .I(N__21254));
    CascadeMux I__2559 (
            .O(N__21266),
            .I(N__21250));
    CascadeMux I__2558 (
            .O(N__21265),
            .I(N__21247));
    LocalMux I__2557 (
            .O(N__21262),
            .I(N__21242));
    InMux I__2556 (
            .O(N__21259),
            .I(N__21237));
    InMux I__2555 (
            .O(N__21258),
            .I(N__21237));
    InMux I__2554 (
            .O(N__21257),
            .I(N__21226));
    InMux I__2553 (
            .O(N__21254),
            .I(N__21226));
    InMux I__2552 (
            .O(N__21253),
            .I(N__21226));
    InMux I__2551 (
            .O(N__21250),
            .I(N__21226));
    InMux I__2550 (
            .O(N__21247),
            .I(N__21226));
    InMux I__2549 (
            .O(N__21246),
            .I(N__21223));
    InMux I__2548 (
            .O(N__21245),
            .I(N__21220));
    Span4Mux_h I__2547 (
            .O(N__21242),
            .I(N__21217));
    LocalMux I__2546 (
            .O(N__21237),
            .I(N__21214));
    LocalMux I__2545 (
            .O(N__21226),
            .I(N__21207));
    LocalMux I__2544 (
            .O(N__21223),
            .I(N__21207));
    LocalMux I__2543 (
            .O(N__21220),
            .I(N__21207));
    Span4Mux_v I__2542 (
            .O(N__21217),
            .I(N__21204));
    Span4Mux_v I__2541 (
            .O(N__21214),
            .I(N__21201));
    Span12Mux_v I__2540 (
            .O(N__21207),
            .I(N__21198));
    Span4Mux_v I__2539 (
            .O(N__21204),
            .I(N__21195));
    Span4Mux_v I__2538 (
            .O(N__21201),
            .I(N__21192));
    Odrv12 I__2537 (
            .O(N__21198),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    Odrv4 I__2536 (
            .O(N__21195),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    Odrv4 I__2535 (
            .O(N__21192),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    InMux I__2534 (
            .O(N__21185),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ));
    CascadeMux I__2533 (
            .O(N__21182),
            .I(N__21179));
    InMux I__2532 (
            .O(N__21179),
            .I(N__21173));
    InMux I__2531 (
            .O(N__21178),
            .I(N__21173));
    LocalMux I__2530 (
            .O(N__21173),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    InMux I__2529 (
            .O(N__21170),
            .I(bfn_4_15_0_));
    InMux I__2528 (
            .O(N__21167),
            .I(N__21161));
    InMux I__2527 (
            .O(N__21166),
            .I(N__21161));
    LocalMux I__2526 (
            .O(N__21161),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    InMux I__2525 (
            .O(N__21158),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ));
    CascadeMux I__2524 (
            .O(N__21155),
            .I(N__21151));
    InMux I__2523 (
            .O(N__21154),
            .I(N__21146));
    InMux I__2522 (
            .O(N__21151),
            .I(N__21146));
    LocalMux I__2521 (
            .O(N__21146),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    InMux I__2520 (
            .O(N__21143),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ));
    CascadeMux I__2519 (
            .O(N__21140),
            .I(N__21137));
    InMux I__2518 (
            .O(N__21137),
            .I(N__21133));
    InMux I__2517 (
            .O(N__21136),
            .I(N__21130));
    LocalMux I__2516 (
            .O(N__21133),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    LocalMux I__2515 (
            .O(N__21130),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    InMux I__2514 (
            .O(N__21125),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ));
    InMux I__2513 (
            .O(N__21122),
            .I(N__21118));
    InMux I__2512 (
            .O(N__21121),
            .I(N__21115));
    LocalMux I__2511 (
            .O(N__21118),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    LocalMux I__2510 (
            .O(N__21115),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    InMux I__2509 (
            .O(N__21110),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ));
    InMux I__2508 (
            .O(N__21107),
            .I(N__21101));
    InMux I__2507 (
            .O(N__21106),
            .I(N__21101));
    LocalMux I__2506 (
            .O(N__21101),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    InMux I__2505 (
            .O(N__21098),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ));
    CascadeMux I__2504 (
            .O(N__21095),
            .I(N__21091));
    CascadeMux I__2503 (
            .O(N__21094),
            .I(N__21088));
    InMux I__2502 (
            .O(N__21091),
            .I(N__21083));
    InMux I__2501 (
            .O(N__21088),
            .I(N__21083));
    LocalMux I__2500 (
            .O(N__21083),
            .I(N__21080));
    Odrv4 I__2499 (
            .O(N__21080),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    InMux I__2498 (
            .O(N__21077),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ));
    InMux I__2497 (
            .O(N__21074),
            .I(N__21068));
    InMux I__2496 (
            .O(N__21073),
            .I(N__21068));
    LocalMux I__2495 (
            .O(N__21068),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ));
    InMux I__2494 (
            .O(N__21065),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ));
    InMux I__2493 (
            .O(N__21062),
            .I(N__21058));
    InMux I__2492 (
            .O(N__21061),
            .I(N__21054));
    LocalMux I__2491 (
            .O(N__21058),
            .I(N__21051));
    InMux I__2490 (
            .O(N__21057),
            .I(N__21048));
    LocalMux I__2489 (
            .O(N__21054),
            .I(N__21045));
    Span12Mux_v I__2488 (
            .O(N__21051),
            .I(N__21042));
    LocalMux I__2487 (
            .O(N__21048),
            .I(N__21037));
    Span4Mux_h I__2486 (
            .O(N__21045),
            .I(N__21037));
    Odrv12 I__2485 (
            .O(N__21042),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    Odrv4 I__2484 (
            .O(N__21037),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    InMux I__2483 (
            .O(N__21032),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ));
    InMux I__2482 (
            .O(N__21029),
            .I(N__21026));
    LocalMux I__2481 (
            .O(N__21026),
            .I(N__21021));
    CascadeMux I__2480 (
            .O(N__21025),
            .I(N__21018));
    InMux I__2479 (
            .O(N__21024),
            .I(N__21015));
    Span4Mux_v I__2478 (
            .O(N__21021),
            .I(N__21012));
    InMux I__2477 (
            .O(N__21018),
            .I(N__21009));
    LocalMux I__2476 (
            .O(N__21015),
            .I(N__21006));
    Span4Mux_v I__2475 (
            .O(N__21012),
            .I(N__21001));
    LocalMux I__2474 (
            .O(N__21009),
            .I(N__21001));
    Span4Mux_h I__2473 (
            .O(N__21006),
            .I(N__20998));
    Span4Mux_h I__2472 (
            .O(N__21001),
            .I(N__20995));
    Odrv4 I__2471 (
            .O(N__20998),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    Odrv4 I__2470 (
            .O(N__20995),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    InMux I__2469 (
            .O(N__20990),
            .I(bfn_4_14_0_));
    InMux I__2468 (
            .O(N__20987),
            .I(N__20984));
    LocalMux I__2467 (
            .O(N__20984),
            .I(N__20981));
    Span4Mux_v I__2466 (
            .O(N__20981),
            .I(N__20977));
    InMux I__2465 (
            .O(N__20980),
            .I(N__20973));
    Span4Mux_v I__2464 (
            .O(N__20977),
            .I(N__20970));
    InMux I__2463 (
            .O(N__20976),
            .I(N__20967));
    LocalMux I__2462 (
            .O(N__20973),
            .I(N__20964));
    Span4Mux_h I__2461 (
            .O(N__20970),
            .I(N__20961));
    LocalMux I__2460 (
            .O(N__20967),
            .I(N__20956));
    Span4Mux_h I__2459 (
            .O(N__20964),
            .I(N__20956));
    Odrv4 I__2458 (
            .O(N__20961),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    Odrv4 I__2457 (
            .O(N__20956),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    InMux I__2456 (
            .O(N__20951),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ));
    InMux I__2455 (
            .O(N__20948),
            .I(N__20942));
    InMux I__2454 (
            .O(N__20947),
            .I(N__20942));
    LocalMux I__2453 (
            .O(N__20942),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ));
    InMux I__2452 (
            .O(N__20939),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ));
    InMux I__2451 (
            .O(N__20936),
            .I(N__20930));
    InMux I__2450 (
            .O(N__20935),
            .I(N__20930));
    LocalMux I__2449 (
            .O(N__20930),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ));
    InMux I__2448 (
            .O(N__20927),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ));
    InMux I__2447 (
            .O(N__20924),
            .I(N__20921));
    LocalMux I__2446 (
            .O(N__20921),
            .I(N__20917));
    InMux I__2445 (
            .O(N__20920),
            .I(N__20914));
    Odrv4 I__2444 (
            .O(N__20917),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    LocalMux I__2443 (
            .O(N__20914),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    InMux I__2442 (
            .O(N__20909),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ));
    InMux I__2441 (
            .O(N__20906),
            .I(N__20900));
    InMux I__2440 (
            .O(N__20905),
            .I(N__20900));
    LocalMux I__2439 (
            .O(N__20900),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    InMux I__2438 (
            .O(N__20897),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ));
    CascadeMux I__2437 (
            .O(N__20894),
            .I(N__20891));
    InMux I__2436 (
            .O(N__20891),
            .I(N__20888));
    LocalMux I__2435 (
            .O(N__20888),
            .I(N__20884));
    InMux I__2434 (
            .O(N__20887),
            .I(N__20881));
    Odrv4 I__2433 (
            .O(N__20884),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    LocalMux I__2432 (
            .O(N__20881),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    InMux I__2431 (
            .O(N__20876),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ));
    InMux I__2430 (
            .O(N__20873),
            .I(N__20869));
    InMux I__2429 (
            .O(N__20872),
            .I(N__20866));
    LocalMux I__2428 (
            .O(N__20869),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    LocalMux I__2427 (
            .O(N__20866),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    CascadeMux I__2426 (
            .O(N__20861),
            .I(N__20851));
    CascadeMux I__2425 (
            .O(N__20860),
            .I(N__20848));
    CascadeMux I__2424 (
            .O(N__20859),
            .I(N__20843));
    CascadeMux I__2423 (
            .O(N__20858),
            .I(N__20840));
    InMux I__2422 (
            .O(N__20857),
            .I(N__20833));
    InMux I__2421 (
            .O(N__20856),
            .I(N__20833));
    InMux I__2420 (
            .O(N__20855),
            .I(N__20833));
    InMux I__2419 (
            .O(N__20854),
            .I(N__20830));
    InMux I__2418 (
            .O(N__20851),
            .I(N__20825));
    InMux I__2417 (
            .O(N__20848),
            .I(N__20825));
    InMux I__2416 (
            .O(N__20847),
            .I(N__20820));
    InMux I__2415 (
            .O(N__20846),
            .I(N__20820));
    InMux I__2414 (
            .O(N__20843),
            .I(N__20815));
    InMux I__2413 (
            .O(N__20840),
            .I(N__20815));
    LocalMux I__2412 (
            .O(N__20833),
            .I(N__20812));
    LocalMux I__2411 (
            .O(N__20830),
            .I(N__20808));
    LocalMux I__2410 (
            .O(N__20825),
            .I(N__20803));
    LocalMux I__2409 (
            .O(N__20820),
            .I(N__20803));
    LocalMux I__2408 (
            .O(N__20815),
            .I(N__20798));
    Span4Mux_v I__2407 (
            .O(N__20812),
            .I(N__20798));
    InMux I__2406 (
            .O(N__20811),
            .I(N__20795));
    Span4Mux_v I__2405 (
            .O(N__20808),
            .I(N__20792));
    Span12Mux_h I__2404 (
            .O(N__20803),
            .I(N__20789));
    Span4Mux_h I__2403 (
            .O(N__20798),
            .I(N__20784));
    LocalMux I__2402 (
            .O(N__20795),
            .I(N__20784));
    Odrv4 I__2401 (
            .O(N__20792),
            .I(pwm_duty_input_6));
    Odrv12 I__2400 (
            .O(N__20789),
            .I(pwm_duty_input_6));
    Odrv4 I__2399 (
            .O(N__20784),
            .I(pwm_duty_input_6));
    InMux I__2398 (
            .O(N__20777),
            .I(N__20763));
    InMux I__2397 (
            .O(N__20776),
            .I(N__20763));
    InMux I__2396 (
            .O(N__20775),
            .I(N__20754));
    InMux I__2395 (
            .O(N__20774),
            .I(N__20754));
    InMux I__2394 (
            .O(N__20773),
            .I(N__20754));
    InMux I__2393 (
            .O(N__20772),
            .I(N__20754));
    InMux I__2392 (
            .O(N__20771),
            .I(N__20747));
    InMux I__2391 (
            .O(N__20770),
            .I(N__20747));
    InMux I__2390 (
            .O(N__20769),
            .I(N__20747));
    InMux I__2389 (
            .O(N__20768),
            .I(N__20744));
    LocalMux I__2388 (
            .O(N__20763),
            .I(N__20737));
    LocalMux I__2387 (
            .O(N__20754),
            .I(N__20737));
    LocalMux I__2386 (
            .O(N__20747),
            .I(N__20737));
    LocalMux I__2385 (
            .O(N__20744),
            .I(N__20734));
    Span4Mux_v I__2384 (
            .O(N__20737),
            .I(N__20731));
    Odrv12 I__2383 (
            .O(N__20734),
            .I(N_28_mux));
    Odrv4 I__2382 (
            .O(N__20731),
            .I(N_28_mux));
    CascadeMux I__2381 (
            .O(N__20726),
            .I(N__20716));
    CascadeMux I__2380 (
            .O(N__20725),
            .I(N__20713));
    CascadeMux I__2379 (
            .O(N__20724),
            .I(N__20709));
    CascadeMux I__2378 (
            .O(N__20723),
            .I(N__20706));
    CascadeMux I__2377 (
            .O(N__20722),
            .I(N__20703));
    InMux I__2376 (
            .O(N__20721),
            .I(N__20697));
    InMux I__2375 (
            .O(N__20720),
            .I(N__20697));
    InMux I__2374 (
            .O(N__20719),
            .I(N__20688));
    InMux I__2373 (
            .O(N__20716),
            .I(N__20688));
    InMux I__2372 (
            .O(N__20713),
            .I(N__20688));
    InMux I__2371 (
            .O(N__20712),
            .I(N__20688));
    InMux I__2370 (
            .O(N__20709),
            .I(N__20685));
    InMux I__2369 (
            .O(N__20706),
            .I(N__20680));
    InMux I__2368 (
            .O(N__20703),
            .I(N__20680));
    InMux I__2367 (
            .O(N__20702),
            .I(N__20677));
    LocalMux I__2366 (
            .O(N__20697),
            .I(N__20668));
    LocalMux I__2365 (
            .O(N__20688),
            .I(N__20668));
    LocalMux I__2364 (
            .O(N__20685),
            .I(N__20668));
    LocalMux I__2363 (
            .O(N__20680),
            .I(N__20668));
    LocalMux I__2362 (
            .O(N__20677),
            .I(N__20665));
    Span4Mux_v I__2361 (
            .O(N__20668),
            .I(N__20662));
    Odrv12 I__2360 (
            .O(N__20665),
            .I(i8_mux));
    Odrv4 I__2359 (
            .O(N__20662),
            .I(i8_mux));
    InMux I__2358 (
            .O(N__20657),
            .I(N__20654));
    LocalMux I__2357 (
            .O(N__20654),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8 ));
    CascadeMux I__2356 (
            .O(N__20651),
            .I(N__20648));
    InMux I__2355 (
            .O(N__20648),
            .I(N__20645));
    LocalMux I__2354 (
            .O(N__20645),
            .I(N__20642));
    Span4Mux_h I__2353 (
            .O(N__20642),
            .I(N__20639));
    Span4Mux_v I__2352 (
            .O(N__20639),
            .I(N__20636));
    Odrv4 I__2351 (
            .O(N__20636),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ));
    InMux I__2350 (
            .O(N__20633),
            .I(N__20630));
    LocalMux I__2349 (
            .O(N__20630),
            .I(N__20627));
    Span4Mux_h I__2348 (
            .O(N__20627),
            .I(N__20624));
    Span4Mux_v I__2347 (
            .O(N__20624),
            .I(N__20621));
    Odrv4 I__2346 (
            .O(N__20621),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ));
    InMux I__2345 (
            .O(N__20618),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ));
    CascadeMux I__2344 (
            .O(N__20615),
            .I(N__20612));
    InMux I__2343 (
            .O(N__20612),
            .I(N__20609));
    LocalMux I__2342 (
            .O(N__20609),
            .I(N__20606));
    Span4Mux_v I__2341 (
            .O(N__20606),
            .I(N__20603));
    Span4Mux_h I__2340 (
            .O(N__20603),
            .I(N__20600));
    Odrv4 I__2339 (
            .O(N__20600),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ));
    InMux I__2338 (
            .O(N__20597),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ));
    CascadeMux I__2337 (
            .O(N__20594),
            .I(N__20591));
    InMux I__2336 (
            .O(N__20591),
            .I(N__20587));
    InMux I__2335 (
            .O(N__20590),
            .I(N__20584));
    LocalMux I__2334 (
            .O(N__20587),
            .I(N__20580));
    LocalMux I__2333 (
            .O(N__20584),
            .I(N__20577));
    InMux I__2332 (
            .O(N__20583),
            .I(N__20574));
    Span4Mux_h I__2331 (
            .O(N__20580),
            .I(N__20569));
    Span4Mux_h I__2330 (
            .O(N__20577),
            .I(N__20569));
    LocalMux I__2329 (
            .O(N__20574),
            .I(N__20566));
    Span4Mux_v I__2328 (
            .O(N__20569),
            .I(N__20563));
    Span4Mux_v I__2327 (
            .O(N__20566),
            .I(N__20560));
    Odrv4 I__2326 (
            .O(N__20563),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    Odrv4 I__2325 (
            .O(N__20560),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    InMux I__2324 (
            .O(N__20555),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ));
    CascadeMux I__2323 (
            .O(N__20552),
            .I(N__20549));
    InMux I__2322 (
            .O(N__20549),
            .I(N__20545));
    InMux I__2321 (
            .O(N__20548),
            .I(N__20542));
    LocalMux I__2320 (
            .O(N__20545),
            .I(N__20537));
    LocalMux I__2319 (
            .O(N__20542),
            .I(N__20534));
    InMux I__2318 (
            .O(N__20541),
            .I(N__20531));
    InMux I__2317 (
            .O(N__20540),
            .I(N__20528));
    Span4Mux_v I__2316 (
            .O(N__20537),
            .I(N__20523));
    Span4Mux_v I__2315 (
            .O(N__20534),
            .I(N__20523));
    LocalMux I__2314 (
            .O(N__20531),
            .I(N__20520));
    LocalMux I__2313 (
            .O(N__20528),
            .I(N__20517));
    Span4Mux_v I__2312 (
            .O(N__20523),
            .I(N__20514));
    Span4Mux_v I__2311 (
            .O(N__20520),
            .I(N__20509));
    Span4Mux_v I__2310 (
            .O(N__20517),
            .I(N__20509));
    Odrv4 I__2309 (
            .O(N__20514),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    Odrv4 I__2308 (
            .O(N__20509),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    InMux I__2307 (
            .O(N__20504),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ));
    InMux I__2306 (
            .O(N__20501),
            .I(N__20498));
    LocalMux I__2305 (
            .O(N__20498),
            .I(N__20495));
    Span4Mux_h I__2304 (
            .O(N__20495),
            .I(N__20490));
    InMux I__2303 (
            .O(N__20494),
            .I(N__20487));
    InMux I__2302 (
            .O(N__20493),
            .I(N__20484));
    Span4Mux_v I__2301 (
            .O(N__20490),
            .I(N__20477));
    LocalMux I__2300 (
            .O(N__20487),
            .I(N__20477));
    LocalMux I__2299 (
            .O(N__20484),
            .I(N__20477));
    Odrv4 I__2298 (
            .O(N__20477),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    InMux I__2297 (
            .O(N__20474),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ));
    InMux I__2296 (
            .O(N__20471),
            .I(N__20468));
    LocalMux I__2295 (
            .O(N__20468),
            .I(N__20464));
    InMux I__2294 (
            .O(N__20467),
            .I(N__20460));
    Span4Mux_h I__2293 (
            .O(N__20464),
            .I(N__20457));
    InMux I__2292 (
            .O(N__20463),
            .I(N__20454));
    LocalMux I__2291 (
            .O(N__20460),
            .I(N__20451));
    Sp12to4 I__2290 (
            .O(N__20457),
            .I(N__20448));
    LocalMux I__2289 (
            .O(N__20454),
            .I(N__20443));
    Span4Mux_h I__2288 (
            .O(N__20451),
            .I(N__20443));
    Odrv12 I__2287 (
            .O(N__20448),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    Odrv4 I__2286 (
            .O(N__20443),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    InMux I__2285 (
            .O(N__20438),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ));
    InMux I__2284 (
            .O(N__20435),
            .I(un5_counter_cry_9));
    InMux I__2283 (
            .O(N__20432),
            .I(N__20428));
    InMux I__2282 (
            .O(N__20431),
            .I(N__20425));
    LocalMux I__2281 (
            .O(N__20428),
            .I(counterZ0Z_11));
    LocalMux I__2280 (
            .O(N__20425),
            .I(counterZ0Z_11));
    InMux I__2279 (
            .O(N__20420),
            .I(un5_counter_cry_10));
    InMux I__2278 (
            .O(N__20417),
            .I(N__20413));
    InMux I__2277 (
            .O(N__20416),
            .I(N__20410));
    LocalMux I__2276 (
            .O(N__20413),
            .I(counterZ0Z_12));
    LocalMux I__2275 (
            .O(N__20410),
            .I(counterZ0Z_12));
    InMux I__2274 (
            .O(N__20405),
            .I(un5_counter_cry_11));
    InMux I__2273 (
            .O(N__20402),
            .I(N__20399));
    LocalMux I__2272 (
            .O(N__20399),
            .I(counter_RNO_0Z0Z_12));
    InMux I__2271 (
            .O(N__20396),
            .I(N__20393));
    LocalMux I__2270 (
            .O(N__20393),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0 ));
    InMux I__2269 (
            .O(N__20390),
            .I(N__20387));
    LocalMux I__2268 (
            .O(N__20387),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4 ));
    InMux I__2267 (
            .O(N__20384),
            .I(N__20381));
    LocalMux I__2266 (
            .O(N__20381),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1 ));
    InMux I__2265 (
            .O(N__20378),
            .I(N__20375));
    LocalMux I__2264 (
            .O(N__20375),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3 ));
    InMux I__2263 (
            .O(N__20372),
            .I(N__20369));
    LocalMux I__2262 (
            .O(N__20369),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6 ));
    InMux I__2261 (
            .O(N__20366),
            .I(N__20363));
    LocalMux I__2260 (
            .O(N__20363),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5 ));
    InMux I__2259 (
            .O(N__20360),
            .I(un5_counter_cry_1));
    InMux I__2258 (
            .O(N__20357),
            .I(N__20353));
    InMux I__2257 (
            .O(N__20356),
            .I(N__20350));
    LocalMux I__2256 (
            .O(N__20353),
            .I(counterZ0Z_3));
    LocalMux I__2255 (
            .O(N__20350),
            .I(counterZ0Z_3));
    InMux I__2254 (
            .O(N__20345),
            .I(un5_counter_cry_2));
    InMux I__2253 (
            .O(N__20342),
            .I(N__20338));
    InMux I__2252 (
            .O(N__20341),
            .I(N__20335));
    LocalMux I__2251 (
            .O(N__20338),
            .I(counterZ0Z_4));
    LocalMux I__2250 (
            .O(N__20335),
            .I(counterZ0Z_4));
    InMux I__2249 (
            .O(N__20330),
            .I(un5_counter_cry_3));
    InMux I__2248 (
            .O(N__20327),
            .I(N__20323));
    InMux I__2247 (
            .O(N__20326),
            .I(N__20320));
    LocalMux I__2246 (
            .O(N__20323),
            .I(counterZ0Z_5));
    LocalMux I__2245 (
            .O(N__20320),
            .I(counterZ0Z_5));
    InMux I__2244 (
            .O(N__20315),
            .I(un5_counter_cry_4));
    CascadeMux I__2243 (
            .O(N__20312),
            .I(N__20308));
    InMux I__2242 (
            .O(N__20311),
            .I(N__20305));
    InMux I__2241 (
            .O(N__20308),
            .I(N__20302));
    LocalMux I__2240 (
            .O(N__20305),
            .I(counterZ0Z_6));
    LocalMux I__2239 (
            .O(N__20302),
            .I(counterZ0Z_6));
    InMux I__2238 (
            .O(N__20297),
            .I(un5_counter_cry_5));
    InMux I__2237 (
            .O(N__20294),
            .I(un5_counter_cry_6));
    CascadeMux I__2236 (
            .O(N__20291),
            .I(N__20287));
    InMux I__2235 (
            .O(N__20290),
            .I(N__20284));
    InMux I__2234 (
            .O(N__20287),
            .I(N__20281));
    LocalMux I__2233 (
            .O(N__20284),
            .I(counterZ0Z_8));
    LocalMux I__2232 (
            .O(N__20281),
            .I(counterZ0Z_8));
    InMux I__2231 (
            .O(N__20276),
            .I(un5_counter_cry_7));
    InMux I__2230 (
            .O(N__20273),
            .I(N__20269));
    InMux I__2229 (
            .O(N__20272),
            .I(N__20266));
    LocalMux I__2228 (
            .O(N__20269),
            .I(counterZ0Z_9));
    LocalMux I__2227 (
            .O(N__20266),
            .I(counterZ0Z_9));
    InMux I__2226 (
            .O(N__20261),
            .I(bfn_4_8_0_));
    InMux I__2225 (
            .O(N__20258),
            .I(N__20255));
    LocalMux I__2224 (
            .O(N__20255),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ));
    CascadeMux I__2223 (
            .O(N__20252),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_ ));
    InMux I__2222 (
            .O(N__20249),
            .I(N__20246));
    LocalMux I__2221 (
            .O(N__20246),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9 ));
    InMux I__2220 (
            .O(N__20243),
            .I(N__20240));
    LocalMux I__2219 (
            .O(N__20240),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ));
    InMux I__2218 (
            .O(N__20237),
            .I(N__20234));
    LocalMux I__2217 (
            .O(N__20234),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ));
    CascadeMux I__2216 (
            .O(N__20231),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_ ));
    InMux I__2215 (
            .O(N__20228),
            .I(N__20225));
    LocalMux I__2214 (
            .O(N__20225),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ));
    InMux I__2213 (
            .O(N__20222),
            .I(N__20219));
    LocalMux I__2212 (
            .O(N__20219),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ));
    InMux I__2211 (
            .O(N__20216),
            .I(N__20213));
    LocalMux I__2210 (
            .O(N__20213),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9 ));
    InMux I__2209 (
            .O(N__20210),
            .I(N__20207));
    LocalMux I__2208 (
            .O(N__20207),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ));
    InMux I__2207 (
            .O(N__20204),
            .I(N__20201));
    LocalMux I__2206 (
            .O(N__20201),
            .I(N__20198));
    Span4Mux_h I__2205 (
            .O(N__20198),
            .I(N__20194));
    InMux I__2204 (
            .O(N__20197),
            .I(N__20191));
    Odrv4 I__2203 (
            .O(N__20194),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ));
    LocalMux I__2202 (
            .O(N__20191),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ));
    InMux I__2201 (
            .O(N__20186),
            .I(N__20183));
    LocalMux I__2200 (
            .O(N__20183),
            .I(N__20179));
    InMux I__2199 (
            .O(N__20182),
            .I(N__20175));
    Span4Mux_h I__2198 (
            .O(N__20179),
            .I(N__20172));
    InMux I__2197 (
            .O(N__20178),
            .I(N__20169));
    LocalMux I__2196 (
            .O(N__20175),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ));
    Odrv4 I__2195 (
            .O(N__20172),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ));
    LocalMux I__2194 (
            .O(N__20169),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ));
    CascadeMux I__2193 (
            .O(N__20162),
            .I(N__20159));
    InMux I__2192 (
            .O(N__20159),
            .I(N__20156));
    LocalMux I__2191 (
            .O(N__20156),
            .I(N__20153));
    Odrv4 I__2190 (
            .O(N__20153),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO ));
    CascadeMux I__2189 (
            .O(N__20150),
            .I(N__20146));
    InMux I__2188 (
            .O(N__20149),
            .I(N__20143));
    InMux I__2187 (
            .O(N__20146),
            .I(N__20140));
    LocalMux I__2186 (
            .O(N__20143),
            .I(N__20127));
    LocalMux I__2185 (
            .O(N__20140),
            .I(N__20127));
    InMux I__2184 (
            .O(N__20139),
            .I(N__20122));
    InMux I__2183 (
            .O(N__20138),
            .I(N__20122));
    InMux I__2182 (
            .O(N__20137),
            .I(N__20111));
    InMux I__2181 (
            .O(N__20136),
            .I(N__20111));
    InMux I__2180 (
            .O(N__20135),
            .I(N__20111));
    InMux I__2179 (
            .O(N__20134),
            .I(N__20111));
    InMux I__2178 (
            .O(N__20133),
            .I(N__20111));
    InMux I__2177 (
            .O(N__20132),
            .I(N__20108));
    Span4Mux_v I__2176 (
            .O(N__20127),
            .I(N__20105));
    LocalMux I__2175 (
            .O(N__20122),
            .I(N__20102));
    LocalMux I__2174 (
            .O(N__20111),
            .I(N__20098));
    LocalMux I__2173 (
            .O(N__20108),
            .I(N__20095));
    Span4Mux_v I__2172 (
            .O(N__20105),
            .I(N__20091));
    Span4Mux_h I__2171 (
            .O(N__20102),
            .I(N__20088));
    InMux I__2170 (
            .O(N__20101),
            .I(N__20085));
    Span4Mux_v I__2169 (
            .O(N__20098),
            .I(N__20080));
    Span4Mux_v I__2168 (
            .O(N__20095),
            .I(N__20080));
    InMux I__2167 (
            .O(N__20094),
            .I(N__20077));
    Odrv4 I__2166 (
            .O(N__20091),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    Odrv4 I__2165 (
            .O(N__20088),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    LocalMux I__2164 (
            .O(N__20085),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    Odrv4 I__2163 (
            .O(N__20080),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    LocalMux I__2162 (
            .O(N__20077),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    InMux I__2161 (
            .O(N__20066),
            .I(N__20063));
    LocalMux I__2160 (
            .O(N__20063),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_4 ));
    CascadeMux I__2159 (
            .O(N__20060),
            .I(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ));
    InMux I__2158 (
            .O(N__20057),
            .I(N__20052));
    InMux I__2157 (
            .O(N__20056),
            .I(N__20049));
    InMux I__2156 (
            .O(N__20055),
            .I(N__20046));
    LocalMux I__2155 (
            .O(N__20052),
            .I(N__20043));
    LocalMux I__2154 (
            .O(N__20049),
            .I(N__20038));
    LocalMux I__2153 (
            .O(N__20046),
            .I(N__20038));
    Span4Mux_v I__2152 (
            .O(N__20043),
            .I(N__20035));
    Span4Mux_v I__2151 (
            .O(N__20038),
            .I(N__20032));
    Odrv4 I__2150 (
            .O(N__20035),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    Odrv4 I__2149 (
            .O(N__20032),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    CascadeMux I__2148 (
            .O(N__20027),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_9_9_cascade_ ));
    CascadeMux I__2147 (
            .O(N__20024),
            .I(N__20021));
    InMux I__2146 (
            .O(N__20021),
            .I(N__20018));
    LocalMux I__2145 (
            .O(N__20018),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ));
    InMux I__2144 (
            .O(N__20015),
            .I(N__20012));
    LocalMux I__2143 (
            .O(N__20012),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ));
    CascadeMux I__2142 (
            .O(N__20009),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9_cascade_ ));
    InMux I__2141 (
            .O(N__20006),
            .I(N__19997));
    InMux I__2140 (
            .O(N__20005),
            .I(N__19986));
    InMux I__2139 (
            .O(N__20004),
            .I(N__19986));
    InMux I__2138 (
            .O(N__20003),
            .I(N__19986));
    InMux I__2137 (
            .O(N__20002),
            .I(N__19986));
    InMux I__2136 (
            .O(N__20001),
            .I(N__19986));
    InMux I__2135 (
            .O(N__20000),
            .I(N__19983));
    LocalMux I__2134 (
            .O(N__19997),
            .I(N__19978));
    LocalMux I__2133 (
            .O(N__19986),
            .I(N__19978));
    LocalMux I__2132 (
            .O(N__19983),
            .I(N__19975));
    Span12Mux_v I__2131 (
            .O(N__19978),
            .I(N__19972));
    Span12Mux_s7_v I__2130 (
            .O(N__19975),
            .I(N__19969));
    Odrv12 I__2129 (
            .O(N__19972),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    Odrv12 I__2128 (
            .O(N__19969),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    InMux I__2127 (
            .O(N__19964),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_3 ));
    InMux I__2126 (
            .O(N__19961),
            .I(N__19958));
    LocalMux I__2125 (
            .O(N__19958),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_5 ));
    InMux I__2124 (
            .O(N__19955),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_4 ));
    InMux I__2123 (
            .O(N__19952),
            .I(N__19949));
    LocalMux I__2122 (
            .O(N__19949),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_6 ));
    InMux I__2121 (
            .O(N__19946),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_5 ));
    InMux I__2120 (
            .O(N__19943),
            .I(N__19940));
    LocalMux I__2119 (
            .O(N__19940),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_7 ));
    InMux I__2118 (
            .O(N__19937),
            .I(N__19934));
    LocalMux I__2117 (
            .O(N__19934),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7 ));
    InMux I__2116 (
            .O(N__19931),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_6 ));
    CascadeMux I__2115 (
            .O(N__19928),
            .I(N__19925));
    InMux I__2114 (
            .O(N__19925),
            .I(N__19922));
    LocalMux I__2113 (
            .O(N__19922),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_8 ));
    InMux I__2112 (
            .O(N__19919),
            .I(bfn_3_10_0_));
    InMux I__2111 (
            .O(N__19916),
            .I(N__19913));
    LocalMux I__2110 (
            .O(N__19913),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO ));
    CascadeMux I__2109 (
            .O(N__19910),
            .I(N__19907));
    InMux I__2108 (
            .O(N__19907),
            .I(N__19904));
    LocalMux I__2107 (
            .O(N__19904),
            .I(N__19901));
    Odrv12 I__2106 (
            .O(N__19901),
            .I(\pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9 ));
    InMux I__2105 (
            .O(N__19898),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_8 ));
    CascadeMux I__2104 (
            .O(N__19895),
            .I(N__19892));
    InMux I__2103 (
            .O(N__19892),
            .I(N__19889));
    LocalMux I__2102 (
            .O(N__19889),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9 ));
    InMux I__2101 (
            .O(N__19886),
            .I(N__19883));
    LocalMux I__2100 (
            .O(N__19883),
            .I(N__19879));
    InMux I__2099 (
            .O(N__19882),
            .I(N__19876));
    Span4Mux_s3_h I__2098 (
            .O(N__19879),
            .I(N__19873));
    LocalMux I__2097 (
            .O(N__19876),
            .I(N__19870));
    Odrv4 I__2096 (
            .O(N__19873),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    Odrv12 I__2095 (
            .O(N__19870),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    InMux I__2094 (
            .O(N__19865),
            .I(N__19862));
    LocalMux I__2093 (
            .O(N__19862),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4 ));
    CascadeMux I__2092 (
            .O(N__19859),
            .I(un2_counter_7_cascade_));
    InMux I__2091 (
            .O(N__19856),
            .I(N__19853));
    LocalMux I__2090 (
            .O(N__19853),
            .I(N__19850));
    Span4Mux_h I__2089 (
            .O(N__19850),
            .I(N__19847));
    Odrv4 I__2088 (
            .O(N__19847),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_0 ));
    CascadeMux I__2087 (
            .O(N__19844),
            .I(N__19841));
    InMux I__2086 (
            .O(N__19841),
            .I(N__19838));
    LocalMux I__2085 (
            .O(N__19838),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_1 ));
    InMux I__2084 (
            .O(N__19835),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_0 ));
    InMux I__2083 (
            .O(N__19832),
            .I(N__19829));
    LocalMux I__2082 (
            .O(N__19829),
            .I(N__19826));
    Span4Mux_v I__2081 (
            .O(N__19826),
            .I(N__19823));
    Odrv4 I__2080 (
            .O(N__19823),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_2 ));
    InMux I__2079 (
            .O(N__19820),
            .I(N__19817));
    LocalMux I__2078 (
            .O(N__19817),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2 ));
    InMux I__2077 (
            .O(N__19814),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_1 ));
    InMux I__2076 (
            .O(N__19811),
            .I(N__19808));
    LocalMux I__2075 (
            .O(N__19808),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_3 ));
    InMux I__2074 (
            .O(N__19805),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_2 ));
    InMux I__2073 (
            .O(N__19802),
            .I(N__19799));
    LocalMux I__2072 (
            .O(N__19799),
            .I(N__19796));
    Span4Mux_v I__2071 (
            .O(N__19796),
            .I(N__19792));
    InMux I__2070 (
            .O(N__19795),
            .I(N__19789));
    Odrv4 I__2069 (
            .O(N__19792),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ));
    LocalMux I__2068 (
            .O(N__19789),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ));
    InMux I__2067 (
            .O(N__19784),
            .I(N__19781));
    LocalMux I__2066 (
            .O(N__19781),
            .I(N__19776));
    CascadeMux I__2065 (
            .O(N__19780),
            .I(N__19773));
    InMux I__2064 (
            .O(N__19779),
            .I(N__19770));
    Span4Mux_v I__2063 (
            .O(N__19776),
            .I(N__19767));
    InMux I__2062 (
            .O(N__19773),
            .I(N__19764));
    LocalMux I__2061 (
            .O(N__19770),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ));
    Odrv4 I__2060 (
            .O(N__19767),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ));
    LocalMux I__2059 (
            .O(N__19764),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ));
    CascadeMux I__2058 (
            .O(N__19757),
            .I(N__19754));
    InMux I__2057 (
            .O(N__19754),
            .I(N__19751));
    LocalMux I__2056 (
            .O(N__19751),
            .I(N__19748));
    Span4Mux_v I__2055 (
            .O(N__19748),
            .I(N__19745));
    Odrv4 I__2054 (
            .O(N__19745),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO ));
    CascadeMux I__2053 (
            .O(N__19742),
            .I(\current_shift_inst.PI_CTRL.N_98_cascade_ ));
    InMux I__2052 (
            .O(N__19739),
            .I(N__19727));
    InMux I__2051 (
            .O(N__19738),
            .I(N__19727));
    InMux I__2050 (
            .O(N__19737),
            .I(N__19727));
    InMux I__2049 (
            .O(N__19736),
            .I(N__19727));
    LocalMux I__2048 (
            .O(N__19727),
            .I(N__19723));
    InMux I__2047 (
            .O(N__19726),
            .I(N__19720));
    Odrv4 I__2046 (
            .O(N__19723),
            .I(\current_shift_inst.PI_CTRL.N_96 ));
    LocalMux I__2045 (
            .O(N__19720),
            .I(\current_shift_inst.PI_CTRL.N_96 ));
    CascadeMux I__2044 (
            .O(N__19715),
            .I(N__19709));
    CascadeMux I__2043 (
            .O(N__19714),
            .I(N__19705));
    InMux I__2042 (
            .O(N__19713),
            .I(N__19700));
    InMux I__2041 (
            .O(N__19712),
            .I(N__19697));
    InMux I__2040 (
            .O(N__19709),
            .I(N__19686));
    InMux I__2039 (
            .O(N__19708),
            .I(N__19686));
    InMux I__2038 (
            .O(N__19705),
            .I(N__19686));
    InMux I__2037 (
            .O(N__19704),
            .I(N__19686));
    InMux I__2036 (
            .O(N__19703),
            .I(N__19686));
    LocalMux I__2035 (
            .O(N__19700),
            .I(N__19682));
    LocalMux I__2034 (
            .O(N__19697),
            .I(N__19676));
    LocalMux I__2033 (
            .O(N__19686),
            .I(N__19676));
    InMux I__2032 (
            .O(N__19685),
            .I(N__19673));
    Span4Mux_v I__2031 (
            .O(N__19682),
            .I(N__19670));
    InMux I__2030 (
            .O(N__19681),
            .I(N__19667));
    Span4Mux_v I__2029 (
            .O(N__19676),
            .I(N__19662));
    LocalMux I__2028 (
            .O(N__19673),
            .I(N__19662));
    Span4Mux_v I__2027 (
            .O(N__19670),
            .I(N__19659));
    LocalMux I__2026 (
            .O(N__19667),
            .I(N__19654));
    Sp12to4 I__2025 (
            .O(N__19662),
            .I(N__19654));
    Odrv4 I__2024 (
            .O(N__19659),
            .I(\current_shift_inst.PI_CTRL.N_178 ));
    Odrv12 I__2023 (
            .O(N__19654),
            .I(\current_shift_inst.PI_CTRL.N_178 ));
    InMux I__2022 (
            .O(N__19649),
            .I(N__19646));
    LocalMux I__2021 (
            .O(N__19646),
            .I(N__19643));
    Odrv4 I__2020 (
            .O(N__19643),
            .I(\current_shift_inst.PI_CTRL.N_91 ));
    CascadeMux I__2019 (
            .O(N__19640),
            .I(N__19637));
    InMux I__2018 (
            .O(N__19637),
            .I(N__19634));
    LocalMux I__2017 (
            .O(N__19634),
            .I(N__19631));
    Odrv4 I__2016 (
            .O(N__19631),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO ));
    CascadeMux I__2015 (
            .O(N__19628),
            .I(N__19624));
    InMux I__2014 (
            .O(N__19627),
            .I(N__19621));
    InMux I__2013 (
            .O(N__19624),
            .I(N__19618));
    LocalMux I__2012 (
            .O(N__19621),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ));
    LocalMux I__2011 (
            .O(N__19618),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ));
    InMux I__2010 (
            .O(N__19613),
            .I(N__19610));
    LocalMux I__2009 (
            .O(N__19610),
            .I(N__19606));
    InMux I__2008 (
            .O(N__19609),
            .I(N__19603));
    Odrv4 I__2007 (
            .O(N__19606),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ));
    LocalMux I__2006 (
            .O(N__19603),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ));
    CascadeMux I__2005 (
            .O(N__19598),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_18_cascade_ ));
    InMux I__2004 (
            .O(N__19595),
            .I(N__19592));
    LocalMux I__2003 (
            .O(N__19592),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO ));
    InMux I__2002 (
            .O(N__19589),
            .I(N__19585));
    InMux I__2001 (
            .O(N__19588),
            .I(N__19582));
    LocalMux I__2000 (
            .O(N__19585),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ));
    LocalMux I__1999 (
            .O(N__19582),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ));
    CascadeMux I__1998 (
            .O(N__19577),
            .I(N__19574));
    InMux I__1997 (
            .O(N__19574),
            .I(N__19571));
    LocalMux I__1996 (
            .O(N__19571),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO ));
    InMux I__1995 (
            .O(N__19568),
            .I(N__19563));
    InMux I__1994 (
            .O(N__19567),
            .I(N__19558));
    InMux I__1993 (
            .O(N__19566),
            .I(N__19558));
    LocalMux I__1992 (
            .O(N__19563),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ));
    LocalMux I__1991 (
            .O(N__19558),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ));
    InMux I__1990 (
            .O(N__19553),
            .I(N__19549));
    InMux I__1989 (
            .O(N__19552),
            .I(N__19546));
    LocalMux I__1988 (
            .O(N__19549),
            .I(N__19543));
    LocalMux I__1987 (
            .O(N__19546),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ));
    Odrv4 I__1986 (
            .O(N__19543),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ));
    InMux I__1985 (
            .O(N__19538),
            .I(N__19533));
    InMux I__1984 (
            .O(N__19537),
            .I(N__19530));
    InMux I__1983 (
            .O(N__19536),
            .I(N__19527));
    LocalMux I__1982 (
            .O(N__19533),
            .I(N__19522));
    LocalMux I__1981 (
            .O(N__19530),
            .I(N__19522));
    LocalMux I__1980 (
            .O(N__19527),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ));
    Odrv12 I__1979 (
            .O(N__19522),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ));
    InMux I__1978 (
            .O(N__19517),
            .I(N__19514));
    LocalMux I__1977 (
            .O(N__19514),
            .I(N__19511));
    Span4Mux_h I__1976 (
            .O(N__19511),
            .I(N__19507));
    InMux I__1975 (
            .O(N__19510),
            .I(N__19504));
    Span4Mux_v I__1974 (
            .O(N__19507),
            .I(N__19501));
    LocalMux I__1973 (
            .O(N__19504),
            .I(N__19498));
    Odrv4 I__1972 (
            .O(N__19501),
            .I(\pwm_generator_inst.O_10 ));
    Odrv4 I__1971 (
            .O(N__19498),
            .I(\pwm_generator_inst.O_10 ));
    InMux I__1970 (
            .O(N__19493),
            .I(N__19490));
    LocalMux I__1969 (
            .O(N__19490),
            .I(N__19486));
    InMux I__1968 (
            .O(N__19489),
            .I(N__19482));
    Span4Mux_v I__1967 (
            .O(N__19486),
            .I(N__19479));
    InMux I__1966 (
            .O(N__19485),
            .I(N__19476));
    LocalMux I__1965 (
            .O(N__19482),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ));
    Odrv4 I__1964 (
            .O(N__19479),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ));
    LocalMux I__1963 (
            .O(N__19476),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ));
    CascadeMux I__1962 (
            .O(N__19469),
            .I(N__19466));
    InMux I__1961 (
            .O(N__19466),
            .I(N__19463));
    LocalMux I__1960 (
            .O(N__19463),
            .I(N__19460));
    Span4Mux_v I__1959 (
            .O(N__19460),
            .I(N__19457));
    Odrv4 I__1958 (
            .O(N__19457),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO ));
    InMux I__1957 (
            .O(N__19454),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_16 ));
    InMux I__1956 (
            .O(N__19451),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_17 ));
    InMux I__1955 (
            .O(N__19448),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_18 ));
    InMux I__1954 (
            .O(N__19445),
            .I(N__19440));
    InMux I__1953 (
            .O(N__19444),
            .I(N__19437));
    InMux I__1952 (
            .O(N__19443),
            .I(N__19434));
    LocalMux I__1951 (
            .O(N__19440),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ));
    LocalMux I__1950 (
            .O(N__19437),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ));
    LocalMux I__1949 (
            .O(N__19434),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ));
    InMux I__1948 (
            .O(N__19427),
            .I(N__19423));
    InMux I__1947 (
            .O(N__19426),
            .I(N__19420));
    LocalMux I__1946 (
            .O(N__19423),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ));
    LocalMux I__1945 (
            .O(N__19420),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ));
    CascadeMux I__1944 (
            .O(N__19415),
            .I(N__19412));
    InMux I__1943 (
            .O(N__19412),
            .I(N__19409));
    LocalMux I__1942 (
            .O(N__19409),
            .I(N__19406));
    Odrv4 I__1941 (
            .O(N__19406),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO ));
    InMux I__1940 (
            .O(N__19403),
            .I(N__19400));
    LocalMux I__1939 (
            .O(N__19400),
            .I(N__19396));
    InMux I__1938 (
            .O(N__19399),
            .I(N__19393));
    Odrv4 I__1937 (
            .O(N__19396),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ));
    LocalMux I__1936 (
            .O(N__19393),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ));
    InMux I__1935 (
            .O(N__19388),
            .I(N__19384));
    InMux I__1934 (
            .O(N__19387),
            .I(N__19381));
    LocalMux I__1933 (
            .O(N__19384),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ));
    LocalMux I__1932 (
            .O(N__19381),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ));
    CascadeMux I__1931 (
            .O(N__19376),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_ ));
    InMux I__1930 (
            .O(N__19373),
            .I(N__19370));
    LocalMux I__1929 (
            .O(N__19370),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO ));
    InMux I__1928 (
            .O(N__19367),
            .I(N__19364));
    LocalMux I__1927 (
            .O(N__19364),
            .I(N__19361));
    Span4Mux_h I__1926 (
            .O(N__19361),
            .I(N__19358));
    Odrv4 I__1925 (
            .O(N__19358),
            .I(\pwm_generator_inst.O_8 ));
    InMux I__1924 (
            .O(N__19355),
            .I(N__19352));
    LocalMux I__1923 (
            .O(N__19352),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_8 ));
    InMux I__1922 (
            .O(N__19349),
            .I(N__19346));
    LocalMux I__1921 (
            .O(N__19346),
            .I(N__19343));
    Span4Mux_h I__1920 (
            .O(N__19343),
            .I(N__19340));
    Odrv4 I__1919 (
            .O(N__19340),
            .I(\pwm_generator_inst.O_9 ));
    InMux I__1918 (
            .O(N__19337),
            .I(N__19334));
    LocalMux I__1917 (
            .O(N__19334),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_9 ));
    InMux I__1916 (
            .O(N__19331),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_9 ));
    InMux I__1915 (
            .O(N__19328),
            .I(N__19325));
    LocalMux I__1914 (
            .O(N__19325),
            .I(N__19321));
    InMux I__1913 (
            .O(N__19324),
            .I(N__19318));
    Span4Mux_v I__1912 (
            .O(N__19321),
            .I(N__19315));
    LocalMux I__1911 (
            .O(N__19318),
            .I(N__19312));
    Odrv4 I__1910 (
            .O(N__19315),
            .I(\pwm_generator_inst.un3_threshold_acc ));
    Odrv4 I__1909 (
            .O(N__19312),
            .I(\pwm_generator_inst.un3_threshold_acc ));
    InMux I__1908 (
            .O(N__19307),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_10 ));
    InMux I__1907 (
            .O(N__19304),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_11 ));
    InMux I__1906 (
            .O(N__19301),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_12 ));
    InMux I__1905 (
            .O(N__19298),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_13 ));
    InMux I__1904 (
            .O(N__19295),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_14 ));
    InMux I__1903 (
            .O(N__19292),
            .I(bfn_2_9_0_));
    InMux I__1902 (
            .O(N__19289),
            .I(N__19286));
    LocalMux I__1901 (
            .O(N__19286),
            .I(N__19283));
    Span4Mux_h I__1900 (
            .O(N__19283),
            .I(N__19280));
    Odrv4 I__1899 (
            .O(N__19280),
            .I(\pwm_generator_inst.O_0 ));
    InMux I__1898 (
            .O(N__19277),
            .I(N__19274));
    LocalMux I__1897 (
            .O(N__19274),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_0 ));
    InMux I__1896 (
            .O(N__19271),
            .I(N__19268));
    LocalMux I__1895 (
            .O(N__19268),
            .I(N__19265));
    Span4Mux_h I__1894 (
            .O(N__19265),
            .I(N__19262));
    Odrv4 I__1893 (
            .O(N__19262),
            .I(\pwm_generator_inst.O_1 ));
    InMux I__1892 (
            .O(N__19259),
            .I(N__19256));
    LocalMux I__1891 (
            .O(N__19256),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_1 ));
    InMux I__1890 (
            .O(N__19253),
            .I(N__19250));
    LocalMux I__1889 (
            .O(N__19250),
            .I(N__19247));
    Span4Mux_v I__1888 (
            .O(N__19247),
            .I(N__19244));
    Odrv4 I__1887 (
            .O(N__19244),
            .I(\pwm_generator_inst.O_2 ));
    InMux I__1886 (
            .O(N__19241),
            .I(N__19238));
    LocalMux I__1885 (
            .O(N__19238),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_2 ));
    InMux I__1884 (
            .O(N__19235),
            .I(N__19232));
    LocalMux I__1883 (
            .O(N__19232),
            .I(N__19229));
    Span4Mux_v I__1882 (
            .O(N__19229),
            .I(N__19226));
    Odrv4 I__1881 (
            .O(N__19226),
            .I(\pwm_generator_inst.O_3 ));
    InMux I__1880 (
            .O(N__19223),
            .I(N__19220));
    LocalMux I__1879 (
            .O(N__19220),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_3 ));
    InMux I__1878 (
            .O(N__19217),
            .I(N__19214));
    LocalMux I__1877 (
            .O(N__19214),
            .I(N__19211));
    Span4Mux_h I__1876 (
            .O(N__19211),
            .I(N__19208));
    Odrv4 I__1875 (
            .O(N__19208),
            .I(\pwm_generator_inst.O_4 ));
    InMux I__1874 (
            .O(N__19205),
            .I(N__19202));
    LocalMux I__1873 (
            .O(N__19202),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_4 ));
    InMux I__1872 (
            .O(N__19199),
            .I(N__19196));
    LocalMux I__1871 (
            .O(N__19196),
            .I(N__19193));
    Span4Mux_h I__1870 (
            .O(N__19193),
            .I(N__19190));
    Odrv4 I__1869 (
            .O(N__19190),
            .I(\pwm_generator_inst.O_5 ));
    InMux I__1868 (
            .O(N__19187),
            .I(N__19184));
    LocalMux I__1867 (
            .O(N__19184),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_5 ));
    InMux I__1866 (
            .O(N__19181),
            .I(N__19178));
    LocalMux I__1865 (
            .O(N__19178),
            .I(N__19175));
    Span4Mux_h I__1864 (
            .O(N__19175),
            .I(N__19172));
    Odrv4 I__1863 (
            .O(N__19172),
            .I(\pwm_generator_inst.O_6 ));
    InMux I__1862 (
            .O(N__19169),
            .I(N__19166));
    LocalMux I__1861 (
            .O(N__19166),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_6 ));
    InMux I__1860 (
            .O(N__19163),
            .I(N__19160));
    LocalMux I__1859 (
            .O(N__19160),
            .I(N__19157));
    Span4Mux_h I__1858 (
            .O(N__19157),
            .I(N__19154));
    Odrv4 I__1857 (
            .O(N__19154),
            .I(\pwm_generator_inst.O_7 ));
    InMux I__1856 (
            .O(N__19151),
            .I(N__19148));
    LocalMux I__1855 (
            .O(N__19148),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_7 ));
    InMux I__1854 (
            .O(N__19145),
            .I(N__19142));
    LocalMux I__1853 (
            .O(N__19142),
            .I(un7_start_stop));
    InMux I__1852 (
            .O(N__19139),
            .I(N__19134));
    InMux I__1851 (
            .O(N__19138),
            .I(N__19129));
    InMux I__1850 (
            .O(N__19137),
            .I(N__19129));
    LocalMux I__1849 (
            .O(N__19134),
            .I(N__19126));
    LocalMux I__1848 (
            .O(N__19129),
            .I(pwm_duty_input_5));
    Odrv4 I__1847 (
            .O(N__19126),
            .I(pwm_duty_input_5));
    CascadeMux I__1846 (
            .O(N__19121),
            .I(N__19117));
    InMux I__1845 (
            .O(N__19120),
            .I(N__19113));
    InMux I__1844 (
            .O(N__19117),
            .I(N__19108));
    InMux I__1843 (
            .O(N__19116),
            .I(N__19108));
    LocalMux I__1842 (
            .O(N__19113),
            .I(N__19105));
    LocalMux I__1841 (
            .O(N__19108),
            .I(pwm_duty_input_9));
    Odrv4 I__1840 (
            .O(N__19105),
            .I(pwm_duty_input_9));
    InMux I__1839 (
            .O(N__19100),
            .I(N__19096));
    CascadeMux I__1838 (
            .O(N__19099),
            .I(N__19092));
    LocalMux I__1837 (
            .O(N__19096),
            .I(N__19089));
    InMux I__1836 (
            .O(N__19095),
            .I(N__19086));
    InMux I__1835 (
            .O(N__19092),
            .I(N__19083));
    Span4Mux_v I__1834 (
            .O(N__19089),
            .I(N__19080));
    LocalMux I__1833 (
            .O(N__19086),
            .I(pwm_duty_input_8));
    LocalMux I__1832 (
            .O(N__19083),
            .I(pwm_duty_input_8));
    Odrv4 I__1831 (
            .O(N__19080),
            .I(pwm_duty_input_8));
    CascadeMux I__1830 (
            .O(N__19073),
            .I(N__19070));
    InMux I__1829 (
            .O(N__19070),
            .I(N__19067));
    LocalMux I__1828 (
            .O(N__19067),
            .I(\current_shift_inst.PI_CTRL.m7_2 ));
    InMux I__1827 (
            .O(N__19064),
            .I(N__19059));
    InMux I__1826 (
            .O(N__19063),
            .I(N__19056));
    InMux I__1825 (
            .O(N__19062),
            .I(N__19053));
    LocalMux I__1824 (
            .O(N__19059),
            .I(N__19050));
    LocalMux I__1823 (
            .O(N__19056),
            .I(pwm_duty_input_7));
    LocalMux I__1822 (
            .O(N__19053),
            .I(pwm_duty_input_7));
    Odrv4 I__1821 (
            .O(N__19050),
            .I(pwm_duty_input_7));
    InMux I__1820 (
            .O(N__19043),
            .I(N__19040));
    LocalMux I__1819 (
            .O(N__19040),
            .I(N__19037));
    Odrv4 I__1818 (
            .O(N__19037),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ));
    CascadeMux I__1817 (
            .O(N__19034),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3_cascade_ ));
    CascadeMux I__1816 (
            .O(N__19031),
            .I(N__19027));
    InMux I__1815 (
            .O(N__19030),
            .I(N__19019));
    InMux I__1814 (
            .O(N__19027),
            .I(N__19019));
    InMux I__1813 (
            .O(N__19026),
            .I(N__19019));
    LocalMux I__1812 (
            .O(N__19019),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_3 ));
    InMux I__1811 (
            .O(N__19016),
            .I(N__19012));
    InMux I__1810 (
            .O(N__19015),
            .I(N__19009));
    LocalMux I__1809 (
            .O(N__19012),
            .I(pwm_duty_input_1));
    LocalMux I__1808 (
            .O(N__19009),
            .I(pwm_duty_input_1));
    InMux I__1807 (
            .O(N__19004),
            .I(N__18999));
    InMux I__1806 (
            .O(N__19003),
            .I(N__18996));
    InMux I__1805 (
            .O(N__19002),
            .I(N__18993));
    LocalMux I__1804 (
            .O(N__18999),
            .I(pwm_duty_input_3));
    LocalMux I__1803 (
            .O(N__18996),
            .I(pwm_duty_input_3));
    LocalMux I__1802 (
            .O(N__18993),
            .I(pwm_duty_input_3));
    CascadeMux I__1801 (
            .O(N__18986),
            .I(N__18983));
    InMux I__1800 (
            .O(N__18983),
            .I(N__18979));
    InMux I__1799 (
            .O(N__18982),
            .I(N__18976));
    LocalMux I__1798 (
            .O(N__18979),
            .I(pwm_duty_input_0));
    LocalMux I__1797 (
            .O(N__18976),
            .I(pwm_duty_input_0));
    InMux I__1796 (
            .O(N__18971),
            .I(N__18967));
    InMux I__1795 (
            .O(N__18970),
            .I(N__18964));
    LocalMux I__1794 (
            .O(N__18967),
            .I(pwm_duty_input_2));
    LocalMux I__1793 (
            .O(N__18964),
            .I(pwm_duty_input_2));
    InMux I__1792 (
            .O(N__18959),
            .I(N__18956));
    LocalMux I__1791 (
            .O(N__18956),
            .I(\current_shift_inst.PI_CTRL.m14_2 ));
    InMux I__1790 (
            .O(N__18953),
            .I(N__18932));
    InMux I__1789 (
            .O(N__18952),
            .I(N__18932));
    InMux I__1788 (
            .O(N__18951),
            .I(N__18915));
    InMux I__1787 (
            .O(N__18950),
            .I(N__18915));
    InMux I__1786 (
            .O(N__18949),
            .I(N__18915));
    InMux I__1785 (
            .O(N__18948),
            .I(N__18915));
    InMux I__1784 (
            .O(N__18947),
            .I(N__18915));
    InMux I__1783 (
            .O(N__18946),
            .I(N__18915));
    InMux I__1782 (
            .O(N__18945),
            .I(N__18915));
    InMux I__1781 (
            .O(N__18944),
            .I(N__18915));
    InMux I__1780 (
            .O(N__18943),
            .I(N__18900));
    InMux I__1779 (
            .O(N__18942),
            .I(N__18900));
    InMux I__1778 (
            .O(N__18941),
            .I(N__18900));
    InMux I__1777 (
            .O(N__18940),
            .I(N__18900));
    InMux I__1776 (
            .O(N__18939),
            .I(N__18900));
    InMux I__1775 (
            .O(N__18938),
            .I(N__18900));
    InMux I__1774 (
            .O(N__18937),
            .I(N__18900));
    LocalMux I__1773 (
            .O(N__18932),
            .I(N__18897));
    LocalMux I__1772 (
            .O(N__18915),
            .I(N__18892));
    LocalMux I__1771 (
            .O(N__18900),
            .I(N__18892));
    Span4Mux_h I__1770 (
            .O(N__18897),
            .I(N__18880));
    Span4Mux_v I__1769 (
            .O(N__18892),
            .I(N__18880));
    InMux I__1768 (
            .O(N__18891),
            .I(N__18875));
    InMux I__1767 (
            .O(N__18890),
            .I(N__18875));
    InMux I__1766 (
            .O(N__18889),
            .I(N__18868));
    InMux I__1765 (
            .O(N__18888),
            .I(N__18868));
    InMux I__1764 (
            .O(N__18887),
            .I(N__18868));
    InMux I__1763 (
            .O(N__18886),
            .I(N__18863));
    InMux I__1762 (
            .O(N__18885),
            .I(N__18863));
    Span4Mux_v I__1761 (
            .O(N__18880),
            .I(N__18856));
    LocalMux I__1760 (
            .O(N__18875),
            .I(N__18856));
    LocalMux I__1759 (
            .O(N__18868),
            .I(N__18856));
    LocalMux I__1758 (
            .O(N__18863),
            .I(pwm_duty_input_10));
    Odrv4 I__1757 (
            .O(N__18856),
            .I(pwm_duty_input_10));
    CascadeMux I__1756 (
            .O(N__18851),
            .I(\current_shift_inst.PI_CTRL.N_19_cascade_ ));
    InMux I__1755 (
            .O(N__18848),
            .I(N__18843));
    InMux I__1754 (
            .O(N__18847),
            .I(N__18840));
    InMux I__1753 (
            .O(N__18846),
            .I(N__18837));
    LocalMux I__1752 (
            .O(N__18843),
            .I(pwm_duty_input_4));
    LocalMux I__1751 (
            .O(N__18840),
            .I(pwm_duty_input_4));
    LocalMux I__1750 (
            .O(N__18837),
            .I(pwm_duty_input_4));
    CascadeMux I__1749 (
            .O(N__18830),
            .I(N__18827));
    InMux I__1748 (
            .O(N__18827),
            .I(N__18824));
    LocalMux I__1747 (
            .O(N__18824),
            .I(N__18821));
    Span4Mux_v I__1746 (
            .O(N__18821),
            .I(N__18818));
    Odrv4 I__1745 (
            .O(N__18818),
            .I(\pwm_generator_inst.un2_threshold_acc_2_10 ));
    InMux I__1744 (
            .O(N__18815),
            .I(N__18812));
    LocalMux I__1743 (
            .O(N__18812),
            .I(N__18809));
    Odrv4 I__1742 (
            .O(N__18809),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0 ));
    InMux I__1741 (
            .O(N__18806),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ));
    InMux I__1740 (
            .O(N__18803),
            .I(N__18800));
    LocalMux I__1739 (
            .O(N__18800),
            .I(N__18797));
    Span4Mux_v I__1738 (
            .O(N__18797),
            .I(N__18794));
    Odrv4 I__1737 (
            .O(N__18794),
            .I(\pwm_generator_inst.un2_threshold_acc_2_11 ));
    CascadeMux I__1736 (
            .O(N__18791),
            .I(N__18788));
    InMux I__1735 (
            .O(N__18788),
            .I(N__18785));
    LocalMux I__1734 (
            .O(N__18785),
            .I(N__18782));
    Odrv4 I__1733 (
            .O(N__18782),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0 ));
    InMux I__1732 (
            .O(N__18779),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ));
    CascadeMux I__1731 (
            .O(N__18776),
            .I(N__18773));
    InMux I__1730 (
            .O(N__18773),
            .I(N__18770));
    LocalMux I__1729 (
            .O(N__18770),
            .I(N__18767));
    Span4Mux_h I__1728 (
            .O(N__18767),
            .I(N__18764));
    Odrv4 I__1727 (
            .O(N__18764),
            .I(\pwm_generator_inst.un2_threshold_acc_2_12 ));
    InMux I__1726 (
            .O(N__18761),
            .I(N__18758));
    LocalMux I__1725 (
            .O(N__18758),
            .I(N__18755));
    Odrv4 I__1724 (
            .O(N__18755),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0 ));
    InMux I__1723 (
            .O(N__18752),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ));
    InMux I__1722 (
            .O(N__18749),
            .I(N__18746));
    LocalMux I__1721 (
            .O(N__18746),
            .I(N__18743));
    Span4Mux_v I__1720 (
            .O(N__18743),
            .I(N__18740));
    Odrv4 I__1719 (
            .O(N__18740),
            .I(\pwm_generator_inst.un2_threshold_acc_2_13 ));
    InMux I__1718 (
            .O(N__18737),
            .I(N__18734));
    LocalMux I__1717 (
            .O(N__18734),
            .I(N__18731));
    Odrv4 I__1716 (
            .O(N__18731),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0 ));
    InMux I__1715 (
            .O(N__18728),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ));
    CascadeMux I__1714 (
            .O(N__18725),
            .I(N__18722));
    InMux I__1713 (
            .O(N__18722),
            .I(N__18719));
    LocalMux I__1712 (
            .O(N__18719),
            .I(N__18716));
    Span4Mux_h I__1711 (
            .O(N__18716),
            .I(N__18713));
    Odrv4 I__1710 (
            .O(N__18713),
            .I(\pwm_generator_inst.un2_threshold_acc_2_14 ));
    InMux I__1709 (
            .O(N__18710),
            .I(N__18707));
    LocalMux I__1708 (
            .O(N__18707),
            .I(N__18704));
    Odrv4 I__1707 (
            .O(N__18704),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0 ));
    InMux I__1706 (
            .O(N__18701),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ));
    InMux I__1705 (
            .O(N__18698),
            .I(N__18695));
    LocalMux I__1704 (
            .O(N__18695),
            .I(N__18692));
    Odrv4 I__1703 (
            .O(N__18692),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0 ));
    CascadeMux I__1702 (
            .O(N__18689),
            .I(N__18682));
    CascadeMux I__1701 (
            .O(N__18688),
            .I(N__18678));
    CascadeMux I__1700 (
            .O(N__18687),
            .I(N__18674));
    InMux I__1699 (
            .O(N__18686),
            .I(N__18668));
    InMux I__1698 (
            .O(N__18685),
            .I(N__18668));
    InMux I__1697 (
            .O(N__18682),
            .I(N__18655));
    InMux I__1696 (
            .O(N__18681),
            .I(N__18655));
    InMux I__1695 (
            .O(N__18678),
            .I(N__18655));
    InMux I__1694 (
            .O(N__18677),
            .I(N__18655));
    InMux I__1693 (
            .O(N__18674),
            .I(N__18655));
    InMux I__1692 (
            .O(N__18673),
            .I(N__18655));
    LocalMux I__1691 (
            .O(N__18668),
            .I(N__18650));
    LocalMux I__1690 (
            .O(N__18655),
            .I(N__18650));
    Span4Mux_v I__1689 (
            .O(N__18650),
            .I(N__18647));
    Odrv4 I__1688 (
            .O(N__18647),
            .I(\pwm_generator_inst.un2_threshold_acc_1_25 ));
    InMux I__1687 (
            .O(N__18644),
            .I(N__18641));
    LocalMux I__1686 (
            .O(N__18641),
            .I(N__18638));
    Odrv4 I__1685 (
            .O(N__18638),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0 ));
    InMux I__1684 (
            .O(N__18635),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ));
    InMux I__1683 (
            .O(N__18632),
            .I(N__18629));
    LocalMux I__1682 (
            .O(N__18629),
            .I(N__18626));
    Odrv4 I__1681 (
            .O(N__18626),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16 ));
    InMux I__1680 (
            .O(N__18623),
            .I(N__18620));
    LocalMux I__1679 (
            .O(N__18620),
            .I(N__18617));
    Odrv4 I__1678 (
            .O(N__18617),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO ));
    InMux I__1677 (
            .O(N__18614),
            .I(bfn_1_14_0_));
    InMux I__1676 (
            .O(N__18611),
            .I(N__18608));
    LocalMux I__1675 (
            .O(N__18608),
            .I(N_110_i_i));
    InMux I__1674 (
            .O(N__18605),
            .I(N__18602));
    LocalMux I__1673 (
            .O(N__18602),
            .I(N__18599));
    Span4Mux_v I__1672 (
            .O(N__18599),
            .I(N__18596));
    Odrv4 I__1671 (
            .O(N__18596),
            .I(\pwm_generator_inst.un2_threshold_acc_1_18 ));
    CascadeMux I__1670 (
            .O(N__18593),
            .I(N__18590));
    InMux I__1669 (
            .O(N__18590),
            .I(N__18587));
    LocalMux I__1668 (
            .O(N__18587),
            .I(N__18584));
    Span4Mux_v I__1667 (
            .O(N__18584),
            .I(N__18581));
    Odrv4 I__1666 (
            .O(N__18581),
            .I(\pwm_generator_inst.un2_threshold_acc_2_3 ));
    CascadeMux I__1665 (
            .O(N__18578),
            .I(N__18575));
    InMux I__1664 (
            .O(N__18575),
            .I(N__18572));
    LocalMux I__1663 (
            .O(N__18572),
            .I(N__18569));
    Odrv4 I__1662 (
            .O(N__18569),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0 ));
    InMux I__1661 (
            .O(N__18566),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ));
    InMux I__1660 (
            .O(N__18563),
            .I(N__18560));
    LocalMux I__1659 (
            .O(N__18560),
            .I(N__18557));
    Span4Mux_v I__1658 (
            .O(N__18557),
            .I(N__18554));
    Odrv4 I__1657 (
            .O(N__18554),
            .I(\pwm_generator_inst.un2_threshold_acc_1_19 ));
    CascadeMux I__1656 (
            .O(N__18551),
            .I(N__18548));
    InMux I__1655 (
            .O(N__18548),
            .I(N__18545));
    LocalMux I__1654 (
            .O(N__18545),
            .I(N__18542));
    Odrv4 I__1653 (
            .O(N__18542),
            .I(\pwm_generator_inst.un2_threshold_acc_2_4 ));
    InMux I__1652 (
            .O(N__18539),
            .I(N__18536));
    LocalMux I__1651 (
            .O(N__18536),
            .I(N__18533));
    Odrv4 I__1650 (
            .O(N__18533),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0 ));
    InMux I__1649 (
            .O(N__18530),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ));
    InMux I__1648 (
            .O(N__18527),
            .I(N__18524));
    LocalMux I__1647 (
            .O(N__18524),
            .I(N__18521));
    Span4Mux_v I__1646 (
            .O(N__18521),
            .I(N__18518));
    Odrv4 I__1645 (
            .O(N__18518),
            .I(\pwm_generator_inst.un2_threshold_acc_1_20 ));
    CascadeMux I__1644 (
            .O(N__18515),
            .I(N__18512));
    InMux I__1643 (
            .O(N__18512),
            .I(N__18509));
    LocalMux I__1642 (
            .O(N__18509),
            .I(N__18506));
    Span4Mux_h I__1641 (
            .O(N__18506),
            .I(N__18503));
    Odrv4 I__1640 (
            .O(N__18503),
            .I(\pwm_generator_inst.un2_threshold_acc_2_5 ));
    InMux I__1639 (
            .O(N__18500),
            .I(N__18497));
    LocalMux I__1638 (
            .O(N__18497),
            .I(N__18494));
    Odrv4 I__1637 (
            .O(N__18494),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0 ));
    InMux I__1636 (
            .O(N__18491),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ));
    InMux I__1635 (
            .O(N__18488),
            .I(N__18485));
    LocalMux I__1634 (
            .O(N__18485),
            .I(N__18482));
    Span4Mux_v I__1633 (
            .O(N__18482),
            .I(N__18479));
    Odrv4 I__1632 (
            .O(N__18479),
            .I(\pwm_generator_inst.un2_threshold_acc_1_21 ));
    CascadeMux I__1631 (
            .O(N__18476),
            .I(N__18473));
    InMux I__1630 (
            .O(N__18473),
            .I(N__18470));
    LocalMux I__1629 (
            .O(N__18470),
            .I(N__18467));
    Span4Mux_h I__1628 (
            .O(N__18467),
            .I(N__18464));
    Odrv4 I__1627 (
            .O(N__18464),
            .I(\pwm_generator_inst.un2_threshold_acc_2_6 ));
    InMux I__1626 (
            .O(N__18461),
            .I(N__18458));
    LocalMux I__1625 (
            .O(N__18458),
            .I(N__18455));
    Odrv4 I__1624 (
            .O(N__18455),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0 ));
    InMux I__1623 (
            .O(N__18452),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ));
    InMux I__1622 (
            .O(N__18449),
            .I(N__18446));
    LocalMux I__1621 (
            .O(N__18446),
            .I(N__18443));
    Span4Mux_v I__1620 (
            .O(N__18443),
            .I(N__18440));
    Odrv4 I__1619 (
            .O(N__18440),
            .I(\pwm_generator_inst.un2_threshold_acc_1_22 ));
    CascadeMux I__1618 (
            .O(N__18437),
            .I(N__18434));
    InMux I__1617 (
            .O(N__18434),
            .I(N__18431));
    LocalMux I__1616 (
            .O(N__18431),
            .I(N__18428));
    Odrv4 I__1615 (
            .O(N__18428),
            .I(\pwm_generator_inst.un2_threshold_acc_2_7 ));
    InMux I__1614 (
            .O(N__18425),
            .I(N__18422));
    LocalMux I__1613 (
            .O(N__18422),
            .I(N__18419));
    Odrv4 I__1612 (
            .O(N__18419),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0 ));
    InMux I__1611 (
            .O(N__18416),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ));
    InMux I__1610 (
            .O(N__18413),
            .I(N__18410));
    LocalMux I__1609 (
            .O(N__18410),
            .I(N__18407));
    Span4Mux_v I__1608 (
            .O(N__18407),
            .I(N__18404));
    Odrv4 I__1607 (
            .O(N__18404),
            .I(\pwm_generator_inst.un2_threshold_acc_1_23 ));
    CascadeMux I__1606 (
            .O(N__18401),
            .I(N__18398));
    InMux I__1605 (
            .O(N__18398),
            .I(N__18395));
    LocalMux I__1604 (
            .O(N__18395),
            .I(N__18392));
    Odrv4 I__1603 (
            .O(N__18392),
            .I(\pwm_generator_inst.un2_threshold_acc_2_8 ));
    CascadeMux I__1602 (
            .O(N__18389),
            .I(N__18386));
    InMux I__1601 (
            .O(N__18386),
            .I(N__18383));
    LocalMux I__1600 (
            .O(N__18383),
            .I(N__18380));
    Odrv4 I__1599 (
            .O(N__18380),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0 ));
    InMux I__1598 (
            .O(N__18377),
            .I(bfn_1_13_0_));
    InMux I__1597 (
            .O(N__18374),
            .I(N__18371));
    LocalMux I__1596 (
            .O(N__18371),
            .I(N__18368));
    Span4Mux_v I__1595 (
            .O(N__18368),
            .I(N__18365));
    Span4Mux_s1_h I__1594 (
            .O(N__18365),
            .I(N__18362));
    Odrv4 I__1593 (
            .O(N__18362),
            .I(\pwm_generator_inst.un2_threshold_acc_1_24 ));
    CascadeMux I__1592 (
            .O(N__18359),
            .I(N__18356));
    InMux I__1591 (
            .O(N__18356),
            .I(N__18353));
    LocalMux I__1590 (
            .O(N__18353),
            .I(N__18350));
    Span4Mux_h I__1589 (
            .O(N__18350),
            .I(N__18347));
    Odrv4 I__1588 (
            .O(N__18347),
            .I(\pwm_generator_inst.un2_threshold_acc_2_9 ));
    InMux I__1587 (
            .O(N__18344),
            .I(N__18341));
    LocalMux I__1586 (
            .O(N__18341),
            .I(N__18338));
    Odrv4 I__1585 (
            .O(N__18338),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0 ));
    InMux I__1584 (
            .O(N__18335),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ));
    InMux I__1583 (
            .O(N__18332),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_19 ));
    InMux I__1582 (
            .O(N__18329),
            .I(N__18326));
    LocalMux I__1581 (
            .O(N__18326),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1_16 ));
    CascadeMux I__1580 (
            .O(N__18323),
            .I(N__18320));
    InMux I__1579 (
            .O(N__18320),
            .I(N__18314));
    InMux I__1578 (
            .O(N__18319),
            .I(N__18314));
    LocalMux I__1577 (
            .O(N__18314),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1_15 ));
    InMux I__1576 (
            .O(N__18311),
            .I(N__18308));
    LocalMux I__1575 (
            .O(N__18308),
            .I(N__18305));
    Odrv4 I__1574 (
            .O(N__18305),
            .I(\pwm_generator_inst.un2_threshold_acc_2_0 ));
    CascadeMux I__1573 (
            .O(N__18302),
            .I(N__18299));
    InMux I__1572 (
            .O(N__18299),
            .I(N__18296));
    LocalMux I__1571 (
            .O(N__18296),
            .I(N__18293));
    Span4Mux_v I__1570 (
            .O(N__18293),
            .I(N__18290));
    Odrv4 I__1569 (
            .O(N__18290),
            .I(\pwm_generator_inst.un2_threshold_acc_1_15 ));
    InMux I__1568 (
            .O(N__18287),
            .I(N__18284));
    LocalMux I__1567 (
            .O(N__18284),
            .I(N__18281));
    Odrv4 I__1566 (
            .O(N__18281),
            .I(\pwm_generator_inst.un3_threshold_acc_axbZ0Z_4 ));
    InMux I__1565 (
            .O(N__18278),
            .I(N__18275));
    LocalMux I__1564 (
            .O(N__18275),
            .I(N__18272));
    Span4Mux_v I__1563 (
            .O(N__18272),
            .I(N__18269));
    Odrv4 I__1562 (
            .O(N__18269),
            .I(\pwm_generator_inst.un2_threshold_acc_1_16 ));
    CascadeMux I__1561 (
            .O(N__18266),
            .I(N__18263));
    InMux I__1560 (
            .O(N__18263),
            .I(N__18260));
    LocalMux I__1559 (
            .O(N__18260),
            .I(N__18257));
    Odrv4 I__1558 (
            .O(N__18257),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1 ));
    CascadeMux I__1557 (
            .O(N__18254),
            .I(N__18251));
    InMux I__1556 (
            .O(N__18251),
            .I(N__18248));
    LocalMux I__1555 (
            .O(N__18248),
            .I(N__18245));
    Odrv4 I__1554 (
            .O(N__18245),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0 ));
    InMux I__1553 (
            .O(N__18242),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ));
    InMux I__1552 (
            .O(N__18239),
            .I(N__18236));
    LocalMux I__1551 (
            .O(N__18236),
            .I(N__18233));
    Span4Mux_v I__1550 (
            .O(N__18233),
            .I(N__18230));
    Odrv4 I__1549 (
            .O(N__18230),
            .I(\pwm_generator_inst.un2_threshold_acc_1_17 ));
    CascadeMux I__1548 (
            .O(N__18227),
            .I(N__18224));
    InMux I__1547 (
            .O(N__18224),
            .I(N__18221));
    LocalMux I__1546 (
            .O(N__18221),
            .I(N__18218));
    Span4Mux_v I__1545 (
            .O(N__18218),
            .I(N__18215));
    Odrv4 I__1544 (
            .O(N__18215),
            .I(\pwm_generator_inst.un2_threshold_acc_2_2 ));
    InMux I__1543 (
            .O(N__18212),
            .I(N__18209));
    LocalMux I__1542 (
            .O(N__18209),
            .I(N__18206));
    Odrv4 I__1541 (
            .O(N__18206),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0 ));
    InMux I__1540 (
            .O(N__18203),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ));
    InMux I__1539 (
            .O(N__18200),
            .I(bfn_1_10_0_));
    InMux I__1538 (
            .O(N__18197),
            .I(N__18194));
    LocalMux I__1537 (
            .O(N__18194),
            .I(N__18191));
    Odrv4 I__1536 (
            .O(N__18191),
            .I(\pwm_generator_inst.O_12 ));
    InMux I__1535 (
            .O(N__18188),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_0 ));
    InMux I__1534 (
            .O(N__18185),
            .I(N__18182));
    LocalMux I__1533 (
            .O(N__18182),
            .I(N__18179));
    Odrv4 I__1532 (
            .O(N__18179),
            .I(\pwm_generator_inst.O_13 ));
    InMux I__1531 (
            .O(N__18176),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_1 ));
    InMux I__1530 (
            .O(N__18173),
            .I(N__18170));
    LocalMux I__1529 (
            .O(N__18170),
            .I(N__18167));
    Span4Mux_h I__1528 (
            .O(N__18167),
            .I(N__18164));
    Odrv4 I__1527 (
            .O(N__18164),
            .I(\pwm_generator_inst.O_14 ));
    InMux I__1526 (
            .O(N__18161),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_2 ));
    InMux I__1525 (
            .O(N__18158),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_3 ));
    InMux I__1524 (
            .O(N__18155),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_4 ));
    InMux I__1523 (
            .O(N__18152),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_5 ));
    InMux I__1522 (
            .O(N__18149),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_6 ));
    InMux I__1521 (
            .O(N__18146),
            .I(N__18137));
    InMux I__1520 (
            .O(N__18145),
            .I(N__18137));
    InMux I__1519 (
            .O(N__18144),
            .I(N__18137));
    LocalMux I__1518 (
            .O(N__18137),
            .I(N__18134));
    Odrv4 I__1517 (
            .O(N__18134),
            .I(\current_shift_inst.PI_CTRL.N_97 ));
    defparam IN_MUX_bfv_8_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_17_0_));
    defparam IN_MUX_bfv_8_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_18_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_0_cry_6 ),
            .carryinitout(bfn_8_18_0_));
    defparam IN_MUX_bfv_8_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_19_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_0_cry_14 ),
            .carryinitout(bfn_8_19_0_));
    defparam IN_MUX_bfv_8_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_20_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_0_cry_22 ),
            .carryinitout(bfn_8_20_0_));
    defparam IN_MUX_bfv_8_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_21_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_0_cry_30 ),
            .carryinitout(bfn_8_21_0_));
    defparam IN_MUX_bfv_4_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_7_0_));
    defparam IN_MUX_bfv_4_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_8_0_ (
            .carryinitin(un5_counter_cry_8),
            .carryinitout(bfn_4_8_0_));
    defparam IN_MUX_bfv_1_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_9_0_));
    defparam IN_MUX_bfv_1_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_10_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_acc_cry_7 ),
            .carryinitout(bfn_1_10_0_));
    defparam IN_MUX_bfv_1_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_11_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_acc_cry_15 ),
            .carryinitout(bfn_1_11_0_));
    defparam IN_MUX_bfv_14_22_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_22_0_));
    defparam IN_MUX_bfv_14_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_23_0_ (
            .carryinitin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_14_23_0_));
    defparam IN_MUX_bfv_14_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_24_0_ (
            .carryinitin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_14_24_0_));
    defparam IN_MUX_bfv_15_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_17_0_));
    defparam IN_MUX_bfv_15_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_18_0_ (
            .carryinitin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_15_18_0_));
    defparam IN_MUX_bfv_15_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_19_0_ (
            .carryinitin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_15_19_0_));
    defparam IN_MUX_bfv_13_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_23_0_));
    defparam IN_MUX_bfv_13_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_24_0_ (
            .carryinitin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_13_24_0_));
    defparam IN_MUX_bfv_13_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_25_0_ (
            .carryinitin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_13_25_0_));
    defparam IN_MUX_bfv_18_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_17_0_));
    defparam IN_MUX_bfv_18_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_18_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_18_18_0_));
    defparam IN_MUX_bfv_18_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_19_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_18_19_0_));
    defparam IN_MUX_bfv_8_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_11_0_));
    defparam IN_MUX_bfv_8_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_12_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_8_12_0_));
    defparam IN_MUX_bfv_8_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_13_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_8_13_0_));
    defparam IN_MUX_bfv_11_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_8_0_));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_11_9_0_));
    defparam IN_MUX_bfv_11_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_10_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_11_10_0_));
    defparam IN_MUX_bfv_10_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_18_0_));
    defparam IN_MUX_bfv_10_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_19_0_ (
            .carryinitin(\current_shift_inst.z_5_cry_8 ),
            .carryinitout(bfn_10_19_0_));
    defparam IN_MUX_bfv_10_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_20_0_ (
            .carryinitin(\current_shift_inst.z_5_cry_16 ),
            .carryinitout(bfn_10_20_0_));
    defparam IN_MUX_bfv_10_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_21_0_ (
            .carryinitin(\current_shift_inst.z_5_cry_24 ),
            .carryinitout(bfn_10_21_0_));
    defparam IN_MUX_bfv_1_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_12_0_));
    defparam IN_MUX_bfv_1_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_13_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7 ),
            .carryinitout(bfn_1_13_0_));
    defparam IN_MUX_bfv_1_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_14_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15 ),
            .carryinitout(bfn_1_14_0_));
    defparam IN_MUX_bfv_2_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_7_0_));
    defparam IN_MUX_bfv_2_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_8_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_acc_1_cry_7 ),
            .carryinitout(bfn_2_8_0_));
    defparam IN_MUX_bfv_2_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_9_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_acc_1_cry_15 ),
            .carryinitout(bfn_2_9_0_));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_8_0_));
    defparam IN_MUX_bfv_9_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_9_0_ (
            .carryinitin(\pwm_generator_inst.un14_counter_cry_7 ),
            .carryinitout(bfn_9_9_0_));
    defparam IN_MUX_bfv_3_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_9_0_));
    defparam IN_MUX_bfv_3_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_10_0_ (
            .carryinitin(\pwm_generator_inst.un19_threshold_acc_cry_7 ),
            .carryinitout(bfn_3_10_0_));
    defparam IN_MUX_bfv_10_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_9_0_));
    defparam IN_MUX_bfv_10_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_10_0_ (
            .carryinitin(\pwm_generator_inst.counter_cry_7 ),
            .carryinitout(bfn_10_10_0_));
    defparam IN_MUX_bfv_13_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_19_0_));
    defparam IN_MUX_bfv_13_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_20_0_ (
            .carryinitin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryinitout(bfn_13_20_0_));
    defparam IN_MUX_bfv_13_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_21_0_ (
            .carryinitin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryinitout(bfn_13_21_0_));
    defparam IN_MUX_bfv_16_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_19_0_));
    defparam IN_MUX_bfv_16_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_20_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryinitout(bfn_16_20_0_));
    defparam IN_MUX_bfv_16_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_21_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryinitout(bfn_16_21_0_));
    defparam IN_MUX_bfv_18_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_13_0_));
    defparam IN_MUX_bfv_18_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_14_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_18_14_0_));
    defparam IN_MUX_bfv_18_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_15_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_18_15_0_));
    defparam IN_MUX_bfv_18_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_16_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_18_16_0_));
    defparam IN_MUX_bfv_17_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_11_0_));
    defparam IN_MUX_bfv_17_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_12_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .carryinitout(bfn_17_12_0_));
    defparam IN_MUX_bfv_17_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_13_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .carryinitout(bfn_17_13_0_));
    defparam IN_MUX_bfv_17_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_14_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .carryinitout(bfn_17_14_0_));
    defparam IN_MUX_bfv_15_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_7_0_));
    defparam IN_MUX_bfv_15_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_8_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_15_8_0_));
    defparam IN_MUX_bfv_15_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_9_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_15_9_0_));
    defparam IN_MUX_bfv_15_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_10_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_15_10_0_));
    defparam IN_MUX_bfv_16_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_7_0_));
    defparam IN_MUX_bfv_16_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_8_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .carryinitout(bfn_16_8_0_));
    defparam IN_MUX_bfv_16_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_9_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .carryinitout(bfn_16_9_0_));
    defparam IN_MUX_bfv_16_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_10_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .carryinitout(bfn_16_10_0_));
    defparam IN_MUX_bfv_10_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_14_0_));
    defparam IN_MUX_bfv_10_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_15_0_ (
            .carryinitin(\current_shift_inst.z_cry_7 ),
            .carryinitout(bfn_10_15_0_));
    defparam IN_MUX_bfv_10_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_16_0_ (
            .carryinitin(\current_shift_inst.z_cry_15 ),
            .carryinitout(bfn_10_16_0_));
    defparam IN_MUX_bfv_10_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_17_0_ (
            .carryinitin(\current_shift_inst.z_cry_23 ),
            .carryinitout(bfn_10_17_0_));
    defparam IN_MUX_bfv_11_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_14_0_));
    defparam IN_MUX_bfv_11_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_15_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_cry_8 ),
            .carryinitout(bfn_11_15_0_));
    defparam IN_MUX_bfv_11_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_16_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_cry_16 ),
            .carryinitout(bfn_11_16_0_));
    defparam IN_MUX_bfv_11_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_17_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_cry_24 ),
            .carryinitout(bfn_11_17_0_));
    defparam IN_MUX_bfv_13_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_13_0_));
    defparam IN_MUX_bfv_13_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_14_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_13_14_0_));
    defparam IN_MUX_bfv_13_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_15_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_13_15_0_));
    defparam IN_MUX_bfv_13_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_16_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_13_16_0_));
    defparam IN_MUX_bfv_15_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_13_0_));
    defparam IN_MUX_bfv_15_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_14_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_7 ),
            .carryinitout(bfn_15_14_0_));
    defparam IN_MUX_bfv_15_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_15_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_15 ),
            .carryinitout(bfn_15_15_0_));
    defparam IN_MUX_bfv_15_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_16_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_23 ),
            .carryinitout(bfn_15_16_0_));
    defparam IN_MUX_bfv_9_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_21_0_));
    defparam IN_MUX_bfv_9_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_22_0_ (
            .carryinitin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_9_22_0_));
    defparam IN_MUX_bfv_9_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_23_0_ (
            .carryinitin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_9_23_0_));
    defparam IN_MUX_bfv_9_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_24_0_ (
            .carryinitin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_9_24_0_));
    defparam IN_MUX_bfv_9_25_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_25_0_));
    defparam IN_MUX_bfv_9_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_26_0_ (
            .carryinitin(\current_shift_inst.timer_phase.counter_cry_7 ),
            .carryinitout(bfn_9_26_0_));
    defparam IN_MUX_bfv_9_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_27_0_ (
            .carryinitin(\current_shift_inst.timer_phase.counter_cry_15 ),
            .carryinitout(bfn_9_27_0_));
    defparam IN_MUX_bfv_9_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_28_0_ (
            .carryinitin(\current_shift_inst.timer_phase.counter_cry_23 ),
            .carryinitout(bfn_9_28_0_));
    defparam IN_MUX_bfv_7_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_17_0_));
    defparam IN_MUX_bfv_7_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_18_0_ (
            .carryinitin(\current_shift_inst.control_input_1_cry_7 ),
            .carryinitout(bfn_7_18_0_));
    defparam IN_MUX_bfv_7_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_19_0_ (
            .carryinitin(\current_shift_inst.control_input_1_cry_15 ),
            .carryinitout(bfn_7_19_0_));
    defparam IN_MUX_bfv_7_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_20_0_ (
            .carryinitin(\current_shift_inst.control_input_1_cry_23 ),
            .carryinitout(bfn_7_20_0_));
    defparam IN_MUX_bfv_4_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_13_0_));
    defparam IN_MUX_bfv_4_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_14_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .carryinitout(bfn_4_14_0_));
    defparam IN_MUX_bfv_4_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_15_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .carryinitout(bfn_4_15_0_));
    defparam IN_MUX_bfv_4_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_16_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .carryinitout(bfn_4_16_0_));
    defparam IN_MUX_bfv_9_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_13_0_));
    defparam IN_MUX_bfv_9_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_14_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ),
            .carryinitout(bfn_9_14_0_));
    defparam IN_MUX_bfv_9_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_15_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ),
            .carryinitout(bfn_9_15_0_));
    defparam IN_MUX_bfv_9_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_16_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ),
            .carryinitout(bfn_9_16_0_));
    ICE_GB \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_0  (
            .USERSIGNALTOGLOBALBUFFER(N__32273),
            .GLOBALBUFFEROUTPUT(\delay_measurement_inst.delay_hc_timer.N_321_i_g ));
    ICE_GB \current_shift_inst.timer_s1.running_RNII51H_0  (
            .USERSIGNALTOGLOBALBUFFER(N__32414),
            .GLOBALBUFFEROUTPUT(\current_shift_inst.timer_s1.N_187_i_g ));
    ICE_GB \current_shift_inst.timer_phase.running_RNIC90O_0  (
            .USERSIGNALTOGLOBALBUFFER(N__33452),
            .GLOBALBUFFEROUTPUT(\current_shift_inst.timer_phase.N_188_i_g ));
    defparam osc.CLKHF_DIV="0b10";
    SB_HFOSC osc (
            .CLKHFPU(N__28547),
            .CLKHFEN(N__28548),
            .CLKHF(clk_12mhz));
    defparam rgb_drv.RGB2_CURRENT="0b111111";
    defparam rgb_drv.CURRENT_MODE="0b0";
    defparam rgb_drv.RGB0_CURRENT="0b111111";
    defparam rgb_drv.RGB1_CURRENT="0b111111";
    SB_RGBA_DRV rgb_drv (
            .RGBLEDEN(N__28528),
            .RGB2PWM(N__18611),
            .RGB1(rgb_g),
            .CURREN(N__28656),
            .RGB2(rgb_b),
            .RGB1PWM(N__19145),
            .RGB0PWM(N__46780),
            .RGB0(rgb_r));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_5_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_5_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_5_0 .LUT_INIT=16'b1010111000001110;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_5_LC_1_5_0  (
            .in0(N__20501),
            .in1(N__19703),
            .in2(N__21265),
            .in3(N__20001),
            .lcout(pwm_duty_input_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47351),
            .ce(N__23648),
            .sr(N__46683));
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_5_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_5_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_5_1 .LUT_INIT=16'b1011101100110000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_7_LC_1_5_1  (
            .in0(N__20003),
            .in1(N__21253),
            .in2(N__19714),
            .in3(N__21062),
            .lcout(pwm_duty_input_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47351),
            .ce(N__23648),
            .sr(N__46683));
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_5_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_5_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_5_2 .LUT_INIT=16'b1010111000001110;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_8_LC_1_5_2  (
            .in0(N__21029),
            .in1(N__19708),
            .in2(N__21267),
            .in3(N__20004),
            .lcout(pwm_duty_input_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47351),
            .ce(N__23648),
            .sr(N__46683));
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_5_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_5_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_5_3 .LUT_INIT=16'b1011101100110000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_9_LC_1_5_3  (
            .in0(N__20005),
            .in1(N__21257),
            .in2(N__19715),
            .in3(N__20987),
            .lcout(pwm_duty_input_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47351),
            .ce(N__23648),
            .sr(N__46683));
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_5_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_5_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_5_4 .LUT_INIT=16'b1010111000001110;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_6_LC_1_5_4  (
            .in0(N__20471),
            .in1(N__19704),
            .in2(N__21266),
            .in3(N__20002),
            .lcout(pwm_duty_input_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47351),
            .ce(N__23648),
            .sr(N__46683));
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_6_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_6_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_6_0 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_0_LC_1_6_0  (
            .in0(N__18144),
            .in1(N__19026),
            .in2(N__20651),
            .in3(N__19736),
            .lcout(pwm_duty_input_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47350),
            .ce(N__23672),
            .sr(N__46693));
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_6_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_6_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_6_1 .LUT_INIT=16'b1111010111110001;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_3_LC_1_6_1  (
            .in0(N__19739),
            .in1(N__19043),
            .in2(N__20594),
            .in3(N__19712),
            .lcout(pwm_duty_input_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47350),
            .ce(N__23672),
            .sr(N__46693));
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_6_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_6_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_6_2 .LUT_INIT=16'b0101000101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_4_LC_1_6_2  (
            .in0(N__19649),
            .in1(N__19886),
            .in2(N__20552),
            .in3(N__20006),
            .lcout(pwm_duty_input_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47350),
            .ce(N__23672),
            .sr(N__46693));
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_6_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_6_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_6_3 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_1_LC_1_6_3  (
            .in0(N__19737),
            .in1(N__20633),
            .in2(N__19031),
            .in3(N__18145),
            .lcout(pwm_duty_input_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47350),
            .ce(N__23672),
            .sr(N__46693));
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_6_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_6_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_6_4 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_2_LC_1_6_4  (
            .in0(N__18146),
            .in1(N__19030),
            .in2(N__20615),
            .in3(N__19738),
            .lcout(pwm_duty_input_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47350),
            .ce(N__23672),
            .sr(N__46693));
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_7_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_7_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_10_LC_1_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21246),
            .lcout(pwm_duty_input_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47349),
            .ce(N__23578),
            .sr(N__46703));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_1_8_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_1_8_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_1_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_1_8_1  (
            .in0(N__19489),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19510),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_1_8_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_1_8_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_1_8_2 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_1_8_2  (
            .in0(N__19685),
            .in1(N__21245),
            .in2(_gnd_net_),
            .in3(N__20057),
            .lcout(\current_shift_inst.PI_CTRL.N_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_1_8_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_1_8_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_1_8_4 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_1_8_4  (
            .in0(_gnd_net_),
            .in1(N__20197),
            .in2(_gnd_net_),
            .in3(N__20182),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_9_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_9_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_9_0  (
            .in0(_gnd_net_),
            .in1(N__19324),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_9_0_),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_9_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_9_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_9_1  (
            .in0(_gnd_net_),
            .in1(N__18197),
            .in2(_gnd_net_),
            .in3(N__18188),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_0 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_9_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_9_2  (
            .in0(_gnd_net_),
            .in1(N__18185),
            .in2(_gnd_net_),
            .in3(N__18176),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_1 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_9_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_9_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_9_3  (
            .in0(_gnd_net_),
            .in1(N__18173),
            .in2(_gnd_net_),
            .in3(N__18161),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_2 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_9_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_9_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_9_4  (
            .in0(_gnd_net_),
            .in1(N__18287),
            .in2(_gnd_net_),
            .in3(N__18158),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_3 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_9_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_9_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_9_5  (
            .in0(_gnd_net_),
            .in1(N__28796),
            .in2(N__18254),
            .in3(N__18155),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_4 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_9_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_9_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_9_6  (
            .in0(_gnd_net_),
            .in1(N__18212),
            .in2(N__28848),
            .in3(N__18152),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_5 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_9_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_9_7  (
            .in0(_gnd_net_),
            .in1(N__28800),
            .in2(N__18578),
            .in3(N__18149),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_6 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_10_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_10_0  (
            .in0(_gnd_net_),
            .in1(N__18539),
            .in2(_gnd_net_),
            .in3(N__18200),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9 ),
            .ltout(),
            .carryin(bfn_1_10_0_),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_10_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_10_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_10_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_10_1  (
            .in0(_gnd_net_),
            .in1(N__18500),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_8 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_10_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_10_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_10_2  (
            .in0(_gnd_net_),
            .in1(N__18461),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_9 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_10_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_10_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_10_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_10_3  (
            .in0(_gnd_net_),
            .in1(N__18425),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_10 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_10_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_10_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_10_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18389),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_11 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_10_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_10_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_10_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_10_5  (
            .in0(_gnd_net_),
            .in1(N__18344),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_12 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_10_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_10_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_10_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_10_6  (
            .in0(_gnd_net_),
            .in1(N__18815),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_13 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_10_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_10_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_10_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18791),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_14 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_11_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(N__18761),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_11_0_),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_11_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_11_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(N__18737),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_16 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_11_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_11_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(N__18710),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_17 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_11_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_11_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(N__18644),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_18 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_11_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18332),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_11_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_11_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_11_5  (
            .in0(N__18686),
            .in1(N__18319),
            .in2(_gnd_net_),
            .in3(N__18952),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_11_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_11_6 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_11_6  (
            .in0(N__18953),
            .in1(N__18329),
            .in2(N__18323),
            .in3(N__18685),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_axb_4_LC_1_12_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_axb_4_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_axb_4_LC_1_12_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_axb_4_LC_1_12_0  (
            .in0(_gnd_net_),
            .in1(N__18311),
            .in2(N__18302),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un3_threshold_acc_axbZ0Z_4 ),
            .ltout(),
            .carryin(bfn_1_12_0_),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_1_12_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_1_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_1_12_1  (
            .in0(_gnd_net_),
            .in1(N__18278),
            .in2(N__18266),
            .in3(N__18242),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_1_12_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_1_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_1_12_2  (
            .in0(_gnd_net_),
            .in1(N__18239),
            .in2(N__18227),
            .in3(N__18203),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_1_12_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_1_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_1_12_3  (
            .in0(_gnd_net_),
            .in1(N__18605),
            .in2(N__18593),
            .in3(N__18566),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_1_12_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_1_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_1_12_4  (
            .in0(_gnd_net_),
            .in1(N__18563),
            .in2(N__18551),
            .in3(N__18530),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_1_12_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_1_12_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_1_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_1_12_5  (
            .in0(_gnd_net_),
            .in1(N__18527),
            .in2(N__18515),
            .in3(N__18491),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_1_12_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_1_12_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_1_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_1_12_6  (
            .in0(_gnd_net_),
            .in1(N__18488),
            .in2(N__18476),
            .in3(N__18452),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_1_12_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_1_12_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_1_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_1_12_7  (
            .in0(_gnd_net_),
            .in1(N__18449),
            .in2(N__18437),
            .in3(N__18416),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_1_13_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_1_13_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_1_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_1_13_0  (
            .in0(_gnd_net_),
            .in1(N__18413),
            .in2(N__18401),
            .in3(N__18377),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0 ),
            .ltout(),
            .carryin(bfn_1_13_0_),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_1_13_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_1_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_1_13_1  (
            .in0(_gnd_net_),
            .in1(N__18374),
            .in2(N__18359),
            .in3(N__18335),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_1_13_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_1_13_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_1_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_1_13_2  (
            .in0(_gnd_net_),
            .in1(N__18673),
            .in2(N__18830),
            .in3(N__18806),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_1_13_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_1_13_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_1_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_1_13_3  (
            .in0(_gnd_net_),
            .in1(N__18803),
            .in2(N__18687),
            .in3(N__18779),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_1_13_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_1_13_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_1_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_1_13_4  (
            .in0(_gnd_net_),
            .in1(N__18677),
            .in2(N__18776),
            .in3(N__18752),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_1_13_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_1_13_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_1_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_1_13_5  (
            .in0(_gnd_net_),
            .in1(N__18749),
            .in2(N__18688),
            .in3(N__18728),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_1_13_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_1_13_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_1_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_1_13_6  (
            .in0(_gnd_net_),
            .in1(N__18681),
            .in2(N__18725),
            .in3(N__18701),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_1_13_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_1_13_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_1_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_1_13_7  (
            .in0(_gnd_net_),
            .in1(N__18698),
            .in2(N__18689),
            .in3(N__18635),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_1_14_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_1_14_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_1_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_1_14_0  (
            .in0(N__18632),
            .in1(N__18623),
            .in2(_gnd_net_),
            .in3(N__18614),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.N_110_i_i_LC_1_29_3 .C_ON=1'b0;
    defparam \current_shift_inst.N_110_i_i_LC_1_29_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.N_110_i_i_LC_1_29_3 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \current_shift_inst.N_110_i_i_LC_1_29_3  (
            .in0(N__46778),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34564),
            .lcout(N_110_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un7_start_stop_LC_1_30_1 .C_ON=1'b0;
    defparam \current_shift_inst.un7_start_stop_LC_1_30_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un7_start_stop_LC_1_30_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \current_shift_inst.un7_start_stop_LC_1_30_1  (
            .in0(N__46779),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34568),
            .lcout(un7_start_stop),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNILM9T_5_LC_2_5_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNILM9T_5_LC_2_5_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNILM9T_5_LC_2_5_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNILM9T_5_LC_2_5_3  (
            .in0(N__19116),
            .in1(N__19137),
            .in2(N__19099),
            .in3(N__19062),
            .lcout(\current_shift_inst.PI_CTRL.m14_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNIDE9T_3_LC_2_5_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNIDE9T_3_LC_2_5_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNIDE9T_3_LC_2_5_7 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNIDE9T_3_LC_2_5_7  (
            .in0(N__19003),
            .in1(N__19138),
            .in2(N__19121),
            .in3(N__18847),
            .lcout(\current_shift_inst.PI_CTRL.m7_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNIVCED1_7_LC_2_6_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNIVCED1_7_LC_2_6_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNIVCED1_7_LC_2_6_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNIVCED1_7_LC_2_6_1  (
            .in0(N__19095),
            .in1(N__18886),
            .in2(N__19073),
            .in3(N__19063),
            .lcout(i8_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_6_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_6_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_6_4 .LUT_INIT=16'b0101010100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_6_4  (
            .in0(N__21269),
            .in1(N__20548),
            .in2(_gnd_net_),
            .in3(N__20055),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_6_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_6_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_6_5 .LUT_INIT=16'b0101010100010000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_6_5  (
            .in0(N__20590),
            .in1(N__19681),
            .in2(N__19034),
            .in3(N__19726),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNIUU8T_0_LC_2_6_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNIUU8T_0_LC_2_6_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNIUU8T_0_LC_2_6_6 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNIUU8T_0_LC_2_6_6  (
            .in0(N__19016),
            .in1(N__19004),
            .in2(N__18986),
            .in3(N__18971),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.N_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNIK2D32_4_LC_2_6_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNIK2D32_4_LC_2_6_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNIK2D32_4_LC_2_6_7 .LUT_INIT=16'b0010001000100000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNIK2D32_4_LC_2_6_7  (
            .in0(N__18959),
            .in1(N__18885),
            .in2(N__18851),
            .in3(N__18848),
            .lcout(N_28_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_2_7_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_2_7_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_2_7_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_2_7_0  (
            .in0(_gnd_net_),
            .in1(N__19277),
            .in2(_gnd_net_),
            .in3(N__19289),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_0 ),
            .ltout(),
            .carryin(bfn_2_7_0_),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_2_7_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_2_7_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_2_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_2_7_1  (
            .in0(_gnd_net_),
            .in1(N__19259),
            .in2(_gnd_net_),
            .in3(N__19271),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_0 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_2_7_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_2_7_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_2_7_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_2_7_2  (
            .in0(_gnd_net_),
            .in1(N__19241),
            .in2(_gnd_net_),
            .in3(N__19253),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_1 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_2_7_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_2_7_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_2_7_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_2_7_3  (
            .in0(_gnd_net_),
            .in1(N__19223),
            .in2(_gnd_net_),
            .in3(N__19235),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_2 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_2_7_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_2_7_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_2_7_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_2_7_4  (
            .in0(_gnd_net_),
            .in1(N__19205),
            .in2(_gnd_net_),
            .in3(N__19217),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_3 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_2_7_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_2_7_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_2_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_2_7_5  (
            .in0(_gnd_net_),
            .in1(N__19187),
            .in2(_gnd_net_),
            .in3(N__19199),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_4 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_2_7_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_2_7_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_2_7_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_2_7_6  (
            .in0(_gnd_net_),
            .in1(N__19169),
            .in2(_gnd_net_),
            .in3(N__19181),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_5 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_2_7_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_2_7_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_2_7_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_2_7_7  (
            .in0(_gnd_net_),
            .in1(N__19151),
            .in2(_gnd_net_),
            .in3(N__19163),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_6 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_2_8_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_2_8_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_2_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_2_8_0  (
            .in0(_gnd_net_),
            .in1(N__19355),
            .in2(_gnd_net_),
            .in3(N__19367),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_8 ),
            .ltout(),
            .carryin(bfn_2_8_0_),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_2_8_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_2_8_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_2_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_2_8_1  (
            .in0(_gnd_net_),
            .in1(N__19337),
            .in2(_gnd_net_),
            .in3(N__19349),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_8 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_2_8_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_2_8_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_2_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_2_8_2  (
            .in0(_gnd_net_),
            .in1(N__19485),
            .in2(_gnd_net_),
            .in3(N__19331),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_9 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_2_8_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_2_8_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_2_8_3 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_2_8_3  (
            .in0(N__20132),
            .in1(N__19328),
            .in2(_gnd_net_),
            .in3(N__19307),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_10 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_2_8_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_2_8_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_2_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_2_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19780),
            .in3(N__19304),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_11 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_2_8_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_2_8_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_2_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_2_8_5  (
            .in0(_gnd_net_),
            .in1(N__19537),
            .in2(_gnd_net_),
            .in3(N__19301),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_12 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_2_8_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_2_8_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_2_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_2_8_6  (
            .in0(_gnd_net_),
            .in1(N__20178),
            .in2(_gnd_net_),
            .in3(N__19298),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_13 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_2_8_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_2_8_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_2_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_2_8_7  (
            .in0(_gnd_net_),
            .in1(N__19443),
            .in2(_gnd_net_),
            .in3(N__19295),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_14 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_2_9_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_2_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_2_9_0  (
            .in0(_gnd_net_),
            .in1(N__19566),
            .in2(_gnd_net_),
            .in3(N__19292),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_2_9_0_),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_2_9_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_2_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_2_9_1  (
            .in0(_gnd_net_),
            .in1(N__19399),
            .in2(_gnd_net_),
            .in3(N__19454),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_16 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_2_9_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_2_9_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_2_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_2_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19628),
            .in3(N__19451),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_17 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_2_9_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_2_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_2_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19448),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_9_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_9_4 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_9_4  (
            .in0(_gnd_net_),
            .in1(N__19795),
            .in2(_gnd_net_),
            .in3(N__19779),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_9_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_9_6 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_9_6  (
            .in0(_gnd_net_),
            .in1(N__19588),
            .in2(_gnd_net_),
            .in3(N__19567),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_9_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_9_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_9_7  (
            .in0(N__19445),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19426),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_10_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_10_0 .LUT_INIT=16'b1010010111001100;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_10_0  (
            .in0(N__19444),
            .in1(N__19427),
            .in2(N__19415),
            .in3(N__20135),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_10_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_10_2  (
            .in0(N__19403),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19387),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ),
            .ltout(\pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_10_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_10_3 .LUT_INIT=16'b1110010001001110;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_10_3  (
            .in0(N__20136),
            .in1(N__19388),
            .in2(N__19376),
            .in3(N__19373),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_10_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_10_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_10_4 .LUT_INIT=16'b1010010111001100;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_10_4  (
            .in0(N__19538),
            .in1(N__19552),
            .in2(N__19640),
            .in3(N__20133),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_10_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_10_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_10_5  (
            .in0(N__19609),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19627),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ),
            .ltout(\pwm_generator_inst.un15_threshold_acc_1_axb_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_10_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_10_6 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_10_6  (
            .in0(N__19613),
            .in1(N__20137),
            .in2(N__19598),
            .in3(N__19595),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_10_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_10_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_10_7 .LUT_INIT=16'b1110010001001110;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_10_7  (
            .in0(N__20134),
            .in1(N__19589),
            .in2(N__19577),
            .in3(N__19568),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_9_LC_2_11_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_9_LC_2_11_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_9_LC_2_11_0 .LUT_INIT=16'b0011000001010000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_9_LC_2_11_0  (
            .in0(N__20702),
            .in1(N__20768),
            .in2(N__19895),
            .in3(N__20854),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47339),
            .ce(),
            .sr(N__46719));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_11_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_11_7  (
            .in0(N__19536),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19553),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_13_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_13_0 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_13_0  (
            .in0(N__19517),
            .in1(N__19493),
            .in2(N__19469),
            .in3(N__20094),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_2_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_2_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_2_13_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_2_LC_2_13_3  (
            .in0(N__44205),
            .in1(N__40328),
            .in2(N__34114),
            .in3(N__43912),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47330),
            .ce(N__31224),
            .sr(N__46727));
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_2_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_2_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_2_13_5 .LUT_INIT=16'b1111111010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_1_LC_2_13_5  (
            .in0(N__44204),
            .in1(N__40327),
            .in2(N__41276),
            .in3(N__43911),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47330),
            .ce(N__31224),
            .sr(N__46727));
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_2_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_2_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_2_13_6 .LUT_INIT=16'b1110111011101100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_3_LC_2_13_6  (
            .in0(N__43913),
            .in1(N__44206),
            .in2(N__40343),
            .in3(N__35522),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47330),
            .ce(N__31224),
            .sr(N__46727));
    defparam \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_2_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_2_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_2_13_7 .LUT_INIT=16'b0000001000000011;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_2_13_7  (
            .in0(N__34169),
            .in1(N__40326),
            .in2(N__44207),
            .in3(N__43910),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ1Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47330),
            .ce(N__31224),
            .sr(N__46727));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_14_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_14_0 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_14_0  (
            .in0(N__19802),
            .in1(N__19784),
            .in2(N__19757),
            .in3(N__20101),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_10_LC_2_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_10_LC_2_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_10_LC_2_15_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_10_LC_2_15_2  (
            .in0(N__20258),
            .in1(N__20228),
            .in2(N__20024),
            .in3(N__20222),
            .lcout(\current_shift_inst.PI_CTRL.N_178 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_3_6_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_3_6_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_3_6_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_3_6_2  (
            .in0(N__20583),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20540),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.N_98_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_3_6_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_3_6_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_3_6_3 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_3_6_3  (
            .in0(N__19882),
            .in1(N__21258),
            .in2(N__19742),
            .in3(N__20000),
            .lcout(\current_shift_inst.PI_CTRL.N_96 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_3_6_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_3_6_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_3_6_6 .LUT_INIT=16'b0000111100000111;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_3_6_6  (
            .in0(N__20541),
            .in1(N__20056),
            .in2(N__21268),
            .in3(N__19713),
            .lcout(\current_shift_inst.PI_CTRL.N_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_1_LC_3_7_0.C_ON=1'b0;
    defparam counter_1_LC_3_7_0.SEQ_MODE=4'b1010;
    defparam counter_1_LC_3_7_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 counter_1_LC_3_7_0 (
            .in0(_gnd_net_),
            .in1(N__21466),
            .in2(_gnd_net_),
            .in3(N__21427),
            .lcout(counterZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47348),
            .ce(),
            .sr(N__46684));
    defparam counter_RNIM6001_12_LC_3_7_1.C_ON=1'b0;
    defparam counter_RNIM6001_12_LC_3_7_1.SEQ_MODE=4'b0000;
    defparam counter_RNIM6001_12_LC_3_7_1.LUT_INIT=16'b0000000100000000;
    LogicCell40 counter_RNIM6001_12_LC_3_7_1 (
            .in0(N__20431),
            .in1(N__20272),
            .in2(N__20291),
            .in3(N__20416),
            .lcout(un2_counter_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNII76D_3_LC_3_7_3.C_ON=1'b0;
    defparam counter_RNII76D_3_LC_3_7_3.SEQ_MODE=4'b0000;
    defparam counter_RNII76D_3_LC_3_7_3.LUT_INIT=16'b0000000000000001;
    LogicCell40 counter_RNII76D_3_LC_3_7_3 (
            .in0(N__20326),
            .in1(N__20341),
            .in2(N__20312),
            .in3(N__20356),
            .lcout(un2_counter_7),
            .ltout(un2_counter_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_0_LC_3_7_4.C_ON=1'b0;
    defparam counter_0_LC_3_7_4.SEQ_MODE=4'b1010;
    defparam counter_0_LC_3_7_4.LUT_INIT=16'b0001001100110011;
    LogicCell40 counter_0_LC_3_7_4 (
            .in0(N__21667),
            .in1(N__21426),
            .in2(N__19859),
            .in3(N__21714),
            .lcout(counterZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47348),
            .ce(),
            .sr(N__46684));
    defparam \pwm_generator_inst.threshold_ACC_7_LC_3_8_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_7_LC_3_8_1 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_7_LC_3_8_1 .LUT_INIT=16'b1111111110101100;
    LogicCell40 \pwm_generator_inst.threshold_ACC_7_LC_3_8_1  (
            .in0(N__20777),
            .in1(N__20721),
            .in2(N__20859),
            .in3(N__19937),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47346),
            .ce(),
            .sr(N__46694));
    defparam counter_12_LC_3_8_2.C_ON=1'b0;
    defparam counter_12_LC_3_8_2.SEQ_MODE=4'b1010;
    defparam counter_12_LC_3_8_2.LUT_INIT=16'b0010101010101010;
    LogicCell40 counter_12_LC_3_8_2 (
            .in0(N__20402),
            .in1(N__21711),
            .in2(N__21674),
            .in3(N__21619),
            .lcout(counterZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47346),
            .ce(),
            .sr(N__46694));
    defparam \pwm_generator_inst.threshold_ACC_2_LC_3_8_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_2_LC_3_8_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_2_LC_3_8_7 .LUT_INIT=16'b0101001100000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_2_LC_3_8_7  (
            .in0(N__20776),
            .in1(N__20720),
            .in2(N__20858),
            .in3(N__19820),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47346),
            .ce(),
            .sr(N__46694));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_3_9_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_3_9_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_3_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_3_9_0  (
            .in0(_gnd_net_),
            .in1(N__19856),
            .in2(N__20150),
            .in3(N__20149),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(bfn_3_9_0_),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_3_9_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_3_9_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_3_9_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_3_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19844),
            .in3(N__19835),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_0 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_3_9_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_3_9_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_3_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_3_9_2  (
            .in0(_gnd_net_),
            .in1(N__19832),
            .in2(_gnd_net_),
            .in3(N__19814),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_1 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_3_9_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_3_9_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_3_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_3_9_3  (
            .in0(_gnd_net_),
            .in1(N__19811),
            .in2(_gnd_net_),
            .in3(N__19805),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_2 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_3_9_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_3_9_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_3_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_3_9_4  (
            .in0(_gnd_net_),
            .in1(N__20066),
            .in2(_gnd_net_),
            .in3(N__19964),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_3 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_3_9_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_3_9_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_3_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_3_9_5  (
            .in0(_gnd_net_),
            .in1(N__19961),
            .in2(_gnd_net_),
            .in3(N__19955),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_4 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_3_9_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_3_9_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_3_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_3_9_6  (
            .in0(_gnd_net_),
            .in1(N__19952),
            .in2(_gnd_net_),
            .in3(N__19946),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_5 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_3_9_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_3_9_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_3_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_3_9_7  (
            .in0(_gnd_net_),
            .in1(N__19943),
            .in2(_gnd_net_),
            .in3(N__19931),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_6 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_3_10_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_3_10_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_3_10_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_3_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19928),
            .in3(N__19919),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(bfn_3_10_0_),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_3_10_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_3_10_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_3_10_1 .LUT_INIT=16'b1000011101111000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_3_10_1  (
            .in0(N__20139),
            .in1(N__19916),
            .in2(N__19910),
            .in3(N__19898),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_3_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_3_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_3_10_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_3_10_2  (
            .in0(N__20494),
            .in1(N__20467),
            .in2(N__21025),
            .in3(N__19865),
            .lcout(\current_shift_inst.PI_CTRL.N_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIU1LD_7_LC_3_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIU1LD_7_LC_3_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIU1LD_7_LC_3_10_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIU1LD_7_LC_3_10_3  (
            .in0(_gnd_net_),
            .in1(N__20980),
            .in2(_gnd_net_),
            .in3(N__21061),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_3_10_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_3_10_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_3_10_4 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_3_10_4  (
            .in0(N__20204),
            .in1(N__20186),
            .in2(N__20162),
            .in3(N__20138),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQTKD_5_LC_3_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQTKD_5_LC_3_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQTKD_5_LC_3_11_4 .LUT_INIT=16'b0111011101110111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIQTKD_5_LC_3_11_4  (
            .in0(N__21057),
            .in1(N__20493),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_3_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_3_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_3_11_5 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_3_11_5  (
            .in0(N__20976),
            .in1(N__21024),
            .in2(N__20060),
            .in3(N__20463),
            .lcout(\current_shift_inst.PI_CTRL.N_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMJ62_12_LC_3_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMJ62_12_LC_3_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMJ62_12_LC_3_14_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMJ62_12_LC_3_14_1  (
            .in0(_gnd_net_),
            .in1(N__21073),
            .in2(_gnd_net_),
            .in3(N__20920),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_9_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIU8H5_14_LC_3_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIU8H5_14_LC_3_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIU8H5_14_LC_3_14_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIU8H5_14_LC_3_14_2  (
            .in0(N__21359),
            .in1(N__21388),
            .in2(N__20027),
            .in3(N__20887),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIEAE4_15_LC_3_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIEAE4_15_LC_3_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIEAE4_15_LC_3_14_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIEAE4_15_LC_3_14_3  (
            .in0(N__20873),
            .in1(N__21107),
            .in2(N__21094),
            .in3(N__21074),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFBE4_19_LC_3_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFBE4_19_LC_3_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFBE4_19_LC_3_14_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIFBE4_19_LC_3_14_5  (
            .in0(N__21121),
            .in1(N__21106),
            .in2(N__21095),
            .in3(N__21136),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_3_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_3_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_3_14_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_3_14_6  (
            .in0(N__20237),
            .in1(N__20015),
            .in2(N__20009),
            .in3(N__20243),
            .lcout(\current_shift_inst.PI_CTRL.N_118 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPM62_13_LC_3_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPM62_13_LC_3_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPM62_13_LC_3_15_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIPM62_13_LC_3_15_0  (
            .in0(_gnd_net_),
            .in1(N__21370),
            .in2(_gnd_net_),
            .in3(N__20905),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRMD4_17_LC_3_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRMD4_17_LC_3_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRMD4_17_LC_3_15_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIRMD4_17_LC_3_15_1  (
            .in0(N__21389),
            .in1(N__21154),
            .in2(N__21358),
            .in3(N__21167),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQJB4_15_LC_3_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQJB4_15_LC_3_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQJB4_15_LC_3_15_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIQJB4_15_LC_3_15_2  (
            .in0(N__21166),
            .in1(N__21178),
            .in2(N__21155),
            .in3(N__20872),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIKAQ8_27_LC_3_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIKAQ8_27_LC_3_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIKAQ8_27_LC_3_15_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIKAQ8_27_LC_3_15_3  (
            .in0(N__21320),
            .in1(N__21335),
            .in2(N__20252),
            .in3(N__20249),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNID9E4_10_LC_3_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNID9E4_10_LC_3_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNID9E4_10_LC_3_15_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNID9E4_10_LC_3_15_4  (
            .in0(N__21304),
            .in1(N__20935),
            .in2(N__21290),
            .in3(N__20947),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPL52_13_LC_3_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPL52_13_LC_3_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPL52_13_LC_3_15_5 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIPL52_13_LC_3_15_5  (
            .in0(N__20906),
            .in1(_gnd_net_),
            .in2(N__21182),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISHP8_10_LC_3_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISHP8_10_LC_3_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISHP8_10_LC_3_15_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISHP8_10_LC_3_15_6  (
            .in0(N__20210),
            .in1(N__20936),
            .in2(N__20231),
            .in3(N__20948),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI9LI5_19_LC_3_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI9LI5_19_LC_3_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI9LI5_19_LC_3_15_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI9LI5_19_LC_3_15_7  (
            .in0(N__21371),
            .in1(N__20216),
            .in2(N__21140),
            .in3(N__21122),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1082_27_LC_3_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1082_27_LC_3_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1082_27_LC_3_16_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI1082_27_LC_3_16_0  (
            .in0(_gnd_net_),
            .in1(N__21319),
            .in2(_gnd_net_),
            .in3(N__21334),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIEE4_12_LC_3_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIEE4_12_LC_3_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIEE4_12_LC_3_16_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIIEE4_12_LC_3_16_7  (
            .in0(N__20924),
            .in1(N__21289),
            .in2(N__20894),
            .in3(N__21305),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_counter_cry_1_c_LC_4_7_0.C_ON=1'b1;
    defparam un5_counter_cry_1_c_LC_4_7_0.SEQ_MODE=4'b0000;
    defparam un5_counter_cry_1_c_LC_4_7_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_counter_cry_1_c_LC_4_7_0 (
            .in0(_gnd_net_),
            .in1(N__21425),
            .in2(N__21467),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_7_0_),
            .carryout(un5_counter_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_2_LC_4_7_1.C_ON=1'b1;
    defparam counter_2_LC_4_7_1.SEQ_MODE=4'b1010;
    defparam counter_2_LC_4_7_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_2_LC_4_7_1 (
            .in0(_gnd_net_),
            .in1(N__21443),
            .in2(_gnd_net_),
            .in3(N__20360),
            .lcout(counterZ0Z_2),
            .ltout(),
            .carryin(un5_counter_cry_1),
            .carryout(un5_counter_cry_2),
            .clk(N__47347),
            .ce(),
            .sr(N__46678));
    defparam counter_3_LC_4_7_2.C_ON=1'b1;
    defparam counter_3_LC_4_7_2.SEQ_MODE=4'b1010;
    defparam counter_3_LC_4_7_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_3_LC_4_7_2 (
            .in0(_gnd_net_),
            .in1(N__20357),
            .in2(_gnd_net_),
            .in3(N__20345),
            .lcout(counterZ0Z_3),
            .ltout(),
            .carryin(un5_counter_cry_2),
            .carryout(un5_counter_cry_3),
            .clk(N__47347),
            .ce(),
            .sr(N__46678));
    defparam counter_4_LC_4_7_3.C_ON=1'b1;
    defparam counter_4_LC_4_7_3.SEQ_MODE=4'b1010;
    defparam counter_4_LC_4_7_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_4_LC_4_7_3 (
            .in0(_gnd_net_),
            .in1(N__20342),
            .in2(_gnd_net_),
            .in3(N__20330),
            .lcout(counterZ0Z_4),
            .ltout(),
            .carryin(un5_counter_cry_3),
            .carryout(un5_counter_cry_4),
            .clk(N__47347),
            .ce(),
            .sr(N__46678));
    defparam counter_5_LC_4_7_4.C_ON=1'b1;
    defparam counter_5_LC_4_7_4.SEQ_MODE=4'b1010;
    defparam counter_5_LC_4_7_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_5_LC_4_7_4 (
            .in0(_gnd_net_),
            .in1(N__20327),
            .in2(_gnd_net_),
            .in3(N__20315),
            .lcout(counterZ0Z_5),
            .ltout(),
            .carryin(un5_counter_cry_4),
            .carryout(un5_counter_cry_5),
            .clk(N__47347),
            .ce(),
            .sr(N__46678));
    defparam counter_6_LC_4_7_5.C_ON=1'b1;
    defparam counter_6_LC_4_7_5.SEQ_MODE=4'b1010;
    defparam counter_6_LC_4_7_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_6_LC_4_7_5 (
            .in0(_gnd_net_),
            .in1(N__20311),
            .in2(_gnd_net_),
            .in3(N__20297),
            .lcout(counterZ0Z_6),
            .ltout(),
            .carryin(un5_counter_cry_5),
            .carryout(un5_counter_cry_6),
            .clk(N__47347),
            .ce(),
            .sr(N__46678));
    defparam counter_RNO_0_7_LC_4_7_6.C_ON=1'b1;
    defparam counter_RNO_0_7_LC_4_7_6.SEQ_MODE=4'b0000;
    defparam counter_RNO_0_7_LC_4_7_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_RNO_0_7_LC_4_7_6 (
            .in0(_gnd_net_),
            .in1(N__21479),
            .in2(_gnd_net_),
            .in3(N__20294),
            .lcout(counter_RNO_0Z0Z_7),
            .ltout(),
            .carryin(un5_counter_cry_6),
            .carryout(un5_counter_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_8_LC_4_7_7.C_ON=1'b1;
    defparam counter_8_LC_4_7_7.SEQ_MODE=4'b1010;
    defparam counter_8_LC_4_7_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_8_LC_4_7_7 (
            .in0(_gnd_net_),
            .in1(N__20290),
            .in2(_gnd_net_),
            .in3(N__20276),
            .lcout(counterZ0Z_8),
            .ltout(),
            .carryin(un5_counter_cry_7),
            .carryout(un5_counter_cry_8),
            .clk(N__47347),
            .ce(),
            .sr(N__46678));
    defparam counter_9_LC_4_8_0.C_ON=1'b1;
    defparam counter_9_LC_4_8_0.SEQ_MODE=4'b1010;
    defparam counter_9_LC_4_8_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_9_LC_4_8_0 (
            .in0(_gnd_net_),
            .in1(N__20273),
            .in2(_gnd_net_),
            .in3(N__20261),
            .lcout(counterZ0Z_9),
            .ltout(),
            .carryin(bfn_4_8_0_),
            .carryout(un5_counter_cry_9),
            .clk(N__47344),
            .ce(),
            .sr(N__46685));
    defparam counter_RNO_0_10_LC_4_8_1.C_ON=1'b1;
    defparam counter_RNO_0_10_LC_4_8_1.SEQ_MODE=4'b0000;
    defparam counter_RNO_0_10_LC_4_8_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_RNO_0_10_LC_4_8_1 (
            .in0(_gnd_net_),
            .in1(N__21593),
            .in2(_gnd_net_),
            .in3(N__20435),
            .lcout(counter_RNO_0Z0Z_10),
            .ltout(),
            .carryin(un5_counter_cry_9),
            .carryout(un5_counter_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_11_LC_4_8_2.C_ON=1'b1;
    defparam counter_11_LC_4_8_2.SEQ_MODE=4'b1010;
    defparam counter_11_LC_4_8_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_11_LC_4_8_2 (
            .in0(_gnd_net_),
            .in1(N__20432),
            .in2(_gnd_net_),
            .in3(N__20420),
            .lcout(counterZ0Z_11),
            .ltout(),
            .carryin(un5_counter_cry_10),
            .carryout(un5_counter_cry_11),
            .clk(N__47344),
            .ce(),
            .sr(N__46685));
    defparam counter_RNO_0_12_LC_4_8_3.C_ON=1'b0;
    defparam counter_RNO_0_12_LC_4_8_3.SEQ_MODE=4'b0000;
    defparam counter_RNO_0_12_LC_4_8_3.LUT_INIT=16'b0011001111001100;
    LogicCell40 counter_RNO_0_12_LC_4_8_3 (
            .in0(_gnd_net_),
            .in1(N__20417),
            .in2(_gnd_net_),
            .in3(N__20405),
            .lcout(counter_RNO_0Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_0_LC_4_9_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_0_LC_4_9_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_0_LC_4_9_0 .LUT_INIT=16'b0100000001001100;
    LogicCell40 \pwm_generator_inst.threshold_ACC_0_LC_4_9_0  (
            .in0(N__20772),
            .in1(N__20396),
            .in2(N__20861),
            .in3(N__20719),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47340),
            .ce(),
            .sr(N__46695));
    defparam \pwm_generator_inst.threshold_ACC_4_LC_4_9_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_4_LC_4_9_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_4_LC_4_9_1 .LUT_INIT=16'b0010011100000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_4_LC_4_9_1  (
            .in0(N__20847),
            .in1(N__20775),
            .in2(N__20726),
            .in3(N__20390),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47340),
            .ce(),
            .sr(N__46695));
    defparam \pwm_generator_inst.threshold_ACC_1_LC_4_9_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_1_LC_4_9_3 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_1_LC_4_9_3 .LUT_INIT=16'b1111111111011000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_1_LC_4_9_3  (
            .in0(N__20846),
            .in1(N__20774),
            .in2(N__20725),
            .in3(N__20384),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47340),
            .ce(),
            .sr(N__46695));
    defparam \pwm_generator_inst.threshold_ACC_3_LC_4_9_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_3_LC_4_9_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_3_LC_4_9_6 .LUT_INIT=16'b0101001100000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_3_LC_4_9_6  (
            .in0(N__20773),
            .in1(N__20712),
            .in2(N__20860),
            .in3(N__20378),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47340),
            .ce(),
            .sr(N__46695));
    defparam \pwm_generator_inst.threshold_ACC_6_LC_4_10_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_6_LC_4_10_2 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_6_LC_4_10_2 .LUT_INIT=16'b1111111111011000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_6_LC_4_10_2  (
            .in0(N__20855),
            .in1(N__20770),
            .in2(N__20722),
            .in3(N__20372),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47336),
            .ce(),
            .sr(N__46704));
    defparam \pwm_generator_inst.threshold_ACC_5_LC_4_10_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_5_LC_4_10_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_5_LC_4_10_5 .LUT_INIT=16'b0100011100000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_5_LC_4_10_5  (
            .in0(N__20769),
            .in1(N__20857),
            .in2(N__20724),
            .in3(N__20366),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47336),
            .ce(),
            .sr(N__46704));
    defparam \pwm_generator_inst.threshold_ACC_8_LC_4_10_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_8_LC_4_10_6 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_8_LC_4_10_6 .LUT_INIT=16'b1111111111011000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_8_LC_4_10_6  (
            .in0(N__20856),
            .in1(N__20771),
            .in2(N__20723),
            .in3(N__20657),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47336),
            .ce(),
            .sr(N__46704));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_4_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_4_13_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_4_13_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_0_LC_4_13_0  (
            .in0(_gnd_net_),
            .in1(N__23888),
            .in2(N__21530),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ),
            .ltout(),
            .carryin(bfn_4_13_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ),
            .clk(N__47315),
            .ce(N__23649),
            .sr(N__46720));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_4_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_4_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_4_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_LC_4_13_1  (
            .in0(_gnd_net_),
            .in1(N__23834),
            .in2(N__21575),
            .in3(N__20618),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .clk(N__47315),
            .ce(N__23649),
            .sr(N__46720));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_4_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_4_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_4_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_2_LC_4_13_2  (
            .in0(_gnd_net_),
            .in1(N__23783),
            .in2(N__21785),
            .in3(N__20597),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .clk(N__47315),
            .ce(N__23649),
            .sr(N__46720));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_4_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_4_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_4_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_3_LC_4_13_3  (
            .in0(_gnd_net_),
            .in1(N__23711),
            .in2(N__21758),
            .in3(N__20555),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .clk(N__47315),
            .ce(N__23649),
            .sr(N__46720));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_4_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_4_13_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_4_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_4_LC_4_13_4  (
            .in0(_gnd_net_),
            .in1(N__23497),
            .in2(N__21521),
            .in3(N__20504),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .clk(N__47315),
            .ce(N__23649),
            .sr(N__46720));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_4_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_4_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_4_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_5_LC_4_13_5  (
            .in0(_gnd_net_),
            .in1(N__24476),
            .in2(N__21539),
            .in3(N__20474),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .clk(N__47315),
            .ce(N__23649),
            .sr(N__46720));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_4_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_4_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_4_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_6_LC_4_13_6  (
            .in0(_gnd_net_),
            .in1(N__24398),
            .in2(N__21767),
            .in3(N__20438),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .clk(N__47315),
            .ce(N__23649),
            .sr(N__46720));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_4_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_4_13_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_4_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_7_LC_4_13_7  (
            .in0(_gnd_net_),
            .in1(N__24302),
            .in2(N__22067),
            .in3(N__21032),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .clk(N__47315),
            .ce(N__23649),
            .sr(N__46720));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_4_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_4_14_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_4_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_8_LC_4_14_0  (
            .in0(_gnd_net_),
            .in1(N__24260),
            .in2(N__21776),
            .in3(N__20990),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ),
            .ltout(),
            .carryin(bfn_4_14_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .clk(N__47303),
            .ce(N__23637),
            .sr(N__46724));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_4_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_4_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_4_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_9_LC_4_14_1  (
            .in0(_gnd_net_),
            .in1(N__24197),
            .in2(N__21551),
            .in3(N__20951),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .clk(N__47303),
            .ce(N__23637),
            .sr(N__46724));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_4_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_4_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_4_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_10_LC_4_14_2  (
            .in0(_gnd_net_),
            .in1(N__24126),
            .in2(N__21734),
            .in3(N__20939),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .clk(N__47303),
            .ce(N__23637),
            .sr(N__46724));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_4_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_4_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_4_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_11_LC_4_14_3  (
            .in0(_gnd_net_),
            .in1(N__21560),
            .in2(N__24064),
            .in3(N__20927),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .clk(N__47303),
            .ce(N__23637),
            .sr(N__46724));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_4_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_4_14_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_4_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_12_LC_4_14_4  (
            .in0(_gnd_net_),
            .in1(N__23989),
            .in2(N__21497),
            .in3(N__20909),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .clk(N__47303),
            .ce(N__23637),
            .sr(N__46724));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_4_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_4_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_4_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_13_LC_4_14_5  (
            .in0(_gnd_net_),
            .in1(N__21725),
            .in2(N__24983),
            .in3(N__20897),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .clk(N__47303),
            .ce(N__23637),
            .sr(N__46724));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_4_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_4_14_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_4_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_14_LC_4_14_6  (
            .in0(_gnd_net_),
            .in1(N__21836),
            .in2(N__24887),
            .in3(N__20876),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .clk(N__47303),
            .ce(N__23637),
            .sr(N__46724));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_4_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_4_14_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_4_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_15_LC_4_14_7  (
            .in0(_gnd_net_),
            .in1(N__21749),
            .in2(N__24836),
            .in3(N__21185),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .clk(N__47303),
            .ce(N__23637),
            .sr(N__46724));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_4_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_4_15_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_4_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_16_LC_4_15_0  (
            .in0(_gnd_net_),
            .in1(N__24754),
            .in2(N__21800),
            .in3(N__21170),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ),
            .ltout(),
            .carryin(bfn_4_15_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .clk(N__47294),
            .ce(N__23676),
            .sr(N__46728));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_4_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_4_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_4_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_17_LC_4_15_1  (
            .in0(_gnd_net_),
            .in1(N__24683),
            .in2(N__21512),
            .in3(N__21158),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .clk(N__47294),
            .ce(N__23676),
            .sr(N__46728));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_4_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_4_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_4_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_18_LC_4_15_2  (
            .in0(_gnd_net_),
            .in1(N__21938),
            .in2(N__24620),
            .in3(N__21143),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .clk(N__47294),
            .ce(N__23676),
            .sr(N__46728));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_4_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_4_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_4_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_19_LC_4_15_3  (
            .in0(_gnd_net_),
            .in1(N__24539),
            .in2(N__21743),
            .in3(N__21125),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .clk(N__47294),
            .ce(N__23676),
            .sr(N__46728));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_4_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_4_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_4_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_20_LC_4_15_4  (
            .in0(_gnd_net_),
            .in1(N__21830),
            .in2(N__25469),
            .in3(N__21110),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .clk(N__47294),
            .ce(N__23676),
            .sr(N__46728));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_4_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_4_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_4_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_21_LC_4_15_5  (
            .in0(_gnd_net_),
            .in1(N__21791),
            .in2(N__25403),
            .in3(N__21098),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .clk(N__47294),
            .ce(N__23676),
            .sr(N__46728));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_4_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_4_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_4_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_22_LC_4_15_6  (
            .in0(_gnd_net_),
            .in1(N__25322),
            .in2(N__21923),
            .in3(N__21077),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .clk(N__47294),
            .ce(N__23676),
            .sr(N__46728));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_4_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_4_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_4_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_23_LC_4_15_7  (
            .in0(_gnd_net_),
            .in1(N__25259),
            .in2(N__21932),
            .in3(N__21065),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .clk(N__47294),
            .ce(N__23676),
            .sr(N__46728));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_4_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_4_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_4_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_24_LC_4_16_0  (
            .in0(_gnd_net_),
            .in1(N__21914),
            .in2(N__25184),
            .in3(N__21374),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ),
            .ltout(),
            .carryin(bfn_4_16_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .clk(N__47286),
            .ce(N__23673),
            .sr(N__46731));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_4_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_4_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_4_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_25_LC_4_16_1  (
            .in0(_gnd_net_),
            .in1(N__25106),
            .in2(N__21906),
            .in3(N__21362),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .clk(N__47286),
            .ce(N__23673),
            .sr(N__46731));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_4_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_4_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_4_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_26_LC_4_16_2  (
            .in0(_gnd_net_),
            .in1(N__21896),
            .in2(N__25055),
            .in3(N__21338),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .clk(N__47286),
            .ce(N__23673),
            .sr(N__46731));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_4_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_4_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_4_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_27_LC_4_16_3  (
            .in0(_gnd_net_),
            .in1(N__25955),
            .in2(N__21907),
            .in3(N__21323),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .clk(N__47286),
            .ce(N__23673),
            .sr(N__46731));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_4_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_4_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_4_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_28_LC_4_16_4  (
            .in0(_gnd_net_),
            .in1(N__21900),
            .in2(N__25906),
            .in3(N__21308),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .clk(N__47286),
            .ce(N__23673),
            .sr(N__46731));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_4_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_4_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_4_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_29_LC_4_16_5  (
            .in0(_gnd_net_),
            .in1(N__25848),
            .in2(N__21908),
            .in3(N__21293),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .clk(N__47286),
            .ce(N__23673),
            .sr(N__46731));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_4_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_4_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_4_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_30_LC_4_16_6  (
            .in0(_gnd_net_),
            .in1(N__21904),
            .in2(N__25791),
            .in3(N__21275),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ),
            .clk(N__47286),
            .ce(N__23673),
            .sr(N__46731));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_4_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_4_16_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_4_16_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_31_LC_4_16_7  (
            .in0(N__21905),
            .in1(N__25658),
            .in2(_gnd_net_),
            .in3(N__21272),
            .lcout(\current_shift_inst.PI_CTRL.un8_enablelto31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47286),
            .ce(N__23673),
            .sr(N__46731));
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_4_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_4_17_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_4_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_12_LC_4_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23956),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47279),
            .ce(N__23678),
            .sr(N__46736));
    defparam CONSTANT_ONE_LUT4_LC_4_30_6.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_4_30_6.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_4_30_6.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_4_30_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_7_LC_5_7_0.C_ON=1'b0;
    defparam counter_7_LC_5_7_0.SEQ_MODE=4'b1010;
    defparam counter_7_LC_5_7_0.LUT_INIT=16'b0010101010101010;
    LogicCell40 counter_7_LC_5_7_0 (
            .in0(N__21485),
            .in1(N__21713),
            .in2(N__21629),
            .in3(N__21655),
            .lcout(counterZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47345),
            .ce(),
            .sr(N__46671));
    defparam counter_RNI800G_7_LC_5_7_2.C_ON=1'b0;
    defparam counter_RNI800G_7_LC_5_7_2.SEQ_MODE=4'b0000;
    defparam counter_RNI800G_7_LC_5_7_2.LUT_INIT=16'b1100110000000000;
    LogicCell40 counter_RNI800G_7_LC_5_7_2 (
            .in0(_gnd_net_),
            .in1(N__21592),
            .in2(_gnd_net_),
            .in3(N__21478),
            .lcout(),
            .ltout(un2_counter_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNI3BSP_1_LC_5_7_3.C_ON=1'b0;
    defparam counter_RNI3BSP_1_LC_5_7_3.SEQ_MODE=4'b0000;
    defparam counter_RNI3BSP_1_LC_5_7_3.LUT_INIT=16'b0000000000010000;
    LogicCell40 counter_RNI3BSP_1_LC_5_7_3 (
            .in0(N__21465),
            .in1(N__21442),
            .in2(N__21431),
            .in3(N__21428),
            .lcout(un2_counter_9),
            .ltout(un2_counter_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_10khz_RNIIENA2_LC_5_7_4.C_ON=1'b0;
    defparam clk_10khz_RNIIENA2_LC_5_7_4.SEQ_MODE=4'b0000;
    defparam clk_10khz_RNIIENA2_LC_5_7_4.LUT_INIT=16'b0110101010101010;
    LogicCell40 clk_10khz_RNIIENA2_LC_5_7_4 (
            .in0(N__21869),
            .in1(N__21712),
            .in2(N__21404),
            .in3(N__21620),
            .lcout(clk_10khz_RNIIENAZ0Z2),
            .ltout(clk_10khz_RNIIENAZ0Z2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_cnv_0_LC_5_7_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_cnv_0_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.prop_term_cnv_0_LC_5_7_5 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_cnv_0_LC_5_7_5  (
            .in0(N__34537),
            .in1(_gnd_net_),
            .in2(N__21401),
            .in3(N__21870),
            .lcout(N_702_g),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_10khz_LC_5_7_7.C_ON=1'b0;
    defparam clk_10khz_LC_5_7_7.SEQ_MODE=4'b1010;
    defparam clk_10khz_LC_5_7_7.LUT_INIT=16'b0110110011001100;
    LogicCell40 clk_10khz_LC_5_7_7 (
            .in0(N__21621),
            .in1(N__21871),
            .in2(N__21665),
            .in3(N__21715),
            .lcout(clk_10khz_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47345),
            .ce(),
            .sr(N__46671));
    defparam \pwm_generator_inst.threshold_2_LC_5_8_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_2_LC_5_8_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_2_LC_5_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_2_LC_5_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21398),
            .lcout(\pwm_generator_inst.thresholdZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47341),
            .ce(),
            .sr(N__46679));
    defparam counter_10_LC_5_8_7.C_ON=1'b0;
    defparam counter_10_LC_5_8_7.SEQ_MODE=4'b1010;
    defparam counter_10_LC_5_8_7.LUT_INIT=16'b0100110011001100;
    LogicCell40 counter_10_LC_5_8_7 (
            .in0(N__21719),
            .in1(N__21680),
            .in2(N__21666),
            .in3(N__21628),
            .lcout(counterZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47341),
            .ce(),
            .sr(N__46679));
    defparam \pwm_generator_inst.threshold_8_LC_5_10_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_8_LC_5_10_5 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_8_LC_5_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_8_LC_5_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21581),
            .lcout(\pwm_generator_inst.thresholdZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47331),
            .ce(),
            .sr(N__46696));
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_5_11_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_5_11_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_5_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_1_LC_5_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23864),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47323),
            .ce(N__23585),
            .sr(N__46705));
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_5_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_5_12_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_5_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_11_LC_5_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24032),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47316),
            .ce(N__23635),
            .sr(N__46709));
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_5_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_5_12_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_5_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_9_LC_5_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24170),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47316),
            .ce(N__23635),
            .sr(N__46709));
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_5_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_5_12_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_5_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_5_LC_5_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24443),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47316),
            .ce(N__23635),
            .sr(N__46709));
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_5_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_5_13_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_5_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_0_LC_5_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23911),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47304),
            .ce(N__23641),
            .sr(N__46713));
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_5_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_5_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_5_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_4_LC_5_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23461),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47304),
            .ce(N__23641),
            .sr(N__46713));
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_5_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_5_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_5_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_17_LC_5_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24659),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47304),
            .ce(N__23641),
            .sr(N__46713));
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_5_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_5_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_5_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_2_LC_5_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23806),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47304),
            .ce(N__23641),
            .sr(N__46713));
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_5_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_5_13_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_5_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_8_LC_5_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24236),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47304),
            .ce(N__23641),
            .sr(N__46713));
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_5_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_5_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_5_13_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_6_LC_5_13_5  (
            .in0(N__24364),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47304),
            .ce(N__23641),
            .sr(N__46713));
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_5_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_5_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_5_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_3_LC_5_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23734),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47304),
            .ce(N__23641),
            .sr(N__46713));
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_5_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_5_14_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_5_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_15_LC_5_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24797),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47295),
            .ce(N__23636),
            .sr(N__46721));
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_5_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_5_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_5_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_19_LC_5_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24515),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47295),
            .ce(N__23636),
            .sr(N__46721));
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_5_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_5_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_5_14_2 .LUT_INIT=16'b1110111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_11_LC_5_14_2  (
            .in0(N__22726),
            .in1(N__25678),
            .in2(N__22625),
            .in3(N__24002),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47295),
            .ce(N__23636),
            .sr(N__46721));
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_5_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_5_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_5_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_10_LC_5_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24100),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47295),
            .ce(N__23636),
            .sr(N__46721));
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_5_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_5_14_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_5_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_13_LC_5_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24946),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47295),
            .ce(N__23636),
            .sr(N__46721));
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_5_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_5_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_5_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_14_LC_5_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24911),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47295),
            .ce(N__23636),
            .sr(N__46721));
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_5_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_5_14_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_5_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_20_LC_5_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25442),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47295),
            .ce(N__23636),
            .sr(N__46721));
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_5_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_5_14_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_5_14_7 .LUT_INIT=16'b1010100011111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_10_LC_5_14_7  (
            .in0(N__24077),
            .in1(N__22725),
            .in2(N__25682),
            .in3(N__22619),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47295),
            .ce(N__23636),
            .sr(N__46721));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_5_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_5_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_5_15_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_5_15_0  (
            .in0(N__25907),
            .in1(N__25954),
            .in2(N__25787),
            .in3(N__23990),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_10_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA53P2_10_LC_5_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA53P2_10_LC_5_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA53P2_10_LC_5_15_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIA53P2_10_LC_5_15_1  (
            .in0(N__21818),
            .in1(N__21812),
            .in2(N__21821),
            .in3(N__21806),
            .lcout(\current_shift_inst.PI_CTRL.N_47_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_5_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_5_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_5_15_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_5_15_2  (
            .in0(N__25105),
            .in1(N__25180),
            .in2(N__25054),
            .in3(N__25396),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_11_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_5_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_5_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_5_15_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_5_15_3  (
            .in0(N__24875),
            .in1(N__24982),
            .in2(N__24755),
            .in3(N__24050),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_9_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_0_10_LC_5_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_0_10_LC_5_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_0_10_LC_5_15_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIB98M_0_10_LC_5_15_5  (
            .in0(N__25257),
            .in1(N__24825),
            .in2(N__25853),
            .in3(N__24119),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_8_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_5_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_5_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_5_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_16_LC_5_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24718),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47280),
            .ce(N__23675),
            .sr(N__46729));
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_5_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_5_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_5_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_21_LC_5_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25361),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47280),
            .ce(N__23675),
            .sr(N__46729));
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_5_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_5_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_5_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_18_LC_5_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24577),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47280),
            .ce(N__23675),
            .sr(N__46729));
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_5_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_5_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_5_16_3 .LUT_INIT=16'b1011101010110000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_30_LC_5_16_3  (
            .in0(N__25745),
            .in1(N__22614),
            .in2(N__25677),
            .in3(N__22741),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47280),
            .ce(N__23675),
            .sr(N__46729));
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_5_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_5_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_5_16_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_23_LC_5_16_4  (
            .in0(N__25222),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47280),
            .ce(N__23675),
            .sr(N__46729));
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_5_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_5_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_5_16_6 .LUT_INIT=16'b1110000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_4_LC_5_16_6  (
            .in0(N__22742),
            .in1(N__25654),
            .in2(N__23438),
            .in3(N__22615),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47280),
            .ce(N__23675),
            .sr(N__46729));
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_5_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_5_16_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_5_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_22_LC_5_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25288),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47280),
            .ce(N__23675),
            .sr(N__46729));
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_5_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_5_17_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_5_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_24_LC_5_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25144),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47267),
            .ce(N__23677),
            .sr(N__46732));
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_5_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_5_17_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_5_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_25_LC_5_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25730),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47267),
            .ce(N__23677),
            .sr(N__46732));
    defparam \current_shift_inst.phase_valid_RNISLOR2_LC_7_7_4 .C_ON=1'b0;
    defparam \current_shift_inst.phase_valid_RNISLOR2_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.phase_valid_RNISLOR2_LC_7_7_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \current_shift_inst.phase_valid_RNISLOR2_LC_7_7_4  (
            .in0(N__32393),
            .in1(N__21875),
            .in2(N__34536),
            .in3(N__21854),
            .lcout(\current_shift_inst.phase_valid_RNISLORZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_7_LC_7_8_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_7_LC_7_8_0 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_7_LC_7_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_7_LC_7_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21845),
            .lcout(\pwm_generator_inst.thresholdZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47332),
            .ce(),
            .sr(N__46660));
    defparam \pwm_generator_inst.threshold_1_LC_7_8_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_1_LC_7_8_4 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_1_LC_7_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_1_LC_7_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21977),
            .lcout(\pwm_generator_inst.thresholdZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47332),
            .ce(),
            .sr(N__46660));
    defparam \pwm_generator_inst.threshold_4_LC_7_9_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_4_LC_7_9_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_4_LC_7_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_4_LC_7_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21965),
            .lcout(\pwm_generator_inst.thresholdZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47324),
            .ce(),
            .sr(N__46672));
    defparam \pwm_generator_inst.threshold_9_LC_7_10_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_9_LC_7_10_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_9_LC_7_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_9_LC_7_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21956),
            .lcout(\pwm_generator_inst.thresholdZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47317),
            .ce(),
            .sr(N__46680));
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_7_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_7_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_7_11_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_8_LC_7_11_1  (
            .in0(N__44157),
            .in1(N__41768),
            .in2(_gnd_net_),
            .in3(N__43851),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47305),
            .ce(N__31226),
            .sr(N__46686));
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_7_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_7_12_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_7_12_0 .LUT_INIT=16'b1000101010001111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_5_LC_7_12_0  (
            .in0(N__24413),
            .in1(N__22604),
            .in2(N__25676),
            .in3(N__22739),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47296),
            .ce(N__23679),
            .sr(N__46697));
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_7_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_7_12_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_7_12_1 .LUT_INIT=16'b1111001100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_6_LC_7_12_1  (
            .in0(N__22740),
            .in1(N__25649),
            .in2(N__22624),
            .in3(N__24338),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47296),
            .ce(N__23679),
            .sr(N__46697));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_7_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_7_13_0 .LUT_INIT=16'b1111111100001101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_7_13_0  (
            .in0(N__23710),
            .in1(N__22406),
            .in2(N__23498),
            .in3(N__22049),
            .lcout(\current_shift_inst.PI_CTRL.N_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_7_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_7_13_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_7_13_1  (
            .in0(N__24190),
            .in1(N__24290),
            .in2(N__24465),
            .in3(N__24386),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_7_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_7_13_2 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_7_13_2  (
            .in0(N__23709),
            .in1(N__23493),
            .in2(N__21941),
            .in3(N__24255),
            .lcout(\current_shift_inst.PI_CTRL.N_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB4HQ_8_LC_7_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB4HQ_8_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB4HQ_8_LC_7_13_4 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIB4HQ_8_LC_7_13_4  (
            .in0(_gnd_net_),
            .in1(N__24189),
            .in2(_gnd_net_),
            .in3(N__24254),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_5_LC_7_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_5_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_5_LC_7_13_5 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI4JA22_5_LC_7_13_5  (
            .in0(N__24459),
            .in1(N__24291),
            .in2(N__22052),
            .in3(N__24387),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIOU8U3_18_LC_7_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIOU8U3_18_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIOU8U3_18_LC_7_13_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIOU8U3_18_LC_7_13_6  (
            .in0(N__24610),
            .in1(N__22447),
            .in2(N__25675),
            .in3(N__21988),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIE7HME_18_LC_7_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIE7HME_18_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIE7HME_18_LC_7_13_7 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIE7HME_18_LC_7_13_7  (
            .in0(N__21998),
            .in1(N__22018),
            .in2(N__22043),
            .in3(N__22040),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNITMGQ3_18_LC_7_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNITMGQ3_18_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNITMGQ3_18_LC_7_14_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNITMGQ3_18_LC_7_14_1  (
            .in0(N__24611),
            .in1(N__25632),
            .in2(N__22465),
            .in3(N__22033),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_7_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_7_14_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_7_14_2  (
            .in0(N__24880),
            .in1(N__24972),
            .in2(N__24753),
            .in3(N__24063),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIBHHP7_18_LC_7_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIBHHP7_18_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIBHHP7_18_LC_7_14_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIBHHP7_18_LC_7_14_4  (
            .in0(N__22034),
            .in1(N__24612),
            .in2(N__22466),
            .in3(N__22019),
            .lcout(\current_shift_inst.PI_CTRL.N_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_7_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_7_14_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_7_14_5  (
            .in0(N__25250),
            .in1(N__24821),
            .in2(N__25852),
            .in3(N__24127),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA53P2_0_10_LC_7_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA53P2_0_10_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA53P2_0_10_LC_7_14_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIA53P2_0_10_LC_7_14_6  (
            .in0(N__22073),
            .in1(N__22082),
            .in2(N__22007),
            .in3(N__22004),
            .lcout(\current_shift_inst.PI_CTRL.N_46_21 ),
            .ltout(\current_shift_inst.PI_CTRL.N_46_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1IOH6_18_LC_7_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1IOH6_18_LC_7_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1IOH6_18_LC_7_14_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI1IOH6_18_LC_7_14_7  (
            .in0(N__24613),
            .in1(N__22448),
            .in2(N__21992),
            .in3(N__21989),
            .lcout(\current_shift_inst.PI_CTRL.N_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_7_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_7_15_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_7_15_2  (
            .in0(N__25886),
            .in1(N__25946),
            .in2(N__25795),
            .in3(N__23981),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_7_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_7_15_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_7_15_3  (
            .in0(N__25091),
            .in1(N__25166),
            .in2(N__25040),
            .in3(N__25385),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_7_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_7_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_7_15_4 .LUT_INIT=16'b1101110011010000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_15_LC_7_15_4  (
            .in0(N__22551),
            .in1(N__24770),
            .in2(N__25667),
            .in3(N__22689),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47268),
            .ce(N__23683),
            .sr(N__46714));
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_7_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_7_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_7_15_5 .LUT_INIT=16'b1110000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_23_LC_7_15_5  (
            .in0(N__22690),
            .in1(N__25614),
            .in2(N__25202),
            .in3(N__22552),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47268),
            .ce(N__23683),
            .sr(N__46714));
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_7_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_7_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_7_16_0 .LUT_INIT=16'b1011101010110000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_27_LC_7_16_0  (
            .in0(N__25922),
            .in1(N__22591),
            .in2(N__25666),
            .in3(N__22735),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47259),
            .ce(N__23671),
            .sr(N__46722));
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_7_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_7_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_7_16_1 .LUT_INIT=16'b1100111110001000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_28_LC_7_16_1  (
            .in0(N__22736),
            .in1(N__25865),
            .in2(N__22621),
            .in3(N__25613),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47259),
            .ce(N__23671),
            .sr(N__46722));
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_7_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_7_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_7_16_2 .LUT_INIT=16'b1011101010110000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_26_LC_7_16_2  (
            .in0(N__25007),
            .in1(N__22590),
            .in2(N__25665),
            .in3(N__22734),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47259),
            .ce(N__23671),
            .sr(N__46722));
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_7_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_7_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_7_16_3 .LUT_INIT=16'b1110111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_31_LC_7_16_3  (
            .in0(N__22738),
            .in1(N__25603),
            .in2(N__22623),
            .in3(N__25490),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47259),
            .ce(N__23671),
            .sr(N__46722));
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_7_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_7_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_7_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_7_LC_7_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24316),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47259),
            .ce(N__23671),
            .sr(N__46722));
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_7_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_7_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_7_16_5 .LUT_INIT=16'b1110111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_29_LC_7_16_5  (
            .in0(N__22737),
            .in1(N__25602),
            .in2(N__22622),
            .in3(N__25808),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47259),
            .ce(N__23671),
            .sr(N__46722));
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_7_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_7_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_7_16_6 .LUT_INIT=16'b1011101010110000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_24_LC_7_16_6  (
            .in0(N__25118),
            .in1(N__22589),
            .in2(N__25664),
            .in3(N__22732),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47259),
            .ce(N__23671),
            .sr(N__46722));
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_7_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_7_16_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_7_16_7 .LUT_INIT=16'b1110111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_25_LC_7_16_7  (
            .in0(N__22733),
            .in1(N__25601),
            .in2(N__22620),
            .in3(N__25070),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47259),
            .ce(N__23671),
            .sr(N__46722));
    defparam \current_shift_inst.control_input_0_LC_7_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_0_LC_7_17_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_0_LC_7_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_0_LC_7_17_0  (
            .in0(_gnd_net_),
            .in1(N__22751),
            .in2(N__31417),
            .in3(N__31418),
            .lcout(\current_shift_inst.control_inputZ0Z_0 ),
            .ltout(),
            .carryin(bfn_7_17_0_),
            .carryout(\current_shift_inst.control_input_1_cry_0 ),
            .clk(N__47251),
            .ce(N__23027),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_1_LC_7_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_1_LC_7_17_1 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_1_LC_7_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_1_LC_7_17_1  (
            .in0(_gnd_net_),
            .in1(N__22871),
            .in2(_gnd_net_),
            .in3(N__22100),
            .lcout(\current_shift_inst.control_inputZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_0 ),
            .carryout(\current_shift_inst.control_input_1_cry_1 ),
            .clk(N__47251),
            .ce(N__23027),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_2_LC_7_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_2_LC_7_17_2 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_2_LC_7_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_2_LC_7_17_2  (
            .in0(_gnd_net_),
            .in1(N__22862),
            .in2(_gnd_net_),
            .in3(N__22097),
            .lcout(\current_shift_inst.control_inputZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_1 ),
            .carryout(\current_shift_inst.control_input_1_cry_2 ),
            .clk(N__47251),
            .ce(N__23027),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_3_LC_7_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_3_LC_7_17_3 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_3_LC_7_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_3_LC_7_17_3  (
            .in0(_gnd_net_),
            .in1(N__22853),
            .in2(_gnd_net_),
            .in3(N__22094),
            .lcout(\current_shift_inst.control_inputZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_2 ),
            .carryout(\current_shift_inst.control_input_1_cry_3 ),
            .clk(N__47251),
            .ce(N__23027),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_4_LC_7_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_4_LC_7_17_4 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_4_LC_7_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_4_LC_7_17_4  (
            .in0(_gnd_net_),
            .in1(N__22844),
            .in2(_gnd_net_),
            .in3(N__22091),
            .lcout(\current_shift_inst.control_inputZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_3 ),
            .carryout(\current_shift_inst.control_input_1_cry_4 ),
            .clk(N__47251),
            .ce(N__23027),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_5_LC_7_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_5_LC_7_17_5 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_5_LC_7_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_5_LC_7_17_5  (
            .in0(_gnd_net_),
            .in1(N__22835),
            .in2(_gnd_net_),
            .in3(N__22088),
            .lcout(\current_shift_inst.control_inputZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_4 ),
            .carryout(\current_shift_inst.control_input_1_cry_5 ),
            .clk(N__47251),
            .ce(N__23027),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_6_LC_7_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_6_LC_7_17_6 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_6_LC_7_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_6_LC_7_17_6  (
            .in0(_gnd_net_),
            .in1(N__22826),
            .in2(_gnd_net_),
            .in3(N__22085),
            .lcout(\current_shift_inst.control_inputZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_5 ),
            .carryout(\current_shift_inst.control_input_1_cry_6 ),
            .clk(N__47251),
            .ce(N__23027),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_7_LC_7_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_7_LC_7_17_7 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_7_LC_7_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_7_LC_7_17_7  (
            .in0(_gnd_net_),
            .in1(N__22817),
            .in2(_gnd_net_),
            .in3(N__22127),
            .lcout(\current_shift_inst.control_inputZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_6 ),
            .carryout(\current_shift_inst.control_input_1_cry_7 ),
            .clk(N__47251),
            .ce(N__23027),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_8_LC_7_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_8_LC_7_18_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_8_LC_7_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_8_LC_7_18_0  (
            .in0(_gnd_net_),
            .in1(N__22796),
            .in2(_gnd_net_),
            .in3(N__22124),
            .lcout(\current_shift_inst.control_inputZ0Z_8 ),
            .ltout(),
            .carryin(bfn_7_18_0_),
            .carryout(\current_shift_inst.control_input_1_cry_8 ),
            .clk(N__47243),
            .ce(N__23026),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_9_LC_7_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_9_LC_7_18_1 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_9_LC_7_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_9_LC_7_18_1  (
            .in0(_gnd_net_),
            .in1(N__22988),
            .in2(_gnd_net_),
            .in3(N__22121),
            .lcout(\current_shift_inst.control_inputZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_8 ),
            .carryout(\current_shift_inst.control_input_1_cry_9 ),
            .clk(N__47243),
            .ce(N__23026),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_10_LC_7_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_10_LC_7_18_2 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_10_LC_7_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_10_LC_7_18_2  (
            .in0(_gnd_net_),
            .in1(N__22979),
            .in2(_gnd_net_),
            .in3(N__22118),
            .lcout(\current_shift_inst.control_inputZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_9 ),
            .carryout(\current_shift_inst.control_input_1_cry_10 ),
            .clk(N__47243),
            .ce(N__23026),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_11_LC_7_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_11_LC_7_18_3 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_11_LC_7_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_11_LC_7_18_3  (
            .in0(_gnd_net_),
            .in1(N__22970),
            .in2(_gnd_net_),
            .in3(N__22115),
            .lcout(\current_shift_inst.control_inputZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_10 ),
            .carryout(\current_shift_inst.control_input_1_cry_11 ),
            .clk(N__47243),
            .ce(N__23026),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_12_LC_7_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_12_LC_7_18_4 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_12_LC_7_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_12_LC_7_18_4  (
            .in0(_gnd_net_),
            .in1(N__22949),
            .in2(_gnd_net_),
            .in3(N__22112),
            .lcout(\current_shift_inst.control_inputZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_11 ),
            .carryout(\current_shift_inst.control_input_1_cry_12 ),
            .clk(N__47243),
            .ce(N__23026),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_13_LC_7_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_13_LC_7_18_5 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_13_LC_7_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_13_LC_7_18_5  (
            .in0(_gnd_net_),
            .in1(N__22928),
            .in2(_gnd_net_),
            .in3(N__22109),
            .lcout(\current_shift_inst.control_inputZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_12 ),
            .carryout(\current_shift_inst.control_input_1_cry_13 ),
            .clk(N__47243),
            .ce(N__23026),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_14_LC_7_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_14_LC_7_18_6 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_14_LC_7_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_14_LC_7_18_6  (
            .in0(_gnd_net_),
            .in1(N__22907),
            .in2(_gnd_net_),
            .in3(N__22106),
            .lcout(\current_shift_inst.control_inputZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_13 ),
            .carryout(\current_shift_inst.control_input_1_cry_14 ),
            .clk(N__47243),
            .ce(N__23026),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_15_LC_7_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_15_LC_7_18_7 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_15_LC_7_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_15_LC_7_18_7  (
            .in0(_gnd_net_),
            .in1(N__22898),
            .in2(_gnd_net_),
            .in3(N__22103),
            .lcout(\current_shift_inst.control_inputZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_14 ),
            .carryout(\current_shift_inst.control_input_1_cry_15 ),
            .clk(N__47243),
            .ce(N__23026),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_16_LC_7_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_16_LC_7_19_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_16_LC_7_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_16_LC_7_19_0  (
            .in0(_gnd_net_),
            .in1(N__22889),
            .in2(_gnd_net_),
            .in3(N__22154),
            .lcout(\current_shift_inst.control_inputZ0Z_16 ),
            .ltout(),
            .carryin(bfn_7_19_0_),
            .carryout(\current_shift_inst.control_input_1_cry_16 ),
            .clk(N__47235),
            .ce(N__23037),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_17_LC_7_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_17_LC_7_19_1 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_17_LC_7_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_17_LC_7_19_1  (
            .in0(_gnd_net_),
            .in1(N__22880),
            .in2(_gnd_net_),
            .in3(N__22151),
            .lcout(\current_shift_inst.control_inputZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_16 ),
            .carryout(\current_shift_inst.control_input_1_cry_17 ),
            .clk(N__47235),
            .ce(N__23037),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_18_LC_7_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_18_LC_7_19_2 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_18_LC_7_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_18_LC_7_19_2  (
            .in0(_gnd_net_),
            .in1(N__23117),
            .in2(_gnd_net_),
            .in3(N__22148),
            .lcout(\current_shift_inst.control_inputZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_17 ),
            .carryout(\current_shift_inst.control_input_1_cry_18 ),
            .clk(N__47235),
            .ce(N__23037),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_19_LC_7_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_19_LC_7_19_3 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_19_LC_7_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_19_LC_7_19_3  (
            .in0(_gnd_net_),
            .in1(N__23108),
            .in2(_gnd_net_),
            .in3(N__22145),
            .lcout(\current_shift_inst.control_inputZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_18 ),
            .carryout(\current_shift_inst.control_input_1_cry_19 ),
            .clk(N__47235),
            .ce(N__23037),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_20_LC_7_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_20_LC_7_19_4 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_20_LC_7_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_20_LC_7_19_4  (
            .in0(_gnd_net_),
            .in1(N__23099),
            .in2(_gnd_net_),
            .in3(N__22142),
            .lcout(\current_shift_inst.control_inputZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_19 ),
            .carryout(\current_shift_inst.control_input_1_cry_20 ),
            .clk(N__47235),
            .ce(N__23037),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_21_LC_7_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_21_LC_7_19_5 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_21_LC_7_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_21_LC_7_19_5  (
            .in0(_gnd_net_),
            .in1(N__23090),
            .in2(_gnd_net_),
            .in3(N__22139),
            .lcout(\current_shift_inst.control_inputZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_20 ),
            .carryout(\current_shift_inst.control_input_1_cry_21 ),
            .clk(N__47235),
            .ce(N__23037),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_22_LC_7_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_22_LC_7_19_6 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_22_LC_7_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_22_LC_7_19_6  (
            .in0(_gnd_net_),
            .in1(N__23081),
            .in2(_gnd_net_),
            .in3(N__22136),
            .lcout(\current_shift_inst.control_inputZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_21 ),
            .carryout(\current_shift_inst.control_input_1_cry_22 ),
            .clk(N__47235),
            .ce(N__23037),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_23_LC_7_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_23_LC_7_19_7 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_23_LC_7_19_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_23_LC_7_19_7  (
            .in0(_gnd_net_),
            .in1(N__23072),
            .in2(_gnd_net_),
            .in3(N__22133),
            .lcout(\current_shift_inst.control_inputZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_22 ),
            .carryout(\current_shift_inst.control_input_1_cry_23 ),
            .clk(N__47235),
            .ce(N__23037),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_24_LC_7_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_24_LC_7_20_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_24_LC_7_20_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_24_LC_7_20_0  (
            .in0(_gnd_net_),
            .in1(N__23063),
            .in2(_gnd_net_),
            .in3(N__22130),
            .lcout(\current_shift_inst.control_inputZ0Z_24 ),
            .ltout(),
            .carryin(bfn_7_20_0_),
            .carryout(\current_shift_inst.control_input_1_cry_24 ),
            .clk(N__47228),
            .ce(N__23038),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_1_cry_24_THRU_LUT4_0_LC_7_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_1_cry_24_THRU_LUT4_0_LC_7_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_1_cry_24_THRU_LUT4_0_LC_7_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.control_input_1_cry_24_THRU_LUT4_0_LC_7_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22226),
            .lcout(\current_shift_inst.control_input_1_cry_24_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MIN_D1_LC_8_5_4.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MIN_D1_LC_8_5_4.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MIN_D1_LC_8_5_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_PH2_MIN_D1_LC_8_5_4 (
            .in0(N__22223),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_min_comp2_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47342),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MAX_D1_LC_8_6_5.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MAX_D1_LC_8_6_5.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MAX_D1_LC_8_6_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_PH2_MAX_D1_LC_8_6_5 (
            .in0(N__22211),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_max_comp2_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47337),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_0_LC_8_8_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_0_LC_8_8_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_0_LC_8_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_0_LC_8_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22196),
            .lcout(\pwm_generator_inst.thresholdZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47325),
            .ce(),
            .sr(N__46651));
    defparam \pwm_generator_inst.threshold_6_LC_8_9_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_6_LC_8_9_0 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_6_LC_8_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_6_LC_8_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22184),
            .lcout(\pwm_generator_inst.thresholdZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47318),
            .ce(),
            .sr(N__46661));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_8_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_8_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_8_9_5 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_8_9_5  (
            .in0(N__39678),
            .in1(N__39846),
            .in2(N__40006),
            .in3(N__28928),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47318),
            .ce(),
            .sr(N__46661));
    defparam \pwm_generator_inst.threshold_3_LC_8_9_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_3_LC_8_9_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_3_LC_8_9_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \pwm_generator_inst.threshold_3_LC_8_9_6  (
            .in0(N__22172),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.thresholdZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47318),
            .ce(),
            .sr(N__46661));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_8_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_8_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_8_9_7 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_8_9_7  (
            .in0(N__39679),
            .in1(N__39847),
            .in2(N__40007),
            .in3(N__29237),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47318),
            .ce(),
            .sr(N__46661));
    defparam \pwm_generator_inst.threshold_5_LC_8_10_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_5_LC_8_10_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_5_LC_8_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_5_LC_8_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22163),
            .lcout(\pwm_generator_inst.thresholdZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47306),
            .ce(),
            .sr(N__46673));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_8_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_8_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_8_10_5 .LUT_INIT=16'b1010101010000010;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_8_10_5  (
            .in0(N__23921),
            .in1(N__39654),
            .in2(N__40018),
            .in3(N__39845),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47306),
            .ce(),
            .sr(N__46673));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_8_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_8_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_8_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23381),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_11_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_8_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_8_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_8_11_1  (
            .in0(_gnd_net_),
            .in1(N__22322),
            .in2(N__22340),
            .in3(N__28377),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_8_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_8_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_8_11_2  (
            .in0(_gnd_net_),
            .in1(N__22298),
            .in2(N__22316),
            .in3(N__28354),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_8_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_8_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_8_11_3  (
            .in0(_gnd_net_),
            .in1(N__22274),
            .in2(N__22292),
            .in3(N__28312),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_8_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_8_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_8_11_4  (
            .in0(_gnd_net_),
            .in1(N__22268),
            .in2(N__23420),
            .in3(N__28279),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_8_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_8_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_8_11_5  (
            .in0(_gnd_net_),
            .in1(N__22262),
            .in2(N__23372),
            .in3(N__29074),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_8_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_8_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_8_11_6  (
            .in0(_gnd_net_),
            .in1(N__22238),
            .in2(N__22256),
            .in3(N__29041),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_8_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_8_11_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_8_11_7  (
            .in0(N__29008),
            .in1(N__22232),
            .in2(N__23930),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_8_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_8_12_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_8_12_0  (
            .in0(N__28978),
            .in1(N__22388),
            .in2(N__22400),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(bfn_8_12_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_8_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_8_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_8_12_1  (
            .in0(_gnd_net_),
            .in1(N__22382),
            .in2(N__27410),
            .in3(N__31142),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_8_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_8_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_8_12_2  (
            .in0(_gnd_net_),
            .in1(N__22376),
            .in2(N__23363),
            .in3(N__28945),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_8_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_8_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_8_12_3  (
            .in0(_gnd_net_),
            .in1(N__22370),
            .in2(N__27422),
            .in3(N__28916),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_8_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_8_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_8_12_4  (
            .in0(_gnd_net_),
            .in1(N__22364),
            .in2(N__23396),
            .in3(N__28886),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_8_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_8_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_8_12_5  (
            .in0(_gnd_net_),
            .in1(N__22358),
            .in2(N__23408),
            .in3(N__29282),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_8_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_8_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_8_12_6  (
            .in0(_gnd_net_),
            .in1(N__22352),
            .in2(N__27437),
            .in3(N__29254),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_8_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_8_12_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_8_12_7  (
            .in0(N__29225),
            .in1(N__22346),
            .in2(N__29354),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_8_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_8_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_8_13_0  (
            .in0(_gnd_net_),
            .in1(N__22433),
            .in2(N__31268),
            .in3(N__29198),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_16 ),
            .ltout(),
            .carryin(bfn_8_13_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_8_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_8_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_8_13_1  (
            .in0(_gnd_net_),
            .in1(N__22427),
            .in2(N__31256),
            .in3(N__29171),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_17 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_8_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_8_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_8_13_2  (
            .in0(_gnd_net_),
            .in1(N__22421),
            .in2(N__29342),
            .in3(N__29144),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_8_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_8_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_8_13_3  (
            .in0(_gnd_net_),
            .in1(N__22415),
            .in2(N__31244),
            .in3(N__29117),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_8_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_8_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_8_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22409),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_8_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_8_13_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_8_13_6  (
            .in0(N__23880),
            .in1(N__23778),
            .in2(_gnd_net_),
            .in3(N__23830),
            .lcout(\current_shift_inst.PI_CTRL.un1_enablelt3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_8_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_8_13_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_8_13_7  (
            .in0(N__39769),
            .in1(N__39962),
            .in2(_gnd_net_),
            .in3(N__39610),
            .lcout(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_8_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_8_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_8_14_1 .LUT_INIT=16'b1110111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_18_LC_8_14_1  (
            .in0(N__22684),
            .in1(N__25634),
            .in2(N__22609),
            .in3(N__24551),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47269),
            .ce(N__23631),
            .sr(N__46706));
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_8_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_8_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_8_14_2 .LUT_INIT=16'b1000101010001111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_9_LC_8_14_2  (
            .in0(N__24140),
            .in1(N__22555),
            .in2(N__25674),
            .in3(N__22688),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47269),
            .ce(N__23631),
            .sr(N__46706));
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_8_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_8_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_8_14_3 .LUT_INIT=16'b1100000011011101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_7_LC_8_14_3  (
            .in0(N__22686),
            .in1(N__24272),
            .in2(N__22611),
            .in3(N__25645),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47269),
            .ce(N__23631),
            .sr(N__46706));
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_8_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_8_14_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_8_14_4 .LUT_INIT=16'b1000101010001111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_8_LC_8_14_4  (
            .in0(N__24206),
            .in1(N__22554),
            .in2(N__25673),
            .in3(N__22687),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47269),
            .ce(N__23631),
            .sr(N__46706));
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_8_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_8_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_8_14_5 .LUT_INIT=16'b1110111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_21_LC_8_14_5  (
            .in0(N__22685),
            .in1(N__25635),
            .in2(N__22610),
            .in3(N__25331),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47269),
            .ce(N__23631),
            .sr(N__46706));
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_8_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_8_14_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_8_14_6 .LUT_INIT=16'b1011101010110000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_12_LC_8_14_6  (
            .in0(N__24992),
            .in1(N__22553),
            .in2(N__25672),
            .in3(N__22682),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47269),
            .ce(N__23631),
            .sr(N__46706));
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_8_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_8_14_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_8_14_7 .LUT_INIT=16'b1110111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_13_LC_8_14_7  (
            .in0(N__22683),
            .in1(N__25633),
            .in2(N__22608),
            .in3(N__24923),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47269),
            .ce(N__23631),
            .sr(N__46706));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_8_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_8_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_8_15_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_8_15_0  (
            .in0(N__25460),
            .in1(N__24533),
            .in2(N__25320),
            .in3(N__24677),
            .lcout(\current_shift_inst.PI_CTRL.N_47_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_8_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_8_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_8_15_1 .LUT_INIT=16'b1100100011111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_17_LC_8_15_1  (
            .in0(N__22721),
            .in1(N__24629),
            .in2(N__25669),
            .in3(N__22575),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47260),
            .ce(N__23684),
            .sr(N__46710));
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_8_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_8_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_8_15_2 .LUT_INIT=16'b1010111010001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_19_LC_8_15_2  (
            .in0(N__24485),
            .in1(N__25619),
            .in2(N__22613),
            .in3(N__22722),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47260),
            .ce(N__23684),
            .sr(N__46710));
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_8_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_8_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_8_15_3 .LUT_INIT=16'b1100100011111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_20_LC_8_15_3  (
            .in0(N__22723),
            .in1(N__25412),
            .in2(N__25670),
            .in3(N__22576),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47260),
            .ce(N__23684),
            .sr(N__46710));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_8_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_8_15_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_8_15_4  (
            .in0(N__25461),
            .in1(N__24534),
            .in2(N__25321),
            .in3(N__24678),
            .lcout(\current_shift_inst.PI_CTRL.N_46_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_8_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_8_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_8_15_5 .LUT_INIT=16'b1100100011111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_22_LC_8_15_5  (
            .in0(N__22724),
            .in1(N__25268),
            .in2(N__25671),
            .in3(N__22577),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47260),
            .ce(N__23684),
            .sr(N__46710));
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_8_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_8_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_8_15_6 .LUT_INIT=16'b1010111010001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_14_LC_8_15_6  (
            .in0(N__24845),
            .in1(N__25618),
            .in2(N__22612),
            .in3(N__22719),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47260),
            .ce(N__23684),
            .sr(N__46710));
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_8_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_8_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_8_15_7 .LUT_INIT=16'b1100100011111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_16_LC_8_15_7  (
            .in0(N__22720),
            .in1(N__24692),
            .in2(N__25668),
            .in3(N__22574),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47260),
            .ce(N__23684),
            .sr(N__46710));
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNO_0_LC_8_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNO_0_LC_8_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNO_0_LC_8_16_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_5_c_RNO_0_LC_8_16_0  (
            .in0(_gnd_net_),
            .in1(N__27487),
            .in2(_gnd_net_),
            .in3(N__29530),
            .lcout(\current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4H5J_19_LC_8_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4H5J_19_LC_8_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4H5J_19_LC_8_16_2 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4H5J_19_LC_8_16_2  (
            .in0(N__30417),
            .in1(N__30463),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI4H5J_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIH6661_17_LC_8_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIH6661_17_LC_8_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIH6661_17_LC_8_16_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIH6661_17_LC_8_16_3  (
            .in0(N__28001),
            .in1(N__29640),
            .in2(N__29684),
            .in3(N__27949),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIH6661_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR0UI_13_LC_8_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR0UI_13_LC_8_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR0UI_13_LC_8_16_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR0UI_13_LC_8_16_4  (
            .in0(_gnd_net_),
            .in1(N__29968),
            .in2(_gnd_net_),
            .in3(N__29929),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIR0UI_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQKU1_5_LC_8_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQKU1_5_LC_8_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQKU1_5_LC_8_16_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQKU1_5_LC_8_16_5  (
            .in0(N__29488),
            .in1(N__27803),
            .in2(N__27857),
            .in3(N__29453),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIVQKU1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNO_LC_8_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNO_LC_8_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNO_LC_8_16_6 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_5_c_RNO_LC_8_16_6  (
            .in0(N__27852),
            .in1(N__27488),
            .in2(N__29534),
            .in3(N__29487),
            .lcout(\current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAL3J_18_LC_8_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAL3J_18_LC_8_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAL3J_18_LC_8_16_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAL3J_18_LC_8_16_7  (
            .in0(_gnd_net_),
            .in1(N__27948),
            .in2(_gnd_net_),
            .in3(N__29641),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIAL3J_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CRY_0_LC_8_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CRY_0_LC_8_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CRY_0_LC_8_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CRY_0_LC_8_17_0  (
            .in0(_gnd_net_),
            .in1(N__30599),
            .in2(N__30605),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_17_0_),
            .carryout(\current_shift_inst.un38_control_input_0_cry_0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_0_c_inv_LC_8_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_0_c_inv_LC_8_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_0_c_inv_LC_8_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_0_c_inv_LC_8_17_1  (
            .in0(_gnd_net_),
            .in1(N__22787),
            .in2(N__29306),
            .in3(N__31435),
            .lcout(\current_shift_inst.z_i_0_31 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_0_c_THRU_CO ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_1_c_LC_8_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_1_c_LC_8_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_1_c_LC_8_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_1_c_LC_8_17_2  (
            .in0(_gnd_net_),
            .in1(N__25481),
            .in2(N__29615),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_0 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_2_c_LC_8_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_2_c_LC_8_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_2_c_LC_8_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_2_c_LC_8_17_3  (
            .in0(_gnd_net_),
            .in1(N__29581),
            .in2(N__26033),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_1 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_3_c_inv_LC_8_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_3_c_inv_LC_8_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_3_c_inv_LC_8_17_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_3_c_inv_LC_8_17_4  (
            .in0(N__25475),
            .in1(N__29555),
            .in2(N__22781),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un38_control_input_0_cry_3_c_invZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_2 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_4_c_LC_8_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_4_c_LC_8_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_4_c_LC_8_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_4_c_LC_8_17_5  (
            .in0(_gnd_net_),
            .in1(N__26012),
            .in2(N__26024),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_3 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_LC_8_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_LC_8_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_LC_8_17_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_5_c_LC_8_17_6  (
            .in0(_gnd_net_),
            .in1(N__22772),
            .in2(N__22766),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_4 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNI7HN13_LC_8_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNI7HN13_LC_8_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_5_c_RNI7HN13_LC_8_17_7 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_5_c_RNI7HN13_LC_8_17_7  (
            .in0(_gnd_net_),
            .in1(N__22757),
            .in2(N__25991),
            .in3(N__22745),
            .lcout(\current_shift_inst.control_input_1_axb_0 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_5 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_6_c_RNIHVR13_LC_8_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_6_c_RNIHVR13_LC_8_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_6_c_RNIHVR13_LC_8_18_0 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_6_c_RNIHVR13_LC_8_18_0  (
            .in0(_gnd_net_),
            .in1(N__26090),
            .in2(N__25967),
            .in3(N__22865),
            .lcout(\current_shift_inst.control_input_1_axb_1 ),
            .ltout(),
            .carryin(bfn_8_18_0_),
            .carryout(\current_shift_inst.un38_control_input_0_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_7_c_RNIRD023_LC_8_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_7_c_RNIRD023_LC_8_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_7_c_RNIRD023_LC_8_18_1 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_7_c_RNIRD023_LC_8_18_1  (
            .in0(_gnd_net_),
            .in1(N__26051),
            .in2(N__26006),
            .in3(N__22856),
            .lcout(\current_shift_inst.control_input_1_axb_2 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_7 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_8_c_RNIC9753_LC_8_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_8_c_RNIC9753_LC_8_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_8_c_RNIC9753_LC_8_18_2 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_8_c_RNIC9753_LC_8_18_2  (
            .in0(_gnd_net_),
            .in1(N__30002),
            .in2(N__29807),
            .in3(N__22847),
            .lcout(\current_shift_inst.control_input_1_axb_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_8 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_9_c_RNII9PR2_LC_8_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_9_c_RNII9PR2_LC_8_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_9_c_RNII9PR2_LC_8_18_3 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_9_c_RNII9PR2_LC_8_18_3  (
            .in0(_gnd_net_),
            .in1(N__26045),
            .in2(N__25982),
            .in3(N__22838),
            .lcout(\current_shift_inst.control_input_1_axb_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_9 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_10_c_RNIV96V1_LC_8_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_10_c_RNIV96V1_LC_8_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_10_c_RNIV96V1_LC_8_18_4 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_10_c_RNIV96V1_LC_8_18_4  (
            .in0(_gnd_net_),
            .in1(N__26096),
            .in2(N__26078),
            .in3(N__22829),
            .lcout(\current_shift_inst.control_input_1_axb_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_10 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_11_c_RNI9OAV1_LC_8_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_11_c_RNI9OAV1_LC_8_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_11_c_RNI9OAV1_LC_8_18_5 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_11_c_RNI9OAV1_LC_8_18_5  (
            .in0(_gnd_net_),
            .in1(N__30647),
            .in2(N__29993),
            .in3(N__22820),
            .lcout(\current_shift_inst.control_input_1_axb_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_11 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_12_c_RNIJ6FV1_LC_8_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_12_c_RNIJ6FV1_LC_8_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_12_c_RNIJ6FV1_LC_8_18_6 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_12_c_RNIJ6FV1_LC_8_18_6  (
            .in0(_gnd_net_),
            .in1(N__29891),
            .in2(N__29981),
            .in3(N__22811),
            .lcout(\current_shift_inst.control_input_1_axb_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_12 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_13_c_RNITKJV1_LC_8_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_13_c_RNITKJV1_LC_8_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_13_c_RNITKJV1_LC_8_18_7 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_13_c_RNITKJV1_LC_8_18_7  (
            .in0(_gnd_net_),
            .in1(N__25997),
            .in2(N__22808),
            .in3(N__22790),
            .lcout(\current_shift_inst.control_input_1_axb_8 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_13 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_14_c_RNI73OV1_LC_8_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_14_c_RNI73OV1_LC_8_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_14_c_RNI73OV1_LC_8_19_0 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_14_c_RNI73OV1_LC_8_19_0  (
            .in0(_gnd_net_),
            .in1(N__30137),
            .in2(N__26066),
            .in3(N__22982),
            .lcout(\current_shift_inst.control_input_1_axb_9 ),
            .ltout(),
            .carryin(bfn_8_19_0_),
            .carryout(\current_shift_inst.un38_control_input_0_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_15_c_RNIHHSV1_LC_8_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_15_c_RNIHHSV1_LC_8_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_15_c_RNIHHSV1_LC_8_19_1 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_15_c_RNIHHSV1_LC_8_19_1  (
            .in0(_gnd_net_),
            .in1(N__30287),
            .in2(N__30374),
            .in3(N__22973),
            .lcout(\current_shift_inst.control_input_1_axb_10 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_15 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_16_c_RNIRV002_LC_8_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_16_c_RNIRV002_LC_8_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_16_c_RNIRV002_LC_8_19_2 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_16_c_RNIRV002_LC_8_19_2  (
            .in0(_gnd_net_),
            .in1(N__26057),
            .in2(N__26117),
            .in3(N__22964),
            .lcout(\current_shift_inst.control_input_1_axb_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_16 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_17_c_RNI5E502_LC_8_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_17_c_RNI5E502_LC_8_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_17_c_RNI5E502_LC_8_19_3 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_17_c_RNI5E502_LC_8_19_3  (
            .in0(_gnd_net_),
            .in1(N__26084),
            .in2(N__22961),
            .in3(N__22943),
            .lcout(\current_shift_inst.control_input_1_axb_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_17 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_18_c_RNI6KA02_LC_8_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_18_c_RNI6KA02_LC_8_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_18_c_RNI6KA02_LC_8_19_4 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_18_c_RNI6KA02_LC_8_19_4  (
            .in0(_gnd_net_),
            .in1(N__25973),
            .in2(N__22940),
            .in3(N__22922),
            .lcout(\current_shift_inst.control_input_1_axb_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_18 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_19_c_RNICO912_LC_8_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_19_c_RNICO912_LC_8_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_19_c_RNICO912_LC_8_19_5 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_19_c_RNICO912_LC_8_19_5  (
            .in0(_gnd_net_),
            .in1(N__30383),
            .in2(N__22919),
            .in3(N__22901),
            .lcout(\current_shift_inst.control_input_1_axb_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_19 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_20_c_RNI92P32_LC_8_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_20_c_RNI92P32_LC_8_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_20_c_RNI92P32_LC_8_19_6 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_20_c_RNI92P32_LC_8_19_6  (
            .in0(_gnd_net_),
            .in1(N__31085),
            .in2(N__31019),
            .in3(N__22892),
            .lcout(\current_shift_inst.control_input_1_axb_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_20 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_21_c_RNIJGT32_LC_8_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_21_c_RNIJGT32_LC_8_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_21_c_RNIJGT32_LC_8_19_7 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_21_c_RNIJGT32_LC_8_19_7  (
            .in0(_gnd_net_),
            .in1(N__26141),
            .in2(N__30938),
            .in3(N__22883),
            .lcout(\current_shift_inst.control_input_1_axb_16 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_21 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_22_c_RNITU142_LC_8_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_22_c_RNITU142_LC_8_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_22_c_RNITU142_LC_8_20_0 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_22_c_RNITU142_LC_8_20_0  (
            .in0(_gnd_net_),
            .in1(N__26147),
            .in2(N__26156),
            .in3(N__22874),
            .lcout(\current_shift_inst.control_input_1_axb_17 ),
            .ltout(),
            .carryin(bfn_8_20_0_),
            .carryout(\current_shift_inst.un38_control_input_0_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_23_c_RNI7D642_LC_8_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_23_c_RNI7D642_LC_8_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_23_c_RNI7D642_LC_8_20_1 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_23_c_RNI7D642_LC_8_20_1  (
            .in0(_gnd_net_),
            .in1(N__31481),
            .in2(N__30923),
            .in3(N__23111),
            .lcout(\current_shift_inst.control_input_1_axb_18 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_23 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_24_c_RNIHRA42_LC_8_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_24_c_RNIHRA42_LC_8_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_24_c_RNIHRA42_LC_8_20_2 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_24_c_RNIHRA42_LC_8_20_2  (
            .in0(_gnd_net_),
            .in1(N__30785),
            .in2(N__31886),
            .in3(N__23102),
            .lcout(\current_shift_inst.control_input_1_axb_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_24 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_25_c_RNIR9F42_LC_8_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_25_c_RNIR9F42_LC_8_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_25_c_RNIR9F42_LC_8_20_3 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_25_c_RNIR9F42_LC_8_20_3  (
            .in0(_gnd_net_),
            .in1(N__31796),
            .in2(N__31730),
            .in3(N__23093),
            .lcout(\current_shift_inst.control_input_1_axb_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_25 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_26_c_RNI5OJ42_LC_8_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_26_c_RNI5OJ42_LC_8_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_26_c_RNI5OJ42_LC_8_20_4 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_26_c_RNI5OJ42_LC_8_20_4  (
            .in0(_gnd_net_),
            .in1(N__26102),
            .in2(N__30911),
            .in3(N__23084),
            .lcout(\current_shift_inst.control_input_1_axb_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_26 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_27_c_RNIF6O42_LC_8_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_27_c_RNIF6O42_LC_8_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_27_c_RNIF6O42_LC_8_20_5 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_27_c_RNIF6O42_LC_8_20_5  (
            .in0(_gnd_net_),
            .in1(N__26039),
            .in2(N__26126),
            .in3(N__23075),
            .lcout(\current_shift_inst.control_input_1_axb_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_27 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_28_c_RNIGCT42_LC_8_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_28_c_RNIGCT42_LC_8_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_28_c_RNIGCT42_LC_8_20_6 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_28_c_RNIGCT42_LC_8_20_6  (
            .in0(_gnd_net_),
            .in1(N__26108),
            .in2(N__30800),
            .in3(N__23066),
            .lcout(\current_shift_inst.control_input_1_axb_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_28 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_29_c_RNIMGS52_LC_8_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_0_cry_29_c_RNIMGS52_LC_8_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_29_c_RNIMGS52_LC_8_20_7 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_29_c_RNIMGS52_LC_8_20_7  (
            .in0(_gnd_net_),
            .in1(N__26132),
            .in2(N__31654),
            .in3(N__23057),
            .lcout(\current_shift_inst.control_input_1_axb_24 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_0_cry_29 ),
            .carryout(\current_shift_inst.un38_control_input_0_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_25_LC_8_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_25_LC_8_21_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_25_LC_8_21_0 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \current_shift_inst.control_input_25_LC_8_21_0  (
            .in0(_gnd_net_),
            .in1(N__30476),
            .in2(N__23054),
            .in3(N__23045),
            .lcout(\current_shift_inst.control_inputZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47221),
            .ce(N__23042),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MIN_D2_LC_9_5_7.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MIN_D2_LC_9_5_7.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MIN_D2_LC_9_5_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MIN_D2_LC_9_5_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23246),
            .lcout(il_min_comp2_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47338),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MAX_D1_LC_9_6_4.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_9_6_4.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_9_6_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MAX_D1_LC_9_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23240),
            .lcout(il_max_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47333),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_9_8_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_9_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_9_8_0  (
            .in0(_gnd_net_),
            .in1(N__23216),
            .in2(N__23225),
            .in3(N__27196),
            .lcout(\pwm_generator_inst.counter_i_0 ),
            .ltout(),
            .carryin(bfn_9_8_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_9_8_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_9_8_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_9_8_1  (
            .in0(N__27174),
            .in1(N__23210),
            .in2(N__23201),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_0 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_9_8_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_9_8_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_9_8_2  (
            .in0(_gnd_net_),
            .in1(N__23180),
            .in2(N__23192),
            .in3(N__27154),
            .lcout(\pwm_generator_inst.counter_i_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_1 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_9_8_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_9_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(N__23174),
            .in2(N__23168),
            .in3(N__27132),
            .lcout(\pwm_generator_inst.counter_i_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_2 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_9_8_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_9_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_9_8_4  (
            .in0(_gnd_net_),
            .in1(N__23159),
            .in2(N__23147),
            .in3(N__27111),
            .lcout(\pwm_generator_inst.counter_i_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_3 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_9_8_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_9_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_9_8_5  (
            .in0(_gnd_net_),
            .in1(N__23123),
            .in2(N__23135),
            .in3(N__27090),
            .lcout(\pwm_generator_inst.counter_i_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_4 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_9_8_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_9_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_9_8_6  (
            .in0(_gnd_net_),
            .in1(N__23339),
            .in2(N__23351),
            .in3(N__27345),
            .lcout(\pwm_generator_inst.counter_i_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_5 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_9_8_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_9_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_9_8_7  (
            .in0(_gnd_net_),
            .in1(N__23333),
            .in2(N__23324),
            .in3(N__27324),
            .lcout(\pwm_generator_inst.counter_i_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_6 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_9_9_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_9_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_9_9_0  (
            .in0(_gnd_net_),
            .in1(N__23300),
            .in2(N__23315),
            .in3(N__27303),
            .lcout(\pwm_generator_inst.counter_i_8 ),
            .ltout(),
            .carryin(bfn_9_9_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_9_9_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_9_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(N__23279),
            .in2(N__23294),
            .in3(N__27228),
            .lcout(\pwm_generator_inst.counter_i_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_8 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.pwm_out_LC_9_9_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.pwm_out_LC_9_9_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.pwm_out_LC_9_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.pwm_out_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23273),
            .lcout(pwm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47307),
            .ce(),
            .sr(N__46652));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_9_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_9_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_9_10_0 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_9_10_0  (
            .in0(N__39823),
            .in1(N__39661),
            .in2(N__40017),
            .in3(N__29030),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47297),
            .ce(),
            .sr(N__46662));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_9_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_9_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_9_10_1 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_9_10_1  (
            .in0(N__39658),
            .in1(N__40002),
            .in2(N__39854),
            .in3(N__28964),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47297),
            .ce(),
            .sr(N__46662));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_9_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_9_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_9_10_2 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_9_10_2  (
            .in0(N__39822),
            .in1(N__39660),
            .in2(N__40016),
            .in3(N__29063),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47297),
            .ce(),
            .sr(N__46662));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_9_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_9_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_9_10_3 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_9_10_3  (
            .in0(N__39656),
            .in1(N__39994),
            .in2(N__39852),
            .in3(N__28268),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47297),
            .ce(),
            .sr(N__46662));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_9_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_9_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_9_10_5 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_9_10_5  (
            .in0(N__39657),
            .in1(N__40001),
            .in2(N__39853),
            .in3(N__28997),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47297),
            .ce(),
            .sr(N__46662));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_9_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_9_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_9_10_6 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_9_10_6  (
            .in0(N__39821),
            .in1(N__39659),
            .in2(N__40015),
            .in3(N__28301),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47297),
            .ce(),
            .sr(N__46662));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_9_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_9_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_9_10_7 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_9_10_7  (
            .in0(N__39655),
            .in1(N__39990),
            .in2(N__39851),
            .in3(N__28343),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47297),
            .ce(),
            .sr(N__46662));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_9_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_9_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_9_11_1 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_LC_9_11_1  (
            .in0(N__43848),
            .in1(N__35432),
            .in2(N__44186),
            .in3(N__40346),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47287),
            .ce(N__31227),
            .sr(N__46674));
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_9_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_9_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_9_11_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_13_LC_9_11_2  (
            .in0(N__44281),
            .in1(N__44144),
            .in2(_gnd_net_),
            .in3(N__43847),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47287),
            .ce(N__31227),
            .sr(N__46674));
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_9_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_9_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_9_11_3 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_12_LC_9_11_3  (
            .in0(N__43846),
            .in1(_gnd_net_),
            .in2(N__44185),
            .in3(N__39407),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47287),
            .ce(N__31227),
            .sr(N__46674));
    defparam \phase_controller_inst1.stoper_hc.target_time_0_LC_9_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_0_LC_9_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_0_LC_9_11_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_0_LC_9_11_4  (
            .in0(N__40345),
            .in1(N__43844),
            .in2(N__42260),
            .in3(N__44139),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47287),
            .ce(N__31227),
            .sr(N__46674));
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_9_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_9_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_9_11_5 .LUT_INIT=16'b0000100000001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_5_LC_9_11_5  (
            .in0(N__43849),
            .in1(N__43956),
            .in2(N__44187),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47287),
            .ce(N__31227),
            .sr(N__46674));
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_9_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_9_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_9_11_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_10_LC_9_11_6  (
            .in0(N__35678),
            .in1(N__44140),
            .in2(_gnd_net_),
            .in3(N__43845),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47287),
            .ce(N__31227),
            .sr(N__46674));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_9_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_9_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_9_11_7 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_LC_9_11_7  (
            .in0(N__43850),
            .in1(_gnd_net_),
            .in2(N__44188),
            .in3(N__41670),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47287),
            .ce(N__31227),
            .sr(N__46674));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_9_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_9_12_2 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_9_12_2  (
            .in0(N__40040),
            .in1(N__27393),
            .in2(_gnd_net_),
            .in3(N__28387),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_9_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_9_12_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_9_12_7  (
            .in0(_gnd_net_),
            .in1(N__27389),
            .in2(_gnd_net_),
            .in3(N__40039),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_9_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_9_13_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_9_13_0 .LUT_INIT=16'b0011110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_0_LC_9_13_0  (
            .in0(_gnd_net_),
            .in1(N__23881),
            .in2(N__23912),
            .in3(N__23755),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ),
            .ltout(),
            .carryin(bfn_9_13_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_0 ),
            .clk(N__47270),
            .ce(N__23674),
            .sr(N__46687));
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_9_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_9_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_9_13_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_LC_9_13_1  (
            .in0(N__23753),
            .in1(N__23829),
            .in2(N__23863),
            .in3(N__23810),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ),
            .clk(N__47270),
            .ce(N__23674),
            .sr(N__46687));
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_9_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_9_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_9_13_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_2_LC_9_13_2  (
            .in0(N__23756),
            .in1(N__23779),
            .in2(N__23807),
            .in3(N__23759),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ),
            .clk(N__47270),
            .ce(N__23674),
            .sr(N__46687));
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_9_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_9_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_9_13_3 .LUT_INIT=16'b1101011101111101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_3_LC_9_13_3  (
            .in0(N__23754),
            .in1(N__23708),
            .in2(N__23735),
            .in3(N__23687),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ),
            .clk(N__47270),
            .ce(N__23674),
            .sr(N__46687));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_9_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_9_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_9_13_4  (
            .in0(_gnd_net_),
            .in1(N__23489),
            .in2(N__23462),
            .in3(N__23423),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_9_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_9_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_9_13_5  (
            .in0(_gnd_net_),
            .in1(N__24472),
            .in2(N__24442),
            .in3(N__24401),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_9_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_9_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_9_13_6  (
            .in0(_gnd_net_),
            .in1(N__24394),
            .in2(N__24365),
            .in3(N__24326),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_9_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_9_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_9_13_7  (
            .in0(_gnd_net_),
            .in1(N__24323),
            .in2(N__24298),
            .in3(N__24263),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_9_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_9_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_9_14_0  (
            .in0(_gnd_net_),
            .in1(N__24256),
            .in2(N__24235),
            .in3(N__24200),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(bfn_9_14_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_9_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_9_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(N__24188),
            .in2(N__24169),
            .in3(N__24134),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_9_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_9_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(N__24131),
            .in2(N__24101),
            .in3(N__24068),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_9_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_9_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(N__24065),
            .in2(N__24031),
            .in3(N__23993),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_9_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_9_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_9_14_4  (
            .in0(_gnd_net_),
            .in1(N__23988),
            .in2(N__23957),
            .in3(N__24986),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_9_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_9_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_9_14_5  (
            .in0(_gnd_net_),
            .in1(N__24971),
            .in2(N__24947),
            .in3(N__24914),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_9_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_9_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(N__24910),
            .in2(N__24879),
            .in3(N__24839),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_9_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_9_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_9_14_7  (
            .in0(_gnd_net_),
            .in1(N__24832),
            .in2(N__24796),
            .in3(N__24758),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_9_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_9_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_9_15_0  (
            .in0(_gnd_net_),
            .in1(N__24746),
            .in2(N__24719),
            .in3(N__24686),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(bfn_9_15_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_9_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_9_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(N__24679),
            .in2(N__24658),
            .in3(N__24623),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_9_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_9_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(N__24599),
            .in2(N__24578),
            .in3(N__24542),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_9_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_9_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(N__24535),
            .in2(N__24514),
            .in3(N__24479),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_9_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_9_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_9_15_4  (
            .in0(_gnd_net_),
            .in1(N__25462),
            .in2(N__25441),
            .in3(N__25406),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_9_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_9_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_9_15_5  (
            .in0(_gnd_net_),
            .in1(N__25386),
            .in2(N__25360),
            .in3(N__25325),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_9_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_9_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_9_15_6  (
            .in0(_gnd_net_),
            .in1(N__25316),
            .in2(N__25292),
            .in3(N__25262),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_9_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_9_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_9_15_7  (
            .in0(_gnd_net_),
            .in1(N__25258),
            .in2(N__25226),
            .in3(N__25187),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_9_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_9_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_9_16_0  (
            .in0(_gnd_net_),
            .in1(N__25176),
            .in2(N__25145),
            .in3(N__25109),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(bfn_9_16_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_9_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_9_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_9_16_1  (
            .in0(_gnd_net_),
            .in1(N__25101),
            .in2(N__25731),
            .in3(N__25058),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_9_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_9_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_9_16_2  (
            .in0(_gnd_net_),
            .in1(N__25720),
            .in2(N__25050),
            .in3(N__24995),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_9_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_9_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_9_16_3  (
            .in0(_gnd_net_),
            .in1(N__25950),
            .in2(N__25732),
            .in3(N__25910),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_9_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_9_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_9_16_4  (
            .in0(_gnd_net_),
            .in1(N__25724),
            .in2(N__25905),
            .in3(N__25856),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_9_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_9_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_9_16_5  (
            .in0(_gnd_net_),
            .in1(N__25847),
            .in2(N__25733),
            .in3(N__25799),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_9_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_9_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_9_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_9_16_6  (
            .in0(_gnd_net_),
            .in1(N__25728),
            .in2(N__25796),
            .in3(N__25736),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_9_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_9_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_9_16_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_9_16_7  (
            .in0(N__25729),
            .in1(N__25653),
            .in2(_gnd_net_),
            .in3(N__25493),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_1_c_RNO_LC_9_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_0_cry_1_c_RNO_LC_9_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_1_c_RNO_LC_9_17_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_1_c_RNO_LC_9_17_0  (
            .in0(N__30594),
            .in1(N__29614),
            .in2(_gnd_net_),
            .in3(N__27596),
            .lcout(\current_shift_inst.un38_control_input_0_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_2_LC_9_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_2_LC_9_17_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_2_LC_9_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_2_LC_9_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26423),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47236),
            .ce(N__26477),
            .sr(N__46715));
    defparam \current_shift_inst.un38_control_input_0_cry_3_c_inv_RNO_LC_9_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_0_cry_3_c_inv_RNO_LC_9_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_3_c_inv_RNO_LC_9_17_2 .LUT_INIT=16'b0101010101100101;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_3_c_inv_RNO_LC_9_17_2  (
            .in0(N__27526),
            .in1(N__27564),
            .in2(N__30603),
            .in3(N__27595),
            .lcout(\current_shift_inst.N_1717_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_1_LC_9_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_1_LC_9_17_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_1_LC_9_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_1_LC_9_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26456),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47236),
            .ce(N__26477),
            .sr(N__46715));
    defparam \current_shift_inst.un38_control_input_0_cry_2_c_RNO_LC_9_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_0_cry_2_c_RNO_LC_9_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_2_c_RNO_LC_9_17_4 .LUT_INIT=16'b1001101010011010;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_2_c_RNO_LC_9_17_4  (
            .in0(N__27568),
            .in1(N__27597),
            .in2(N__30604),
            .in3(N__29582),
            .lcout(\current_shift_inst.un38_control_input_0_cry_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5LGN1_3_LC_9_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5LGN1_3_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5LGN1_3_LC_9_17_5 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5LGN1_3_LC_9_17_5  (
            .in0(N__27598),
            .in1(N__27527),
            .in2(N__27569),
            .in3(N__30598),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3 ),
            .ltout(\current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_0_cry_4_c_RNO_LC_9_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_0_cry_4_c_RNO_LC_9_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_0_cry_4_c_RNO_LC_9_17_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.un38_control_input_0_cry_4_c_RNO_LC_9_17_6  (
            .in0(_gnd_net_),
            .in1(N__27486),
            .in2(N__26015),
            .in3(N__29529),
            .lcout(\current_shift_inst.un38_control_input_0_cry_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIK3CV_7_LC_9_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIK3CV_7_LC_9_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIK3CV_7_LC_9_18_0 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIK3CV_7_LC_9_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27758),
            .in3(N__29403),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIK3CV_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIP5T51_13_LC_9_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIP5T51_13_LC_9_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIP5T51_13_LC_9_18_1 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIP5T51_13_LC_9_18_1  (
            .in0(N__30271),
            .in1(N__29969),
            .in2(N__29933),
            .in3(N__30207),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIP5T51_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIER9V_5_LC_9_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIER9V_5_LC_9_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIER9V_5_LC_9_18_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIER9V_5_LC_9_18_2  (
            .in0(_gnd_net_),
            .in1(N__27853),
            .in2(_gnd_net_),
            .in3(N__29489),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIER9V_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJDBL1_10_LC_9_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJDBL1_10_LC_9_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJDBL1_10_LC_9_18_3 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJDBL1_10_LC_9_18_3  (
            .in0(N__27676),
            .in1(N__30074),
            .in2(N__30041),
            .in3(N__29736),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJDBL1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIE6961_18_LC_9_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIE6961_18_LC_9_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIE6961_18_LC_9_18_4 .LUT_INIT=16'b1001100110011001;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIE6961_18_LC_9_18_4  (
            .in0(N__30462),
            .in1(N__30424),
            .in2(N__27953),
            .in3(N__29645),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIE6961_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHVAV_6_LC_9_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHVAV_6_LC_9_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHVAV_6_LC_9_18_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHVAV_6_LC_9_18_5  (
            .in0(N__27798),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29451),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIHVAV_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7DM51_10_LC_9_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7DM51_10_LC_9_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7DM51_10_LC_9_18_6 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7DM51_10_LC_9_18_6  (
            .in0(N__29737),
            .in1(N__27677),
            .in2(N__30773),
            .in3(N__30715),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI7DM51_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI53NU1_6_LC_9_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI53NU1_6_LC_9_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI53NU1_6_LC_9_18_7 .LUT_INIT=16'b1100001111000011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI53NU1_6_LC_9_18_7  (
            .in0(N__27799),
            .in1(N__27752),
            .in2(N__29407),
            .in3(N__29452),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI53NU1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7H2J_17_LC_9_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7H2J_17_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7H2J_17_LC_9_19_0 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7H2J_17_LC_9_19_0  (
            .in0(N__29679),
            .in1(_gnd_net_),
            .in2(N__28000),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI7H2J_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIIKQI_10_LC_9_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIIKQI_10_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIIKQI_10_LC_9_19_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIIKQI_10_LC_9_19_1  (
            .in0(N__27675),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29738),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIIKQI_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU4VI_14_LC_9_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU4VI_14_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU4VI_14_LC_9_19_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU4VI_14_LC_9_19_2  (
            .in0(_gnd_net_),
            .in1(N__30270),
            .in2(_gnd_net_),
            .in3(N__30211),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIU4VI_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBU361_16_LC_9_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBU361_16_LC_9_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBU361_16_LC_9_19_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBU361_16_LC_9_19_3  (
            .in0(N__30320),
            .in1(N__27993),
            .in2(N__30358),
            .in3(N__29680),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIBU361_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBBPU1_7_LC_9_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBBPU1_7_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBBPU1_7_LC_9_19_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBBPU1_7_LC_9_19_5  (
            .in0(N__27756),
            .in1(N__29846),
            .in2(N__29414),
            .in3(N__29880),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIBBPU1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1PG21_9_LC_9_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1PG21_9_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1PG21_9_LC_9_19_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1PG21_9_LC_9_19_6  (
            .in0(_gnd_net_),
            .in1(N__30069),
            .in2(_gnd_net_),
            .in3(N__30037),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI1PG21_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNINKG81_27_LC_9_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNINKG81_27_LC_9_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNINKG81_27_LC_9_19_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNINKG81_27_LC_9_19_7  (
            .in0(N__28144),
            .in1(N__30879),
            .in2(N__30128),
            .in3(N__30838),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNINKG81_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR32K_22_LC_9_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR32K_22_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR32K_22_LC_9_20_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR32K_22_LC_9_20_0  (
            .in0(_gnd_net_),
            .in1(N__28249),
            .in2(_gnd_net_),
            .in3(N__29779),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIR32K_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPB581_22_LC_9_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPB581_22_LC_9_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPB581_22_LC_9_20_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPB581_22_LC_9_20_1  (
            .in0(N__28250),
            .in1(N__31544),
            .in2(N__29783),
            .in3(N__31588),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPB581_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJ3381_21_LC_9_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJ3381_21_LC_9_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJ3381_21_LC_9_20_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJ3381_21_LC_9_20_2  (
            .in0(N__30968),
            .in1(N__28248),
            .in2(N__31007),
            .in3(N__29778),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJ3381_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQF91_30_LC_9_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQF91_30_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQF91_30_LC_9_20_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQF91_30_LC_9_20_3  (
            .in0(N__31655),
            .in1(N__30631),
            .in2(_gnd_net_),
            .in3(N__30500),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIVQF91_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAO7K_27_LC_9_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAO7K_27_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAO7K_27_LC_9_20_4 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAO7K_27_LC_9_20_4  (
            .in0(N__30120),
            .in1(_gnd_net_),
            .in2(N__28145),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIAO7K_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4D1J_16_LC_9_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4D1J_16_LC_9_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4D1J_16_LC_9_20_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4D1J_16_LC_9_20_5  (
            .in0(_gnd_net_),
            .in1(N__30350),
            .in2(_gnd_net_),
            .in3(N__30319),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI4D1J_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIKKJ81_29_LC_9_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIKKJ81_29_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIKKJ81_29_LC_9_20_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIKKJ81_29_LC_9_20_6  (
            .in0(N__30883),
            .in1(N__31679),
            .in2(N__30842),
            .in3(N__31705),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIKKJ81_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHCE81_26_LC_9_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHCE81_26_LC_9_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHCE81_26_LC_9_20_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHCE81_26_LC_9_20_7  (
            .in0(N__31866),
            .in1(N__28140),
            .in2(N__31832),
            .in3(N__30121),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIHCE81_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_3_LC_9_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_3_LC_9_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_3_LC_9_21_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_3_LC_9_21_0  (
            .in0(_gnd_net_),
            .in1(N__26455),
            .in2(N__26398),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_3 ),
            .ltout(),
            .carryin(bfn_9_21_0_),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_2 ),
            .clk(N__47215),
            .ce(N__26476),
            .sr(N__46733));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_4_LC_9_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_4_LC_9_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_4_LC_9_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_4_LC_9_21_1  (
            .in0(_gnd_net_),
            .in1(N__26422),
            .in2(N__26371),
            .in3(N__26183),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_2 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_3 ),
            .clk(N__47215),
            .ce(N__26476),
            .sr(N__46733));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_5_LC_9_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_5_LC_9_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_5_LC_9_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_5_LC_9_21_2  (
            .in0(_gnd_net_),
            .in1(N__26341),
            .in2(N__26399),
            .in3(N__26180),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_3 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_4 ),
            .clk(N__47215),
            .ce(N__26476),
            .sr(N__46733));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_6_LC_9_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_6_LC_9_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_6_LC_9_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_6_LC_9_21_3  (
            .in0(_gnd_net_),
            .in1(N__26320),
            .in2(N__26372),
            .in3(N__26177),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_4 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_5 ),
            .clk(N__47215),
            .ce(N__26476),
            .sr(N__46733));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_7_LC_9_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_7_LC_9_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_7_LC_9_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_7_LC_9_21_4  (
            .in0(_gnd_net_),
            .in1(N__26342),
            .in2(N__26297),
            .in3(N__26174),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_5 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_6 ),
            .clk(N__47215),
            .ce(N__26476),
            .sr(N__46733));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_8_LC_9_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_8_LC_9_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_8_LC_9_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_8_LC_9_21_5  (
            .in0(_gnd_net_),
            .in1(N__26321),
            .in2(N__26263),
            .in3(N__26171),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_8 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_6 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_7 ),
            .clk(N__47215),
            .ce(N__26476),
            .sr(N__46733));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_9_LC_9_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_9_LC_9_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_9_LC_9_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_9_LC_9_21_6  (
            .in0(_gnd_net_),
            .in1(N__26296),
            .in2(N__26696),
            .in3(N__26168),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_7 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_8 ),
            .clk(N__47215),
            .ce(N__26476),
            .sr(N__46733));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_10_LC_9_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_10_LC_9_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_10_LC_9_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_10_LC_9_21_7  (
            .in0(_gnd_net_),
            .in1(N__26665),
            .in2(N__26264),
            .in3(N__26165),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_8 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_9 ),
            .clk(N__47215),
            .ce(N__26476),
            .sr(N__46733));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_11_LC_9_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_11_LC_9_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_11_LC_9_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_11_LC_9_22_0  (
            .in0(_gnd_net_),
            .in1(N__26695),
            .in2(N__26638),
            .in3(N__26162),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_11 ),
            .ltout(),
            .carryin(bfn_9_22_0_),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_10 ),
            .clk(N__47211),
            .ce(N__26475),
            .sr(N__46737));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_12_LC_9_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_12_LC_9_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_12_LC_9_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_12_LC_9_22_1  (
            .in0(_gnd_net_),
            .in1(N__26666),
            .in2(N__26608),
            .in3(N__26159),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_10 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_11 ),
            .clk(N__47211),
            .ce(N__26475),
            .sr(N__46737));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_13_LC_9_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_13_LC_9_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_13_LC_9_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_13_LC_9_22_2  (
            .in0(_gnd_net_),
            .in1(N__26581),
            .in2(N__26639),
            .in3(N__26210),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_11 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_12 ),
            .clk(N__47211),
            .ce(N__26475),
            .sr(N__46737));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_14_LC_9_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_14_LC_9_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_14_LC_9_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_14_LC_9_22_3  (
            .in0(_gnd_net_),
            .in1(N__26560),
            .in2(N__26609),
            .in3(N__26207),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_12 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_13 ),
            .clk(N__47211),
            .ce(N__26475),
            .sr(N__46737));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_15_LC_9_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_15_LC_9_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_15_LC_9_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_15_LC_9_22_4  (
            .in0(_gnd_net_),
            .in1(N__26582),
            .in2(N__26536),
            .in3(N__26204),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_13 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_14 ),
            .clk(N__47211),
            .ce(N__26475),
            .sr(N__46737));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_16_LC_9_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_16_LC_9_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_16_LC_9_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_16_LC_9_22_5  (
            .in0(_gnd_net_),
            .in1(N__26561),
            .in2(N__26509),
            .in3(N__26201),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_16 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_14 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_15 ),
            .clk(N__47211),
            .ce(N__26475),
            .sr(N__46737));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_17_LC_9_22_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_17_LC_9_22_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_17_LC_9_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_17_LC_9_22_6  (
            .in0(_gnd_net_),
            .in1(N__26914),
            .in2(N__26537),
            .in3(N__26198),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_15 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_16 ),
            .clk(N__47211),
            .ce(N__26475),
            .sr(N__46737));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_18_LC_9_22_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_18_LC_9_22_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_18_LC_9_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_18_LC_9_22_7  (
            .in0(_gnd_net_),
            .in1(N__26887),
            .in2(N__26510),
            .in3(N__26195),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_16 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_17 ),
            .clk(N__47211),
            .ce(N__26475),
            .sr(N__46737));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_19_LC_9_23_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_19_LC_9_23_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_19_LC_9_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_19_LC_9_23_0  (
            .in0(_gnd_net_),
            .in1(N__26915),
            .in2(N__26860),
            .in3(N__26192),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_19 ),
            .ltout(),
            .carryin(bfn_9_23_0_),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_18 ),
            .clk(N__47208),
            .ce(N__26474),
            .sr(N__46738));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_20_LC_9_23_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_20_LC_9_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_20_LC_9_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_20_LC_9_23_1  (
            .in0(_gnd_net_),
            .in1(N__26888),
            .in2(N__26830),
            .in3(N__26189),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_18 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_19 ),
            .clk(N__47208),
            .ce(N__26474),
            .sr(N__46738));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_21_LC_9_23_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_21_LC_9_23_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_21_LC_9_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_21_LC_9_23_2  (
            .in0(_gnd_net_),
            .in1(N__26800),
            .in2(N__26861),
            .in3(N__26186),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_19 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_20 ),
            .clk(N__47208),
            .ce(N__26474),
            .sr(N__46738));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_22_LC_9_23_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_22_LC_9_23_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_22_LC_9_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_22_LC_9_23_3  (
            .in0(_gnd_net_),
            .in1(N__26776),
            .in2(N__26831),
            .in3(N__26237),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_20 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_21 ),
            .clk(N__47208),
            .ce(N__26474),
            .sr(N__46738));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_23_LC_9_23_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_23_LC_9_23_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_23_LC_9_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_23_LC_9_23_4  (
            .in0(_gnd_net_),
            .in1(N__26801),
            .in2(N__26752),
            .in3(N__26234),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_21 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_22 ),
            .clk(N__47208),
            .ce(N__26474),
            .sr(N__46738));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_24_LC_9_23_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_24_LC_9_23_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_24_LC_9_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_24_LC_9_23_5  (
            .in0(_gnd_net_),
            .in1(N__26777),
            .in2(N__26722),
            .in3(N__26231),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_24 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_22 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_23 ),
            .clk(N__47208),
            .ce(N__26474),
            .sr(N__46738));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_25_LC_9_23_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_25_LC_9_23_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_25_LC_9_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_25_LC_9_23_6  (
            .in0(_gnd_net_),
            .in1(N__27070),
            .in2(N__26753),
            .in3(N__26228),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_23 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_24 ),
            .clk(N__47208),
            .ce(N__26474),
            .sr(N__46738));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_26_LC_9_23_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_26_LC_9_23_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_26_LC_9_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_26_LC_9_23_7  (
            .in0(_gnd_net_),
            .in1(N__27043),
            .in2(N__26723),
            .in3(N__26225),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_24 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_25 ),
            .clk(N__47208),
            .ce(N__26474),
            .sr(N__46738));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_27_LC_9_24_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_27_LC_9_24_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_27_LC_9_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_27_LC_9_24_0  (
            .in0(_gnd_net_),
            .in1(N__27071),
            .in2(N__27016),
            .in3(N__26222),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_27 ),
            .ltout(),
            .carryin(bfn_9_24_0_),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_26 ),
            .clk(N__47204),
            .ce(N__26473),
            .sr(N__46740));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_28_LC_9_24_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_28_LC_9_24_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_28_LC_9_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_28_LC_9_24_1  (
            .in0(_gnd_net_),
            .in1(N__27044),
            .in2(N__26986),
            .in3(N__26219),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_26 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_27 ),
            .clk(N__47204),
            .ce(N__26473),
            .sr(N__46740));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_29_LC_9_24_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_29_LC_9_24_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_29_LC_9_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_29_LC_9_24_2  (
            .in0(_gnd_net_),
            .in1(N__26960),
            .in2(N__27017),
            .in3(N__26216),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_29 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_27 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_28 ),
            .clk(N__47204),
            .ce(N__26473),
            .sr(N__46740));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_30_LC_9_24_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_30_LC_9_24_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_30_LC_9_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_30_LC_9_24_3  (
            .in0(_gnd_net_),
            .in1(N__26936),
            .in2(N__26987),
            .in3(N__26213),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_30 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_28 ),
            .carryout(\current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_29 ),
            .clk(N__47204),
            .ce(N__26473),
            .sr(N__46740));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_31_LC_9_24_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_31_LC_9_24_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_31_LC_9_24_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_31_LC_9_24_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26480),
            .lcout(\current_shift_inst.elapsed_time_ns_phase_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47204),
            .ce(N__26473),
            .sr(N__46740));
    defparam \current_shift_inst.timer_phase.counter_0_LC_9_25_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_0_LC_9_25_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_0_LC_9_25_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_0_LC_9_25_0  (
            .in0(N__32081),
            .in1(N__26442),
            .in2(_gnd_net_),
            .in3(N__26426),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_9_25_0_),
            .carryout(\current_shift_inst.timer_phase.counter_cry_0 ),
            .clk(N__47199),
            .ce(N__32134),
            .sr(N__46741));
    defparam \current_shift_inst.timer_phase.counter_1_LC_9_25_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_1_LC_9_25_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_1_LC_9_25_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_1_LC_9_25_1  (
            .in0(N__32077),
            .in1(N__26415),
            .in2(_gnd_net_),
            .in3(N__26402),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_0 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_1 ),
            .clk(N__47199),
            .ce(N__32134),
            .sr(N__46741));
    defparam \current_shift_inst.timer_phase.counter_2_LC_9_25_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_2_LC_9_25_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_2_LC_9_25_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_2_LC_9_25_2  (
            .in0(N__32082),
            .in1(N__26391),
            .in2(_gnd_net_),
            .in3(N__26375),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_1 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_2 ),
            .clk(N__47199),
            .ce(N__32134),
            .sr(N__46741));
    defparam \current_shift_inst.timer_phase.counter_3_LC_9_25_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_3_LC_9_25_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_3_LC_9_25_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_3_LC_9_25_3  (
            .in0(N__32078),
            .in1(N__26359),
            .in2(_gnd_net_),
            .in3(N__26345),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_2 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_3 ),
            .clk(N__47199),
            .ce(N__32134),
            .sr(N__46741));
    defparam \current_shift_inst.timer_phase.counter_4_LC_9_25_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_4_LC_9_25_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_4_LC_9_25_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_4_LC_9_25_4  (
            .in0(N__32083),
            .in1(N__26340),
            .in2(_gnd_net_),
            .in3(N__26324),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_3 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_4 ),
            .clk(N__47199),
            .ce(N__32134),
            .sr(N__46741));
    defparam \current_shift_inst.timer_phase.counter_5_LC_9_25_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_5_LC_9_25_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_5_LC_9_25_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_5_LC_9_25_5  (
            .in0(N__32079),
            .in1(N__26314),
            .in2(_gnd_net_),
            .in3(N__26300),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_4 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_5 ),
            .clk(N__47199),
            .ce(N__32134),
            .sr(N__46741));
    defparam \current_shift_inst.timer_phase.counter_6_LC_9_25_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_6_LC_9_25_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_6_LC_9_25_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_6_LC_9_25_6  (
            .in0(N__32084),
            .in1(N__26286),
            .in2(_gnd_net_),
            .in3(N__26267),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_5 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_6 ),
            .clk(N__47199),
            .ce(N__32134),
            .sr(N__46741));
    defparam \current_shift_inst.timer_phase.counter_7_LC_9_25_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_7_LC_9_25_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_7_LC_9_25_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_7_LC_9_25_7  (
            .in0(N__32080),
            .in1(N__26256),
            .in2(_gnd_net_),
            .in3(N__26240),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_6 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_7 ),
            .clk(N__47199),
            .ce(N__32134),
            .sr(N__46741));
    defparam \current_shift_inst.timer_phase.counter_8_LC_9_26_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_8_LC_9_26_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_8_LC_9_26_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_8_LC_9_26_0  (
            .in0(N__32064),
            .in1(N__26685),
            .in2(_gnd_net_),
            .in3(N__26669),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_9_26_0_),
            .carryout(\current_shift_inst.timer_phase.counter_cry_8 ),
            .clk(N__47197),
            .ce(N__32126),
            .sr(N__46742));
    defparam \current_shift_inst.timer_phase.counter_9_LC_9_26_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_9_LC_9_26_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_9_LC_9_26_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_9_LC_9_26_1  (
            .in0(N__32068),
            .in1(N__26658),
            .in2(_gnd_net_),
            .in3(N__26642),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_8 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_9 ),
            .clk(N__47197),
            .ce(N__32126),
            .sr(N__46742));
    defparam \current_shift_inst.timer_phase.counter_10_LC_9_26_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_10_LC_9_26_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_10_LC_9_26_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_10_LC_9_26_2  (
            .in0(N__32061),
            .in1(N__26626),
            .in2(_gnd_net_),
            .in3(N__26612),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_9 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_10 ),
            .clk(N__47197),
            .ce(N__32126),
            .sr(N__46742));
    defparam \current_shift_inst.timer_phase.counter_11_LC_9_26_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_11_LC_9_26_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_11_LC_9_26_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_11_LC_9_26_3  (
            .in0(N__32065),
            .in1(N__26601),
            .in2(_gnd_net_),
            .in3(N__26585),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_10 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_11 ),
            .clk(N__47197),
            .ce(N__32126),
            .sr(N__46742));
    defparam \current_shift_inst.timer_phase.counter_12_LC_9_26_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_12_LC_9_26_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_12_LC_9_26_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_12_LC_9_26_4  (
            .in0(N__32062),
            .in1(N__26580),
            .in2(_gnd_net_),
            .in3(N__26564),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_11 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_12 ),
            .clk(N__47197),
            .ce(N__32126),
            .sr(N__46742));
    defparam \current_shift_inst.timer_phase.counter_13_LC_9_26_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_13_LC_9_26_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_13_LC_9_26_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_13_LC_9_26_5  (
            .in0(N__32066),
            .in1(N__26554),
            .in2(_gnd_net_),
            .in3(N__26540),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_12 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_13 ),
            .clk(N__47197),
            .ce(N__32126),
            .sr(N__46742));
    defparam \current_shift_inst.timer_phase.counter_14_LC_9_26_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_14_LC_9_26_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_14_LC_9_26_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_14_LC_9_26_6  (
            .in0(N__32063),
            .in1(N__26529),
            .in2(_gnd_net_),
            .in3(N__26513),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_13 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_14 ),
            .clk(N__47197),
            .ce(N__32126),
            .sr(N__46742));
    defparam \current_shift_inst.timer_phase.counter_15_LC_9_26_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_15_LC_9_26_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_15_LC_9_26_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_15_LC_9_26_7  (
            .in0(N__32067),
            .in1(N__26497),
            .in2(_gnd_net_),
            .in3(N__26483),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_14 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_15 ),
            .clk(N__47197),
            .ce(N__32126),
            .sr(N__46742));
    defparam \current_shift_inst.timer_phase.counter_16_LC_9_27_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_16_LC_9_27_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_16_LC_9_27_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_16_LC_9_27_0  (
            .in0(N__32069),
            .in1(N__26907),
            .in2(_gnd_net_),
            .in3(N__26891),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_9_27_0_),
            .carryout(\current_shift_inst.timer_phase.counter_cry_16 ),
            .clk(N__47195),
            .ce(N__32135),
            .sr(N__46744));
    defparam \current_shift_inst.timer_phase.counter_17_LC_9_27_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_17_LC_9_27_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_17_LC_9_27_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_17_LC_9_27_1  (
            .in0(N__32073),
            .in1(N__26880),
            .in2(_gnd_net_),
            .in3(N__26864),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_16 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_17 ),
            .clk(N__47195),
            .ce(N__32135),
            .sr(N__46744));
    defparam \current_shift_inst.timer_phase.counter_18_LC_9_27_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_18_LC_9_27_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_18_LC_9_27_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_18_LC_9_27_2  (
            .in0(N__32070),
            .in1(N__26848),
            .in2(_gnd_net_),
            .in3(N__26834),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_17 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_18 ),
            .clk(N__47195),
            .ce(N__32135),
            .sr(N__46744));
    defparam \current_shift_inst.timer_phase.counter_19_LC_9_27_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_19_LC_9_27_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_19_LC_9_27_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_19_LC_9_27_3  (
            .in0(N__32074),
            .in1(N__26818),
            .in2(_gnd_net_),
            .in3(N__26804),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_18 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_19 ),
            .clk(N__47195),
            .ce(N__32135),
            .sr(N__46744));
    defparam \current_shift_inst.timer_phase.counter_20_LC_9_27_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_20_LC_9_27_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_20_LC_9_27_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_20_LC_9_27_4  (
            .in0(N__32071),
            .in1(N__26794),
            .in2(_gnd_net_),
            .in3(N__26780),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_19 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_20 ),
            .clk(N__47195),
            .ce(N__32135),
            .sr(N__46744));
    defparam \current_shift_inst.timer_phase.counter_21_LC_9_27_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_21_LC_9_27_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_21_LC_9_27_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_21_LC_9_27_5  (
            .in0(N__32075),
            .in1(N__26770),
            .in2(_gnd_net_),
            .in3(N__26756),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_20 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_21 ),
            .clk(N__47195),
            .ce(N__32135),
            .sr(N__46744));
    defparam \current_shift_inst.timer_phase.counter_22_LC_9_27_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_22_LC_9_27_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_22_LC_9_27_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_22_LC_9_27_6  (
            .in0(N__32072),
            .in1(N__26740),
            .in2(_gnd_net_),
            .in3(N__26726),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_21 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_22 ),
            .clk(N__47195),
            .ce(N__32135),
            .sr(N__46744));
    defparam \current_shift_inst.timer_phase.counter_23_LC_9_27_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_23_LC_9_27_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_23_LC_9_27_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_23_LC_9_27_7  (
            .in0(N__32076),
            .in1(N__26715),
            .in2(_gnd_net_),
            .in3(N__26699),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_22 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_23 ),
            .clk(N__47195),
            .ce(N__32135),
            .sr(N__46744));
    defparam \current_shift_inst.timer_phase.counter_24_LC_9_28_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_24_LC_9_28_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_24_LC_9_28_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_24_LC_9_28_0  (
            .in0(N__32085),
            .in1(N__27063),
            .in2(_gnd_net_),
            .in3(N__27047),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_9_28_0_),
            .carryout(\current_shift_inst.timer_phase.counter_cry_24 ),
            .clk(N__47193),
            .ce(N__32133),
            .sr(N__46745));
    defparam \current_shift_inst.timer_phase.counter_25_LC_9_28_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_25_LC_9_28_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_25_LC_9_28_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_25_LC_9_28_1  (
            .in0(N__32089),
            .in1(N__27036),
            .in2(_gnd_net_),
            .in3(N__27020),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_24 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_25 ),
            .clk(N__47193),
            .ce(N__32133),
            .sr(N__46745));
    defparam \current_shift_inst.timer_phase.counter_26_LC_9_28_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_26_LC_9_28_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_26_LC_9_28_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_26_LC_9_28_2  (
            .in0(N__32086),
            .in1(N__27004),
            .in2(_gnd_net_),
            .in3(N__26990),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_25 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_26 ),
            .clk(N__47193),
            .ce(N__32133),
            .sr(N__46745));
    defparam \current_shift_inst.timer_phase.counter_27_LC_9_28_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_27_LC_9_28_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_27_LC_9_28_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_27_LC_9_28_3  (
            .in0(N__32090),
            .in1(N__26979),
            .in2(_gnd_net_),
            .in3(N__26963),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_26 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_27 ),
            .clk(N__47193),
            .ce(N__32133),
            .sr(N__46745));
    defparam \current_shift_inst.timer_phase.counter_28_LC_9_28_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_phase.counter_28_LC_9_28_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_28_LC_9_28_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_phase.counter_28_LC_9_28_4  (
            .in0(N__32087),
            .in1(N__26956),
            .in2(_gnd_net_),
            .in3(N__26942),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_phase.counter_cry_27 ),
            .carryout(\current_shift_inst.timer_phase.counter_cry_28 ),
            .clk(N__47193),
            .ce(N__32133),
            .sr(N__46745));
    defparam \current_shift_inst.timer_phase.counter_29_LC_9_28_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.counter_29_LC_9_28_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.counter_29_LC_9_28_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \current_shift_inst.timer_phase.counter_29_LC_9_28_5  (
            .in0(N__26935),
            .in1(N__32088),
            .in2(_gnd_net_),
            .in3(N__26939),
            .lcout(\current_shift_inst.timer_phase.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47193),
            .ce(N__32133),
            .sr(N__46745));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_10_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_10_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_10_7_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_10_7_0  (
            .in0(_gnd_net_),
            .in1(N__27397),
            .in2(_gnd_net_),
            .in3(N__40067),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MAX_D2_LC_10_7_7.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_10_7_7.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_10_7_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MAX_D2_LC_10_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26921),
            .lcout(il_max_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47308),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_10_8_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_10_8_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pwm_generator_inst.counter_RNISQD2_0_LC_10_8_0  (
            .in0(_gnd_net_),
            .in1(N__27153),
            .in2(_gnd_net_),
            .in3(N__27195),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlto2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_10_8_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_10_8_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_10_8_1 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \pwm_generator_inst.counter_RNIBO26_1_LC_10_8_1  (
            .in0(N__27112),
            .in1(N__27133),
            .in2(N__27209),
            .in3(N__27175),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlt9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_10_8_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_10_8_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIFA6C_5_LC_10_8_2  (
            .in0(N__27203),
            .in1(N__27347),
            .in2(N__27206),
            .in3(N__27092),
            .lcout(\pwm_generator_inst.un1_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_10_8_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_10_8_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_10_8_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIVDL3_9_LC_10_8_7  (
            .in0(N__27230),
            .in1(N__27305),
            .in2(_gnd_net_),
            .in3(N__27325),
            .lcout(\pwm_generator_inst.un1_counterlto9_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_0_LC_10_9_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_0_LC_10_9_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_0_LC_10_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_0_LC_10_9_0  (
            .in0(N__27276),
            .in1(N__27197),
            .in2(_gnd_net_),
            .in3(N__27179),
            .lcout(\pwm_generator_inst.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_10_9_0_),
            .carryout(\pwm_generator_inst.counter_cry_0 ),
            .clk(N__47288),
            .ce(),
            .sr(N__46638));
    defparam \pwm_generator_inst.counter_1_LC_10_9_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_1_LC_10_9_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_1_LC_10_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_1_LC_10_9_1  (
            .in0(N__27272),
            .in1(N__27176),
            .in2(_gnd_net_),
            .in3(N__27158),
            .lcout(\pwm_generator_inst.counterZ0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_0 ),
            .carryout(\pwm_generator_inst.counter_cry_1 ),
            .clk(N__47288),
            .ce(),
            .sr(N__46638));
    defparam \pwm_generator_inst.counter_2_LC_10_9_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_2_LC_10_9_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_2_LC_10_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_2_LC_10_9_2  (
            .in0(N__27277),
            .in1(N__27155),
            .in2(_gnd_net_),
            .in3(N__27137),
            .lcout(\pwm_generator_inst.counterZ0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_1 ),
            .carryout(\pwm_generator_inst.counter_cry_2 ),
            .clk(N__47288),
            .ce(),
            .sr(N__46638));
    defparam \pwm_generator_inst.counter_3_LC_10_9_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_3_LC_10_9_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_3_LC_10_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_3_LC_10_9_3  (
            .in0(N__27273),
            .in1(N__27134),
            .in2(_gnd_net_),
            .in3(N__27116),
            .lcout(\pwm_generator_inst.counterZ0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_2 ),
            .carryout(\pwm_generator_inst.counter_cry_3 ),
            .clk(N__47288),
            .ce(),
            .sr(N__46638));
    defparam \pwm_generator_inst.counter_4_LC_10_9_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_4_LC_10_9_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_4_LC_10_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_4_LC_10_9_4  (
            .in0(N__27278),
            .in1(N__27113),
            .in2(_gnd_net_),
            .in3(N__27095),
            .lcout(\pwm_generator_inst.counterZ0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_3 ),
            .carryout(\pwm_generator_inst.counter_cry_4 ),
            .clk(N__47288),
            .ce(),
            .sr(N__46638));
    defparam \pwm_generator_inst.counter_5_LC_10_9_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_5_LC_10_9_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_5_LC_10_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_5_LC_10_9_5  (
            .in0(N__27274),
            .in1(N__27091),
            .in2(_gnd_net_),
            .in3(N__27074),
            .lcout(\pwm_generator_inst.counterZ0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_4 ),
            .carryout(\pwm_generator_inst.counter_cry_5 ),
            .clk(N__47288),
            .ce(),
            .sr(N__46638));
    defparam \pwm_generator_inst.counter_6_LC_10_9_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_6_LC_10_9_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_6_LC_10_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_6_LC_10_9_6  (
            .in0(N__27279),
            .in1(N__27346),
            .in2(_gnd_net_),
            .in3(N__27329),
            .lcout(\pwm_generator_inst.counterZ0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_5 ),
            .carryout(\pwm_generator_inst.counter_cry_6 ),
            .clk(N__47288),
            .ce(),
            .sr(N__46638));
    defparam \pwm_generator_inst.counter_7_LC_10_9_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_7_LC_10_9_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_7_LC_10_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_7_LC_10_9_7  (
            .in0(N__27275),
            .in1(N__27326),
            .in2(_gnd_net_),
            .in3(N__27308),
            .lcout(\pwm_generator_inst.counterZ0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_6 ),
            .carryout(\pwm_generator_inst.counter_cry_7 ),
            .clk(N__47288),
            .ce(),
            .sr(N__46638));
    defparam \pwm_generator_inst.counter_8_LC_10_10_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_8_LC_10_10_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_8_LC_10_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_8_LC_10_10_0  (
            .in0(N__27281),
            .in1(N__27304),
            .in2(_gnd_net_),
            .in3(N__27284),
            .lcout(\pwm_generator_inst.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_10_10_0_),
            .carryout(\pwm_generator_inst.counter_cry_8 ),
            .clk(N__47281),
            .ce(),
            .sr(N__46645));
    defparam \pwm_generator_inst.counter_9_LC_10_10_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_9_LC_10_10_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_9_LC_10_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_9_LC_10_10_1  (
            .in0(N__27280),
            .in1(N__27229),
            .in2(_gnd_net_),
            .in3(N__27233),
            .lcout(\pwm_generator_inst.counterZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47281),
            .ce(),
            .sr(N__46645));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_10_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_10_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_10_10_2 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_10_10_2  (
            .in0(N__39662),
            .in1(N__39978),
            .in2(N__39848),
            .in3(N__28895),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47281),
            .ce(),
            .sr(N__46645));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_10_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_10_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_10_10_3 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_10_10_3  (
            .in0(N__39820),
            .in1(N__39667),
            .in2(N__40014),
            .in3(N__29207),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47281),
            .ce(),
            .sr(N__46645));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_10_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_10_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_10_10_4 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_10_10_4  (
            .in0(N__39663),
            .in1(N__39988),
            .in2(N__39849),
            .in3(N__29180),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47281),
            .ce(),
            .sr(N__46645));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_10_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_10_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_10_10_5 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_10_10_5  (
            .in0(N__39819),
            .in1(N__39666),
            .in2(N__40013),
            .in3(N__29264),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47281),
            .ce(),
            .sr(N__46645));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_10_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_10_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_10_10_6 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_10_10_6  (
            .in0(N__39664),
            .in1(N__39989),
            .in2(N__39850),
            .in3(N__29096),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47281),
            .ce(),
            .sr(N__46645));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_10_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_10_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_10_10_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_10_10_7  (
            .in0(N__39818),
            .in1(N__39665),
            .in2(N__40012),
            .in3(N__28865),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47281),
            .ce(),
            .sr(N__46645));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_10_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_10_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_10_11_2 .LUT_INIT=16'b1100100010001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_10_11_2  (
            .in0(N__39811),
            .in1(N__29126),
            .in2(N__39680),
            .in3(N__39932),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47272),
            .ce(),
            .sr(N__46653));
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_10_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_10_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_10_11_4 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_LC_10_11_4  (
            .in0(N__31106),
            .in1(N__27398),
            .in2(N__27368),
            .in3(N__40064),
            .lcout(\phase_controller_inst1.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47272),
            .ce(),
            .sr(N__46653));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_10_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_10_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_10_11_5 .LUT_INIT=16'b1100110010000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_10_11_5  (
            .in0(N__39669),
            .in1(N__29153),
            .in2(N__39977),
            .in3(N__39812),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47272),
            .ce(),
            .sr(N__46653));
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_10_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_10_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_10_12_1 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_14_LC_10_12_1  (
            .in0(N__43899),
            .in1(N__44087),
            .in2(_gnd_net_),
            .in3(N__33878),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47262),
            .ce(N__31225),
            .sr(N__46663));
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_10_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_10_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_10_12_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_11_LC_10_12_4  (
            .in0(N__44086),
            .in1(N__39352),
            .in2(_gnd_net_),
            .in3(N__43898),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47262),
            .ce(N__31225),
            .sr(N__46663));
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_10_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_10_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_10_12_6 .LUT_INIT=16'b0000010000000101;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_9_LC_10_12_6  (
            .in0(N__40344),
            .in1(N__34048),
            .in2(N__44155),
            .in3(N__43900),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47262),
            .ce(N__31225),
            .sr(N__46663));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_10_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_10_13_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_10_13_1  (
            .in0(_gnd_net_),
            .in1(N__39608),
            .in2(_gnd_net_),
            .in3(N__39766),
            .lcout(\phase_controller_inst1.stoper_hc.time_passed11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_10_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_10_13_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_10_13_3  (
            .in0(N__39961),
            .in1(N__39609),
            .in2(_gnd_net_),
            .in3(N__39767),
            .lcout(\phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_0_c_inv_LC_10_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_0_c_inv_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_0_c_inv_LC_10_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_0_c_inv_LC_10_14_0  (
            .in0(_gnd_net_),
            .in1(N__29293),
            .in2(N__27356),
            .in3(N__29325),
            .lcout(G_407),
            .ltout(),
            .carryin(bfn_10_14_0_),
            .carryout(\current_shift_inst.z_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_1_c_inv_LC_10_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_1_c_inv_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_1_c_inv_LC_10_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_1_c_inv_LC_10_14_1  (
            .in0(_gnd_net_),
            .in1(N__27443),
            .in2(N__29604),
            .in3(N__27599),
            .lcout(G_406),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_0 ),
            .carryout(\current_shift_inst.z_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_2_c_LC_10_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_2_c_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_2_c_LC_10_14_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_2_c_LC_10_14_2  (
            .in0(_gnd_net_),
            .in1(N__29569),
            .in2(N__27545),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_1 ),
            .carryout(\current_shift_inst.z_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_3_c_LC_10_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_3_c_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_3_c_LC_10_14_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_3_c_LC_10_14_3  (
            .in0(_gnd_net_),
            .in1(N__29548),
            .in2(N__27506),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_2 ),
            .carryout(\current_shift_inst.z_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_4_c_LC_10_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_4_c_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_4_c_LC_10_14_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_4_c_LC_10_14_4  (
            .in0(_gnd_net_),
            .in1(N__27458),
            .in2(N__29519),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_3 ),
            .carryout(\current_shift_inst.z_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_5_c_LC_10_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_5_c_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_5_c_LC_10_14_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_5_c_LC_10_14_5  (
            .in0(_gnd_net_),
            .in1(N__29472),
            .in2(N__27821),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_4 ),
            .carryout(\current_shift_inst.z_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_6_c_LC_10_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_6_c_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_6_c_LC_10_14_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_6_c_LC_10_14_6  (
            .in0(_gnd_net_),
            .in1(N__27773),
            .in2(N__29442),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_5 ),
            .carryout(\current_shift_inst.z_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_7_c_LC_10_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_7_c_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_7_c_LC_10_14_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_7_c_LC_10_14_7  (
            .in0(_gnd_net_),
            .in1(N__27722),
            .in2(N__29391),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_6 ),
            .carryout(\current_shift_inst.z_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_8_c_LC_10_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_8_c_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_8_c_LC_10_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_8_c_LC_10_15_0  (
            .in0(_gnd_net_),
            .in1(N__27707),
            .in2(N__29837),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_15_0_),
            .carryout(\current_shift_inst.z_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_9_c_LC_10_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_9_c_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_9_c_LC_10_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_9_c_LC_10_15_1  (
            .in0(_gnd_net_),
            .in1(N__27692),
            .in2(N__30029),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_8 ),
            .carryout(\current_shift_inst.z_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_10_c_LC_10_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_10_c_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_10_c_LC_10_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_10_c_LC_10_15_2  (
            .in0(_gnd_net_),
            .in1(N__29721),
            .in2(N__27650),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_9 ),
            .carryout(\current_shift_inst.z_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_11_c_LC_10_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_11_c_LC_10_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_11_c_LC_10_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_11_c_LC_10_15_3  (
            .in0(_gnd_net_),
            .in1(N__27632),
            .in2(N__30707),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_10 ),
            .carryout(\current_shift_inst.z_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_12_c_LC_10_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_12_c_LC_10_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_12_c_LC_10_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_12_c_LC_10_15_4  (
            .in0(_gnd_net_),
            .in1(N__27617),
            .in2(N__30737),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_11 ),
            .carryout(\current_shift_inst.z_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_13_c_LC_10_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_13_c_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_13_c_LC_10_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_13_c_LC_10_15_5  (
            .in0(_gnd_net_),
            .in1(N__28064),
            .in2(N__29921),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_12 ),
            .carryout(\current_shift_inst.z_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_14_c_LC_10_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_14_c_LC_10_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_14_c_LC_10_15_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_14_c_LC_10_15_6  (
            .in0(_gnd_net_),
            .in1(N__28049),
            .in2(N__30197),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_13 ),
            .carryout(\current_shift_inst.z_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_15_c_LC_10_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_15_c_LC_10_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_15_c_LC_10_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_15_c_LC_10_15_7  (
            .in0(_gnd_net_),
            .in1(N__28034),
            .in2(N__30233),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_14 ),
            .carryout(\current_shift_inst.z_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_16_c_LC_10_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_16_c_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_16_c_LC_10_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_16_c_LC_10_16_0  (
            .in0(_gnd_net_),
            .in1(N__30303),
            .in2(N__28019),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_16_0_),
            .carryout(\current_shift_inst.z_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_17_c_LC_10_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_17_c_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_17_c_LC_10_16_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_17_c_LC_10_16_1  (
            .in0(_gnd_net_),
            .in1(N__27968),
            .in2(N__29670),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_16 ),
            .carryout(\current_shift_inst.z_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_18_c_LC_10_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_18_c_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_18_c_LC_10_16_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_18_c_LC_10_16_2  (
            .in0(_gnd_net_),
            .in1(N__29631),
            .in2(N__27920),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_17 ),
            .carryout(\current_shift_inst.z_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_19_c_LC_10_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_19_c_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_19_c_LC_10_16_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_19_c_LC_10_16_3  (
            .in0(_gnd_net_),
            .in1(N__27902),
            .in2(N__30416),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_18 ),
            .carryout(\current_shift_inst.z_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_20_c_LC_10_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_20_c_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_20_c_LC_10_16_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_20_c_LC_10_16_4  (
            .in0(_gnd_net_),
            .in1(N__27887),
            .in2(N__31070),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_19 ),
            .carryout(\current_shift_inst.z_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_21_c_LC_10_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_21_c_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_21_c_LC_10_16_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_21_c_LC_10_16_5  (
            .in0(_gnd_net_),
            .in1(N__30954),
            .in2(N__27872),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_20 ),
            .carryout(\current_shift_inst.z_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_22_c_LC_10_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_22_c_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_22_c_LC_10_16_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_22_c_LC_10_16_6  (
            .in0(_gnd_net_),
            .in1(N__28226),
            .in2(N__29770),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_21 ),
            .carryout(\current_shift_inst.z_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_23_c_LC_10_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_23_c_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_23_c_LC_10_16_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_23_c_LC_10_16_7  (
            .in0(_gnd_net_),
            .in1(N__31572),
            .in2(N__28211),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_22 ),
            .carryout(\current_shift_inst.z_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_24_c_LC_10_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_24_c_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_24_c_LC_10_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_24_c_LC_10_17_0  (
            .in0(_gnd_net_),
            .in1(N__28193),
            .in2(N__31507),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_17_0_),
            .carryout(\current_shift_inst.z_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_25_c_LC_10_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_25_c_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_25_c_LC_10_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_25_c_LC_10_17_1  (
            .in0(_gnd_net_),
            .in1(N__31748),
            .in2(N__28178),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_24 ),
            .carryout(\current_shift_inst.z_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_26_c_LC_10_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_26_c_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_26_c_LC_10_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_26_c_LC_10_17_2  (
            .in0(_gnd_net_),
            .in1(N__28160),
            .in2(N__31824),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_25 ),
            .carryout(\current_shift_inst.z_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_27_c_LC_10_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_27_c_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_27_c_LC_10_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_27_c_LC_10_17_3  (
            .in0(_gnd_net_),
            .in1(N__28112),
            .in2(N__30111),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_26 ),
            .carryout(\current_shift_inst.z_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_28_c_LC_10_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_28_c_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_28_c_LC_10_17_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_28_c_LC_10_17_4  (
            .in0(_gnd_net_),
            .in1(N__28097),
            .in2(N__30831),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_27 ),
            .carryout(\current_shift_inst.z_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_29_c_LC_10_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_29_c_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_29_c_LC_10_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_29_c_LC_10_17_5  (
            .in0(_gnd_net_),
            .in1(N__31671),
            .in2(N__28082),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_28 ),
            .carryout(\current_shift_inst.z_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_cry_30_c_LC_10_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_cry_30_c_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_cry_30_c_LC_10_17_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_cry_30_c_LC_10_17_6  (
            .in0(_gnd_net_),
            .in1(N__30489),
            .in2(N__28469),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.z_cry_29 ),
            .carryout(\current_shift_inst.z_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_s_31_LC_10_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_z_s_31_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_s_31_LC_10_17_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \current_shift_inst.un10_control_input_z_s_31_LC_10_17_7  (
            .in0(N__30574),
            .in1(N__28448),
            .in2(N__30529),
            .in3(N__27602),
            .lcout(\current_shift_inst.z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_1_c_LC_10_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_1_c_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_1_c_LC_10_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_1_c_LC_10_18_0  (
            .in0(_gnd_net_),
            .in1(N__27591),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_18_0_),
            .carryout(\current_shift_inst.z_5_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_2_s_LC_10_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_2_s_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_2_s_LC_10_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_2_s_LC_10_18_1  (
            .in0(_gnd_net_),
            .in1(N__27563),
            .in2(N__28693),
            .in3(N__27530),
            .lcout(\current_shift_inst.z_5_2 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_1 ),
            .carryout(\current_shift_inst.z_5_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_3_s_LC_10_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_3_s_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_3_s_LC_10_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_3_s_LC_10_18_2  (
            .in0(_gnd_net_),
            .in1(N__27520),
            .in2(N__28697),
            .in3(N__27491),
            .lcout(\current_shift_inst.z_5_3 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_2 ),
            .carryout(\current_shift_inst.z_5_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_4_s_LC_10_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_4_s_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_4_s_LC_10_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_4_s_LC_10_18_3  (
            .in0(_gnd_net_),
            .in1(N__27485),
            .in2(N__28694),
            .in3(N__27446),
            .lcout(\current_shift_inst.z_5_4 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_3 ),
            .carryout(\current_shift_inst.z_5_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_5_s_LC_10_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_5_s_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_5_s_LC_10_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_5_s_LC_10_18_4  (
            .in0(_gnd_net_),
            .in1(N__27842),
            .in2(N__28698),
            .in3(N__27806),
            .lcout(\current_shift_inst.z_5_5 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_4 ),
            .carryout(\current_shift_inst.z_5_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_6_s_LC_10_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_6_s_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_6_s_LC_10_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_6_s_LC_10_18_5  (
            .in0(_gnd_net_),
            .in1(N__27797),
            .in2(N__28695),
            .in3(N__27761),
            .lcout(\current_shift_inst.z_5_6 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_5 ),
            .carryout(\current_shift_inst.z_5_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_7_s_LC_10_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_7_s_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_7_s_LC_10_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_7_s_LC_10_18_6  (
            .in0(_gnd_net_),
            .in1(N__27757),
            .in2(N__28699),
            .in3(N__27710),
            .lcout(\current_shift_inst.z_5_7 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_6 ),
            .carryout(\current_shift_inst.z_5_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_8_s_LC_10_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_8_s_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_8_s_LC_10_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_8_s_LC_10_18_7  (
            .in0(_gnd_net_),
            .in1(N__29873),
            .in2(N__28696),
            .in3(N__27695),
            .lcout(\current_shift_inst.z_5_8 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_7 ),
            .carryout(\current_shift_inst.z_5_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_9_s_LC_10_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_9_s_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_9_s_LC_10_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_9_s_LC_10_19_0  (
            .in0(_gnd_net_),
            .in1(N__30065),
            .in2(N__28847),
            .in3(N__27680),
            .lcout(\current_shift_inst.z_5_9 ),
            .ltout(),
            .carryin(bfn_10_19_0_),
            .carryout(\current_shift_inst.z_5_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_10_s_LC_10_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_10_s_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_10_s_LC_10_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_10_s_LC_10_19_1  (
            .in0(_gnd_net_),
            .in1(N__27674),
            .in2(N__28841),
            .in3(N__27635),
            .lcout(\current_shift_inst.z_5_10 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_9 ),
            .carryout(\current_shift_inst.z_5_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_11_s_LC_10_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_11_s_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_11_s_LC_10_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_11_s_LC_10_19_2  (
            .in0(_gnd_net_),
            .in1(N__30762),
            .in2(N__28844),
            .in3(N__27620),
            .lcout(\current_shift_inst.z_5_11 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_10 ),
            .carryout(\current_shift_inst.z_5_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_12_s_LC_10_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_12_s_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_12_s_LC_10_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_12_s_LC_10_19_3  (
            .in0(_gnd_net_),
            .in1(N__30663),
            .in2(N__28842),
            .in3(N__27605),
            .lcout(\current_shift_inst.z_5_12 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_11 ),
            .carryout(\current_shift_inst.z_5_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_13_s_LC_10_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_13_s_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_13_s_LC_10_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_13_s_LC_10_19_4  (
            .in0(_gnd_net_),
            .in1(N__29957),
            .in2(N__28845),
            .in3(N__28052),
            .lcout(\current_shift_inst.z_5_13 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_12 ),
            .carryout(\current_shift_inst.z_5_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_14_s_LC_10_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_14_s_LC_10_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_14_s_LC_10_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_14_s_LC_10_19_5  (
            .in0(_gnd_net_),
            .in1(N__30269),
            .in2(N__28843),
            .in3(N__28037),
            .lcout(\current_shift_inst.z_5_14 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_13 ),
            .carryout(\current_shift_inst.z_5_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_15_s_LC_10_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_15_s_LC_10_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_15_s_LC_10_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_15_s_LC_10_19_6  (
            .in0(_gnd_net_),
            .in1(N__30164),
            .in2(N__28846),
            .in3(N__28022),
            .lcout(\current_shift_inst.z_5_15 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_14 ),
            .carryout(\current_shift_inst.z_5_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_16_s_LC_10_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_16_s_LC_10_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_16_s_LC_10_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_16_s_LC_10_19_7  (
            .in0(_gnd_net_),
            .in1(N__28792),
            .in2(N__30357),
            .in3(N__28004),
            .lcout(\current_shift_inst.z_5_16 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_15 ),
            .carryout(\current_shift_inst.z_5_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_17_s_LC_10_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_17_s_LC_10_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_17_s_LC_10_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_17_s_LC_10_20_0  (
            .in0(_gnd_net_),
            .in1(N__27992),
            .in2(N__28833),
            .in3(N__27956),
            .lcout(\current_shift_inst.z_5_17 ),
            .ltout(),
            .carryin(bfn_10_20_0_),
            .carryout(\current_shift_inst.z_5_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_18_s_LC_10_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_18_s_LC_10_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_18_s_LC_10_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_18_s_LC_10_20_1  (
            .in0(_gnd_net_),
            .in1(N__27939),
            .in2(N__28837),
            .in3(N__27905),
            .lcout(\current_shift_inst.z_5_18 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_17 ),
            .carryout(\current_shift_inst.z_5_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_19_s_LC_10_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_19_s_LC_10_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_19_s_LC_10_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_19_s_LC_10_20_2  (
            .in0(_gnd_net_),
            .in1(N__30452),
            .in2(N__28834),
            .in3(N__27890),
            .lcout(\current_shift_inst.z_5_19 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_18 ),
            .carryout(\current_shift_inst.z_5_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_20_s_LC_10_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_20_s_LC_10_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_20_s_LC_10_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_20_s_LC_10_20_3  (
            .in0(_gnd_net_),
            .in1(N__31033),
            .in2(N__28838),
            .in3(N__27875),
            .lcout(\current_shift_inst.z_5_20 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_19 ),
            .carryout(\current_shift_inst.z_5_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_21_s_LC_10_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_21_s_LC_10_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_21_s_LC_10_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_21_s_LC_10_20_4  (
            .in0(_gnd_net_),
            .in1(N__30992),
            .in2(N__28835),
            .in3(N__28253),
            .lcout(\current_shift_inst.z_5_21 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_20 ),
            .carryout(\current_shift_inst.z_5_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_22_s_LC_10_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_22_s_LC_10_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_22_s_LC_10_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_22_s_LC_10_20_5  (
            .in0(_gnd_net_),
            .in1(N__28247),
            .in2(N__28839),
            .in3(N__28214),
            .lcout(\current_shift_inst.z_5_22 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_21 ),
            .carryout(\current_shift_inst.z_5_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_23_s_LC_10_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_23_s_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_23_s_LC_10_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_23_s_LC_10_20_6  (
            .in0(_gnd_net_),
            .in1(N__31548),
            .in2(N__28836),
            .in3(N__28196),
            .lcout(\current_shift_inst.z_5_23 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_22 ),
            .carryout(\current_shift_inst.z_5_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_24_s_LC_10_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_24_s_LC_10_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_24_s_LC_10_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_24_s_LC_10_20_7  (
            .in0(_gnd_net_),
            .in1(N__31622),
            .in2(N__28840),
            .in3(N__28181),
            .lcout(\current_shift_inst.z_5_24 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_23 ),
            .carryout(\current_shift_inst.z_5_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_25_s_LC_10_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_25_s_LC_10_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_25_s_LC_10_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_25_s_LC_10_21_0  (
            .in0(_gnd_net_),
            .in1(N__31768),
            .in2(N__28827),
            .in3(N__28163),
            .lcout(\current_shift_inst.z_5_25 ),
            .ltout(),
            .carryin(bfn_10_21_0_),
            .carryout(\current_shift_inst.z_5_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_26_s_LC_10_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_26_s_LC_10_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_26_s_LC_10_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_26_s_LC_10_21_1  (
            .in0(_gnd_net_),
            .in1(N__31859),
            .in2(N__28830),
            .in3(N__28148),
            .lcout(\current_shift_inst.z_5_26 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_25 ),
            .carryout(\current_shift_inst.z_5_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_27_s_LC_10_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_27_s_LC_10_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_27_s_LC_10_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_27_s_LC_10_21_2  (
            .in0(_gnd_net_),
            .in1(N__28139),
            .in2(N__28828),
            .in3(N__28100),
            .lcout(\current_shift_inst.z_5_27 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_26 ),
            .carryout(\current_shift_inst.z_5_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_28_s_LC_10_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_28_s_LC_10_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_28_s_LC_10_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_28_s_LC_10_21_3  (
            .in0(_gnd_net_),
            .in1(N__30869),
            .in2(N__28831),
            .in3(N__28085),
            .lcout(\current_shift_inst.z_5_28 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_27 ),
            .carryout(\current_shift_inst.z_5_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_29_s_LC_10_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_29_s_LC_10_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_29_s_LC_10_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_29_s_LC_10_21_4  (
            .in0(_gnd_net_),
            .in1(N__31704),
            .in2(N__28829),
            .in3(N__28067),
            .lcout(\current_shift_inst.z_5_29 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_28 ),
            .carryout(\current_shift_inst.z_5_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_5_cry_30_s_LC_10_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_z_5_cry_30_s_LC_10_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_5_cry_30_s_LC_10_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un10_control_input_z_5_cry_30_s_LC_10_21_5  (
            .in0(_gnd_net_),
            .in1(N__30630),
            .in2(N__28832),
            .in3(N__28454),
            .lcout(\current_shift_inst.z_5_30 ),
            .ltout(),
            .carryin(\current_shift_inst.z_5_cry_29 ),
            .carryout(\current_shift_inst.z_5_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.z_5_cry_30_THRU_LUT4_0_LC_10_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.z_5_cry_30_THRU_LUT4_0_LC_10_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.z_5_cry_30_THRU_LUT4_0_LC_10_21_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.z_5_cry_30_THRU_LUT4_0_LC_10_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28451),
            .lcout(\current_shift_inst.z_5_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.S2_LC_10_28_3 .C_ON=1'b0;
    defparam \phase_controller_slave.S2_LC_10_28_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.S2_LC_10_28_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.S2_LC_10_28_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32255),
            .lcout(s4_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47190),
            .ce(),
            .sr(N__46743));
    defparam SB_DFF_inst_PH1_MIN_D1_LC_11_6_6.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_11_6_6.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_11_6_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MIN_D1_LC_11_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28421),
            .lcout(il_min_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47309),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_11_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_11_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_11_8_0  (
            .in0(_gnd_net_),
            .in1(N__28406),
            .in2(N__28391),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_8_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_11_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_11_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(N__28361),
            .in2(_gnd_net_),
            .in3(N__28331),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_11_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_11_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_11_8_2  (
            .in0(_gnd_net_),
            .in1(N__28328),
            .in2(N__28322),
            .in3(N__28289),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_11_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_11_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_11_8_3  (
            .in0(_gnd_net_),
            .in1(N__28286),
            .in2(_gnd_net_),
            .in3(N__28256),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_11_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_11_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_11_8_4  (
            .in0(_gnd_net_),
            .in1(N__29081),
            .in2(_gnd_net_),
            .in3(N__29051),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_11_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_11_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_11_8_5  (
            .in0(_gnd_net_),
            .in1(N__29048),
            .in2(_gnd_net_),
            .in3(N__29018),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_11_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_11_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_11_8_6  (
            .in0(_gnd_net_),
            .in1(N__29015),
            .in2(_gnd_net_),
            .in3(N__28985),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_11_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_11_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_11_8_7  (
            .in0(_gnd_net_),
            .in1(N__28982),
            .in2(_gnd_net_),
            .in3(N__28952),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_11_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_11_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(N__31138),
            .in2(_gnd_net_),
            .in3(N__28949),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_11_9_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_11_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_11_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(N__28946),
            .in2(_gnd_net_),
            .in3(N__28919),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_11_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_11_9_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_11_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28915),
            .in3(N__28889),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_11_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_11_9_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28885),
            .in3(N__28859),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_11_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_11_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(N__29278),
            .in2(_gnd_net_),
            .in3(N__29258),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_11_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_11_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_11_9_5  (
            .in0(_gnd_net_),
            .in1(N__29255),
            .in2(_gnd_net_),
            .in3(N__29228),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_11_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_11_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_11_9_6  (
            .in0(_gnd_net_),
            .in1(N__29221),
            .in2(_gnd_net_),
            .in3(N__29201),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_11_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_11_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_11_9_7  (
            .in0(_gnd_net_),
            .in1(N__29194),
            .in2(_gnd_net_),
            .in3(N__29174),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_11_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_11_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_11_10_0  (
            .in0(_gnd_net_),
            .in1(N__29167),
            .in2(_gnd_net_),
            .in3(N__29147),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(bfn_11_10_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_11_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_11_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_11_10_1  (
            .in0(_gnd_net_),
            .in1(N__29140),
            .in2(_gnd_net_),
            .in3(N__29120),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_11_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_11_10_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_11_10_2  (
            .in0(_gnd_net_),
            .in1(N__29113),
            .in2(_gnd_net_),
            .in3(N__29099),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MIN_D2_LC_11_10_6.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_11_10_6.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_11_10_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MIN_D2_LC_11_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29090),
            .lcout(il_min_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47273),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_6_LC_11_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_6_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_6_LC_11_11_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_6_LC_11_11_2  (
            .in0(N__34150),
            .in1(N__34047),
            .in2(_gnd_net_),
            .in3(N__35431),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_10_LC_11_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_10_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_10_LC_11_11_3 .LUT_INIT=16'b0101000001110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_10_LC_11_11_3  (
            .in0(N__35513),
            .in1(N__34107),
            .in2(N__29357),
            .in3(N__41253),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_11_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_11_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_11_12_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_15_LC_11_12_2  (
            .in0(N__44084),
            .in1(N__33916),
            .in2(_gnd_net_),
            .in3(N__43878),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47253),
            .ce(N__31229),
            .sr(N__46654));
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_11_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_11_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_11_12_7 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_18_LC_11_12_7  (
            .in0(N__43879),
            .in1(N__44085),
            .in2(_gnd_net_),
            .in3(N__42191),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47253),
            .ce(N__31229),
            .sr(N__46654));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_11_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_11_13_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_11_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_11_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35854),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47245),
            .ce(N__32738),
            .sr(N__46664));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_11_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_11_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_11_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_11_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35827),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47245),
            .ce(N__32738),
            .sr(N__46664));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_11_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_11_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_11_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_11_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32716),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47245),
            .ce(N__32738),
            .sr(N__46664));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_11_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_11_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_11_13_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_11_13_3  (
            .in0(N__32717),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_1_fast_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47245),
            .ce(N__32738),
            .sr(N__46664));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_RNI48NB_31_LC_11_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_RNI48NB_31_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_RNI48NB_31_LC_11_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_RNI48NB_31_LC_11_14_0  (
            .in0(_gnd_net_),
            .in1(N__31328),
            .in2(N__29327),
            .in3(N__29326),
            .lcout(\current_shift_inst.un38_control_input_0 ),
            .ltout(),
            .carryin(bfn_11_14_0_),
            .carryout(\current_shift_inst.un4_control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_1_c_RNIJF2G_LC_11_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_1_c_RNIJF2G_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_1_c_RNIJF2G_LC_11_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_1_c_RNIJF2G_LC_11_14_1  (
            .in0(_gnd_net_),
            .in1(N__31316),
            .in2(_gnd_net_),
            .in3(N__29585),
            .lcout(\current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_1 ),
            .carryout(\current_shift_inst.un4_control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_2_c_RNILI3G_LC_11_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_2_c_RNILI3G_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_2_c_RNILI3G_LC_11_14_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.un4_control_input_cry_2_c_RNILI3G_LC_11_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31163),
            .in3(N__29558),
            .lcout(\current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_2 ),
            .carryout(\current_shift_inst.un4_control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_3_c_RNINL4G_LC_11_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_3_c_RNINL4G_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_3_c_RNINL4G_LC_11_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_3_c_RNINL4G_LC_11_14_3  (
            .in0(_gnd_net_),
            .in1(N__31154),
            .in2(_gnd_net_),
            .in3(N__29537),
            .lcout(\current_shift_inst.un4_control_input_cry_3_c_RNINL4GZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_3 ),
            .carryout(\current_shift_inst.un4_control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_4_c_RNIPO5G_LC_11_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_4_c_RNIPO5G_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_4_c_RNIPO5G_LC_11_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_4_c_RNIPO5G_LC_11_14_4  (
            .in0(_gnd_net_),
            .in1(N__31298),
            .in2(_gnd_net_),
            .in3(N__29492),
            .lcout(\current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_4 ),
            .carryout(\current_shift_inst.un4_control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_5_c_RNIRR6G_LC_11_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_5_c_RNIRR6G_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_5_c_RNIRR6G_LC_11_14_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.un4_control_input_cry_5_c_RNIRR6G_LC_11_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31289),
            .in3(N__29456),
            .lcout(\current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_5 ),
            .carryout(\current_shift_inst.un4_control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_6_c_RNITU7G_LC_11_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_6_c_RNITU7G_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_6_c_RNITU7G_LC_11_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_6_c_RNITU7G_LC_11_14_6  (
            .in0(_gnd_net_),
            .in1(N__31277),
            .in2(_gnd_net_),
            .in3(N__29417),
            .lcout(\current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_6 ),
            .carryout(\current_shift_inst.un4_control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_7_c_RNIV19G_LC_11_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_7_c_RNIV19G_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_7_c_RNIV19G_LC_11_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_7_c_RNIV19G_LC_11_14_7  (
            .in0(_gnd_net_),
            .in1(N__33749),
            .in2(_gnd_net_),
            .in3(N__29366),
            .lcout(\current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_7 ),
            .carryout(\current_shift_inst.un4_control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_8_c_RNI15AG_LC_11_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_8_c_RNI15AG_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_8_c_RNI15AG_LC_11_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_8_c_RNI15AG_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(N__33980),
            .in2(_gnd_net_),
            .in3(N__29363),
            .lcout(\current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0 ),
            .ltout(),
            .carryin(bfn_11_15_0_),
            .carryout(\current_shift_inst.un4_control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_9_c_RNIALDJ_LC_11_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_9_c_RNIALDJ_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_9_c_RNIALDJ_LC_11_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_9_c_RNIALDJ_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(N__31376),
            .in2(_gnd_net_),
            .in3(N__29360),
            .lcout(\current_shift_inst.un4_control_input_cry_9_c_RNIALDJZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_9 ),
            .carryout(\current_shift_inst.un4_control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_10_c_RNIJLTG_LC_11_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_10_c_RNIJLTG_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_10_c_RNIJLTG_LC_11_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_10_c_RNIJLTG_LC_11_15_2  (
            .in0(_gnd_net_),
            .in1(N__31391),
            .in2(_gnd_net_),
            .in3(N__29705),
            .lcout(\current_shift_inst.un4_control_input_cry_10_c_RNIJLTGZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_10 ),
            .carryout(\current_shift_inst.un4_control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_11_c_RNILOUG_LC_11_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_11_c_RNILOUG_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_11_c_RNILOUG_LC_11_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_11_c_RNILOUG_LC_11_15_3  (
            .in0(_gnd_net_),
            .in1(N__31370),
            .in2(_gnd_net_),
            .in3(N__29702),
            .lcout(\current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_11 ),
            .carryout(\current_shift_inst.un4_control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_12_c_RNINRVG_LC_11_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_12_c_RNINRVG_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_12_c_RNINRVG_LC_11_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_12_c_RNINRVG_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(N__33926),
            .in2(_gnd_net_),
            .in3(N__29699),
            .lcout(\current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_12 ),
            .carryout(\current_shift_inst.un4_control_input_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_13_c_RNIPU0H_LC_11_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_13_c_RNIPU0H_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_13_c_RNIPU0H_LC_11_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_13_c_RNIPU0H_LC_11_15_5  (
            .in0(_gnd_net_),
            .in1(N__31364),
            .in2(_gnd_net_),
            .in3(N__29696),
            .lcout(\current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_13 ),
            .carryout(\current_shift_inst.un4_control_input_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_14_c_RNIR12H_LC_11_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_14_c_RNIR12H_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_14_c_RNIR12H_LC_11_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_14_c_RNIR12H_LC_11_15_6  (
            .in0(_gnd_net_),
            .in1(N__31304),
            .in2(_gnd_net_),
            .in3(N__29693),
            .lcout(\current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_14 ),
            .carryout(\current_shift_inst.un4_control_input_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_15_c_RNIT43H_LC_11_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_15_c_RNIT43H_LC_11_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_15_c_RNIT43H_LC_11_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_15_c_RNIT43H_LC_11_15_7  (
            .in0(_gnd_net_),
            .in1(N__33962),
            .in2(_gnd_net_),
            .in3(N__29690),
            .lcout(\current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_15 ),
            .carryout(\current_shift_inst.un4_control_input_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_16_c_RNIV74H_LC_11_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_16_c_RNIV74H_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_16_c_RNIV74H_LC_11_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_16_c_RNIV74H_LC_11_16_0  (
            .in0(_gnd_net_),
            .in1(N__33944),
            .in2(_gnd_net_),
            .in3(N__29687),
            .lcout(\current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0 ),
            .ltout(),
            .carryin(bfn_11_16_0_),
            .carryout(\current_shift_inst.un4_control_input_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_17_c_RNI1B5H_LC_11_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_17_c_RNI1B5H_LC_11_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_17_c_RNI1B5H_LC_11_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_17_c_RNI1B5H_LC_11_16_1  (
            .in0(_gnd_net_),
            .in1(N__31358),
            .in2(_gnd_net_),
            .in3(N__29648),
            .lcout(\current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_17 ),
            .carryout(\current_shift_inst.un4_control_input_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_18_c_RNI3E6H_LC_11_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_18_c_RNI3E6H_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_18_c_RNI3E6H_LC_11_16_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.un4_control_input_cry_18_c_RNI3E6H_LC_11_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31385),
            .in3(N__29795),
            .lcout(\current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_18 ),
            .carryout(\current_shift_inst.un4_control_input_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_19_c_RNIS88H_LC_11_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_19_c_RNIS88H_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_19_c_RNIS88H_LC_11_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_19_c_RNIS88H_LC_11_16_3  (
            .in0(_gnd_net_),
            .in1(N__31442),
            .in2(_gnd_net_),
            .in3(N__29792),
            .lcout(\current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_19 ),
            .carryout(\current_shift_inst.un4_control_input_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_20_c_RNILQ1I_LC_11_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_20_c_RNILQ1I_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_20_c_RNILQ1I_LC_11_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_20_c_RNILQ1I_LC_11_16_4  (
            .in0(_gnd_net_),
            .in1(N__31454),
            .in2(_gnd_net_),
            .in3(N__29789),
            .lcout(\current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_20 ),
            .carryout(\current_shift_inst.un4_control_input_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_21_c_RNINT2I_LC_11_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_21_c_RNINT2I_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_21_c_RNINT2I_LC_11_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_21_c_RNINT2I_LC_11_16_5  (
            .in0(_gnd_net_),
            .in1(N__31346),
            .in2(_gnd_net_),
            .in3(N__29786),
            .lcout(\current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_21 ),
            .carryout(\current_shift_inst.un4_control_input_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_22_c_RNIP04I_LC_11_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_22_c_RNIP04I_LC_11_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_22_c_RNIP04I_LC_11_16_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_22_c_RNIP04I_LC_11_16_6  (
            .in0(_gnd_net_),
            .in1(N__33734),
            .in2(_gnd_net_),
            .in3(N__29753),
            .lcout(\current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_22 ),
            .carryout(\current_shift_inst.un4_control_input_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_23_c_RNIR35I_LC_11_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_23_c_RNIR35I_LC_11_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_23_c_RNIR35I_LC_11_16_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_23_c_RNIR35I_LC_11_16_7  (
            .in0(_gnd_net_),
            .in1(N__31310),
            .in2(_gnd_net_),
            .in3(N__29750),
            .lcout(\current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_23 ),
            .carryout(\current_shift_inst.un4_control_input_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_24_c_RNIT66I_LC_11_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_24_c_RNIT66I_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_24_c_RNIT66I_LC_11_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_24_c_RNIT66I_LC_11_17_0  (
            .in0(_gnd_net_),
            .in1(N__31448),
            .in2(_gnd_net_),
            .in3(N__29747),
            .lcout(\current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0 ),
            .ltout(),
            .carryin(bfn_11_17_0_),
            .carryout(\current_shift_inst.un4_control_input_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_25_c_RNIV97I_LC_11_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_25_c_RNIV97I_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_25_c_RNIV97I_LC_11_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_25_c_RNIV97I_LC_11_17_1  (
            .in0(_gnd_net_),
            .in1(N__31340),
            .in2(_gnd_net_),
            .in3(N__29744),
            .lcout(\current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_25 ),
            .carryout(\current_shift_inst.un4_control_input_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_26_c_RNI1D8I_LC_11_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_26_c_RNI1D8I_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_26_c_RNI1D8I_LC_11_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_26_c_RNI1D8I_LC_11_17_2  (
            .in0(_gnd_net_),
            .in1(N__31466),
            .in2(_gnd_net_),
            .in3(N__29741),
            .lcout(\current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_26 ),
            .carryout(\current_shift_inst.un4_control_input_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_27_c_RNI3G9I_LC_11_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_27_c_RNI3G9I_LC_11_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_27_c_RNI3G9I_LC_11_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_27_c_RNI3G9I_LC_11_17_3  (
            .in0(_gnd_net_),
            .in1(N__31397),
            .in2(_gnd_net_),
            .in3(N__30086),
            .lcout(\current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_27 ),
            .carryout(\current_shift_inst.un4_control_input_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_28_c_RNI5JAI_LC_11_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_28_c_RNI5JAI_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_28_c_RNI5JAI_LC_11_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_28_c_RNI5JAI_LC_11_17_4  (
            .in0(_gnd_net_),
            .in1(N__31352),
            .in2(_gnd_net_),
            .in3(N__30083),
            .lcout(\current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_28 ),
            .carryout(\current_shift_inst.un4_control_input_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_29_c_RNIUDCI_LC_11_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_cry_29_c_RNIUDCI_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_29_c_RNIUDCI_LC_11_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_cry_29_c_RNIUDCI_LC_11_17_5  (
            .in0(_gnd_net_),
            .in1(N__31460),
            .in2(_gnd_net_),
            .in3(N__30080),
            .lcout(\current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_cry_29 ),
            .carryout(\current_shift_inst.un4_control_input_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_cry_30_c_RNINV5J_LC_11_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_cry_30_c_RNINV5J_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_cry_30_c_RNINV5J_LC_11_17_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.un4_control_input_cry_30_c_RNINV5J_LC_11_17_6  (
            .in0(_gnd_net_),
            .in1(N__30560),
            .in2(_gnd_net_),
            .in3(N__30077),
            .lcout(\current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIO0U12_8_LC_11_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIO0U12_8_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIO0U12_8_LC_11_18_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIO0U12_8_LC_11_18_0  (
            .in0(N__29882),
            .in1(N__30073),
            .in2(N__29845),
            .in3(N__30030),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIO0U12_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILORI_11_LC_11_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILORI_11_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILORI_11_LC_11_18_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILORI_11_LC_11_18_1  (
            .in0(N__30771),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30708),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNILORI_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOSSI_12_LC_11_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOSSI_12_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOSSI_12_LC_11_18_2 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOSSI_12_LC_11_18_2  (
            .in0(N__30739),
            .in1(_gnd_net_),
            .in2(N__30679),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIOSSI_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJTQ51_12_LC_11_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJTQ51_12_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJTQ51_12_LC_11_18_3 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJTQ51_12_LC_11_18_3  (
            .in0(N__29967),
            .in1(N__30740),
            .in2(N__30680),
            .in3(N__29925),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJTQ51_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIN7DV_8_LC_11_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIN7DV_8_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIN7DV_8_LC_11_18_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIN7DV_8_LC_11_18_4  (
            .in0(_gnd_net_),
            .in1(N__29881),
            .in2(_gnd_net_),
            .in3(N__29838),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIN7DV_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDS8K_28_LC_11_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDS8K_28_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDS8K_28_LC_11_18_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDS8K_28_LC_11_18_5  (
            .in0(_gnd_net_),
            .in1(N__30884),
            .in2(_gnd_net_),
            .in3(N__30827),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIDS8K_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5S981_24_LC_11_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5S981_24_LC_11_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5S981_24_LC_11_18_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5S981_24_LC_11_18_6  (
            .in0(N__31628),
            .in1(N__31749),
            .in2(N__31508),
            .in3(N__31784),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5S981_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDLO51_11_LC_11_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDLO51_11_LC_11_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDLO51_11_LC_11_18_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDLO51_11_LC_11_18_7  (
            .in0(N__30772),
            .in1(N__30738),
            .in2(N__30716),
            .in3(N__30672),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIDLO51_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_RNO_0_25_LC_11_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_RNO_0_25_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_RNO_0_25_LC_11_19_0 .LUT_INIT=16'b1100001110010110;
    LogicCell40 \current_shift_inst.control_input_RNO_0_25_LC_11_19_0  (
            .in0(N__30638),
            .in1(N__30590),
            .in2(N__30533),
            .in3(N__30499),
            .lcout(\current_shift_inst.un38_control_input_0_axb_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPC571_19_LC_11_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPC571_19_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPC571_19_LC_11_19_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPC571_19_LC_11_19_1  (
            .in0(N__30464),
            .in1(N__31041),
            .in2(N__30425),
            .in3(N__31071),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPC571_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI190J_15_LC_11_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI190J_15_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI190J_15_LC_11_19_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI190J_15_LC_11_19_2  (
            .in0(_gnd_net_),
            .in1(N__30166),
            .in2(_gnd_net_),
            .in3(N__30234),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI190J_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5M161_15_LC_11_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5M161_15_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5M161_15_LC_11_19_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5M161_15_LC_11_19_3  (
            .in0(N__30167),
            .in1(N__30359),
            .in2(N__30239),
            .in3(N__30312),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5M161_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVDV51_14_LC_11_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVDV51_14_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVDV51_14_LC_11_19_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVDV51_14_LC_11_19_4  (
            .in0(N__30278),
            .in1(N__30235),
            .in2(N__30212),
            .in3(N__30165),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIVDV51_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDR081_20_LC_11_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDR081_20_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDR081_20_LC_11_19_5 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDR081_20_LC_11_19_5  (
            .in0(N__31003),
            .in1(N__31045),
            .in2(N__31076),
            .in3(N__30963),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIDR081_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILRVJ_20_LC_11_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILRVJ_20_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILRVJ_20_LC_11_19_6 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILRVJ_20_LC_11_19_6  (
            .in0(N__31072),
            .in1(_gnd_net_),
            .in2(N__31046),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNILRVJ_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOV0K_21_LC_11_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOV0K_21_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOV0K_21_LC_11_19_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOV0K_21_LC_11_19_7  (
            .in0(_gnd_net_),
            .in1(N__31002),
            .in2(_gnd_net_),
            .in3(N__30964),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIOV0K_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU73K_23_LC_11_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU73K_23_LC_11_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU73K_23_LC_11_20_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU73K_23_LC_11_20_2  (
            .in0(_gnd_net_),
            .in1(N__31549),
            .in2(_gnd_net_),
            .in3(N__31592),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIU73K_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.start_timer_tr_RNO_1_LC_11_20_3 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_tr_RNO_1_LC_11_20_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.start_timer_tr_RNO_1_LC_11_20_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.start_timer_tr_RNO_1_LC_11_20_3  (
            .in0(_gnd_net_),
            .in1(N__32250),
            .in2(_gnd_net_),
            .in3(N__32217),
            .lcout(\phase_controller_slave.start_timer_tr_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7K6K_26_LC_11_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7K6K_26_LC_11_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7K6K_26_LC_11_20_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7K6K_26_LC_11_20_5  (
            .in0(_gnd_net_),
            .in1(N__31867),
            .in2(_gnd_net_),
            .in3(N__31825),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI7K6K_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MAX_D2_LC_11_21_7.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MAX_D2_LC_11_21_7.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MAX_D2_LC_11_21_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MAX_D2_LC_11_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30899),
            .lcout(il_max_comp2_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47205),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.state_1_LC_11_22_2 .C_ON=1'b0;
    defparam \phase_controller_slave.state_1_LC_11_22_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.state_1_LC_11_22_2 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \phase_controller_slave.state_1_LC_11_22_2  (
            .in0(N__32218),
            .in1(N__47637),
            .in2(N__32251),
            .in3(N__47665),
            .lcout(\phase_controller_slave.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47201),
            .ce(),
            .sr(N__46725));
    defparam \delay_measurement_inst.delay_hc_reg_6_LC_12_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_6_LC_12_9_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_6_LC_12_9_0 .LUT_INIT=16'b1011100011111111;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_6_LC_12_9_0  (
            .in0(N__35129),
            .in1(N__42648),
            .in2(N__34158),
            .in3(N__42102),
            .lcout(measured_delay_hc_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47271),
            .ce(),
            .sr(N__46627));
    defparam \phase_controller_inst1.state_1_LC_12_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_1_LC_12_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_1_LC_12_10_0 .LUT_INIT=16'b1100000011101010;
    LogicCell40 \phase_controller_inst1.state_1_LC_12_10_0  (
            .in0(N__43076),
            .in1(N__31115),
            .in2(N__33787),
            .in3(N__43023),
            .lcout(\phase_controller_inst1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47261),
            .ce(),
            .sr(N__46633));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_12_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_12_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_12_10_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_12_10_2  (
            .in0(N__39668),
            .in1(N__39768),
            .in2(N__39928),
            .in3(N__31148),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47261),
            .ce(),
            .sr(N__46633));
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_12_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_12_11_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_1_LC_12_11_0  (
            .in0(_gnd_net_),
            .in1(N__32504),
            .in2(_gnd_net_),
            .in3(N__32538),
            .lcout(),
            .ltout(\phase_controller_inst1.start_timer_hc_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_LC_12_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_LC_12_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_hc_LC_12_11_1 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \phase_controller_inst1.start_timer_hc_LC_12_11_1  (
            .in0(N__43153),
            .in1(N__39910),
            .in2(N__31124),
            .in3(N__31121),
            .lcout(\phase_controller_inst1.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47252),
            .ce(),
            .sr(N__46639));
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_12_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_12_11_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_0_LC_12_11_2  (
            .in0(_gnd_net_),
            .in1(N__33773),
            .in2(_gnd_net_),
            .in3(N__31110),
            .lcout(\phase_controller_inst1.N_88 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_2_LC_12_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_2_LC_12_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_2_LC_12_11_3 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \phase_controller_inst1.state_2_LC_12_11_3  (
            .in0(N__31111),
            .in1(N__32505),
            .in2(N__33783),
            .in3(N__32539),
            .lcout(\phase_controller_inst1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47252),
            .ce(),
            .sr(N__46639));
    defparam \phase_controller_slave.stoper_tr.target_time_10_LC_12_12_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_10_LC_12_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_10_LC_12_12_0 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_10_LC_12_12_0  (
            .in0(N__47598),
            .in1(N__39473),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47244),
            .ce(N__44417),
            .sr(N__46646));
    defparam \phase_controller_slave.stoper_tr.target_time_11_LC_12_12_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_11_LC_12_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_11_LC_12_12_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_11_LC_12_12_1  (
            .in0(_gnd_net_),
            .in1(N__47595),
            .in2(_gnd_net_),
            .in3(N__41531),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47244),
            .ce(N__44417),
            .sr(N__46646));
    defparam \phase_controller_slave.stoper_tr.target_time_12_LC_12_12_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_12_LC_12_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_12_LC_12_12_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_12_LC_12_12_2  (
            .in0(N__47596),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39500),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47244),
            .ce(N__44417),
            .sr(N__46646));
    defparam \phase_controller_slave.stoper_tr.target_time_13_LC_12_12_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_13_LC_12_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_13_LC_12_12_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_13_LC_12_12_3  (
            .in0(N__41999),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47597),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47244),
            .ce(N__44417),
            .sr(N__46646));
    defparam \phase_controller_slave.stoper_tr.target_time_15_LC_12_12_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_15_LC_12_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_15_LC_12_12_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_15_LC_12_12_4  (
            .in0(_gnd_net_),
            .in1(N__41489),
            .in2(_gnd_net_),
            .in3(N__47520),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47244),
            .ce(N__44417),
            .sr(N__46646));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_12_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_12_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_12_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32471),
            .lcout(\current_shift_inst.un4_control_input_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_12_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_12_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_12_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32462),
            .lcout(\current_shift_inst.un4_control_input_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_12_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_12_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_12_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_12_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32453),
            .lcout(\current_shift_inst.un4_control_input_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_12_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_12_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_12_13_2 .LUT_INIT=16'b0100010001010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_16_LC_12_13_2  (
            .in0(N__44061),
            .in1(N__40453),
            .in2(_gnd_net_),
            .in3(N__43887),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47237),
            .ce(N__31228),
            .sr(N__46655));
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_12_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_12_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_12_13_3 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_17_LC_12_13_3  (
            .in0(N__43888),
            .in1(N__44062),
            .in2(_gnd_net_),
            .in3(N__42346),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47237),
            .ce(N__31228),
            .sr(N__46655));
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_12_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_12_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_12_13_5 .LUT_INIT=16'b0001000100110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_19_LC_12_13_5  (
            .in0(N__41887),
            .in1(N__44060),
            .in2(_gnd_net_),
            .in3(N__40389),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47237),
            .ce(N__31228),
            .sr(N__46655));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_12_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_12_13_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_12_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32486),
            .lcout(\current_shift_inst.un4_control_input_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_12_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_12_13_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_12_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32480),
            .lcout(\current_shift_inst.un4_control_input_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.stoper_state_1_LC_12_14_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.stoper_state_1_LC_12_14_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_slave.stoper_hc.stoper_state_1_LC_12_14_0 .LUT_INIT=16'b0010000001100100;
    LogicCell40 \phase_controller_slave.stoper_hc.stoper_state_1_LC_12_14_0  (
            .in0(N__40981),
            .in1(N__40655),
            .in2(N__40916),
            .in3(N__40739),
            .lcout(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47229),
            .ce(N__40514),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.stoper_state_0_LC_12_14_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.stoper_state_0_LC_12_14_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_slave.stoper_tr.stoper_state_0_LC_12_14_1 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \phase_controller_slave.stoper_tr.stoper_state_0_LC_12_14_1  (
            .in0(N__37793),
            .in1(N__38103),
            .in2(N__38051),
            .in3(N__34417),
            .lcout(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47229),
            .ce(N__40514),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.stoper_state_1_LC_12_14_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.stoper_state_1_LC_12_14_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_slave.stoper_tr.stoper_state_1_LC_12_14_2 .LUT_INIT=16'b0000110001010000;
    LogicCell40 \phase_controller_slave.stoper_tr.stoper_state_1_LC_12_14_2  (
            .in0(N__34418),
            .in1(N__38039),
            .in2(N__38144),
            .in3(N__37794),
            .lcout(\phase_controller_slave.stoper_tr.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47229),
            .ce(N__40514),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.tr_state_0_LC_12_14_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.tr_state_0_LC_12_14_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.tr_state_0_LC_12_14_4 .LUT_INIT=16'b1100110001100110;
    LogicCell40 \delay_measurement_inst.tr_state_0_LC_12_14_4  (
            .in0(N__34910),
            .in1(N__33826),
            .in2(_gnd_net_),
            .in3(N__33812),
            .lcout(\delay_measurement_inst.tr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47229),
            .ce(N__40514),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.hc_state_0_LC_12_14_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.hc_state_0_LC_12_14_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.hc_state_0_LC_12_14_5 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \delay_measurement_inst.hc_state_0_LC_12_14_5  (
            .in0(N__35881),
            .in1(N__35916),
            .in2(_gnd_net_),
            .in3(N__41939),
            .lcout(\delay_measurement_inst.hc_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47229),
            .ce(N__40514),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_12_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_12_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_12_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_12_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31334),
            .lcout(\current_shift_inst.un4_control_input_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_12_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_12_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_12_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31322),
            .lcout(\current_shift_inst.un4_control_input_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_12_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_12_15_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_12_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32621),
            .lcout(\current_shift_inst.un4_control_input_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_12_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_12_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_12_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32555),
            .lcout(\current_shift_inst.un4_control_input_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_12_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_12_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_12_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32585),
            .lcout(\current_shift_inst.un4_control_input_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_12_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_12_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_12_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32660),
            .lcout(\current_shift_inst.un4_control_input_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_12_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_12_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_12_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32597),
            .lcout(\current_shift_inst.un4_control_input_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_12_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_12_15_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_12_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32576),
            .lcout(\current_shift_inst.un4_control_input_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_12_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_12_15_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_12_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32564),
            .lcout(\current_shift_inst.un4_control_input_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_12_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_12_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_12_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32669),
            .lcout(\current_shift_inst.un4_control_input_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_12_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_12_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_12_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32759),
            .lcout(\current_shift_inst.un4_control_input_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_12_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_12_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_12_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32633),
            .lcout(\current_shift_inst.un4_control_input_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_12_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_12_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_12_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32786),
            .lcout(\current_shift_inst.un4_control_input_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_12_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_12_16_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_12_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32777),
            .lcout(\current_shift_inst.un4_control_input_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_12_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_12_16_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_12_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32750),
            .lcout(\current_shift_inst.un4_control_input_axb_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_12_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_12_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_12_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32642),
            .lcout(\current_shift_inst.un4_control_input_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_12_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_12_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_12_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32612),
            .lcout(\current_shift_inst.un4_control_input_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_12_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_12_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_12_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_12_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32651),
            .lcout(\current_shift_inst.un4_control_input_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_LC_12_17_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_LC_12_17_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_LC_12_17_0  (
            .in0(N__32426),
            .in1(N__40393),
            .in2(_gnd_net_),
            .in3(N__41886),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlt31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_z_i_31_LC_12_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_z_i_31_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_z_i_31_LC_12_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_z_i_31_LC_12_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31436),
            .lcout(\current_shift_inst.z_i_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_12_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_12_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_12_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32768),
            .lcout(\current_shift_inst.un4_control_input_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam reset_ibuf_gb_io_RNI79U7_LC_12_17_6.C_ON=1'b0;
    defparam reset_ibuf_gb_io_RNI79U7_LC_12_17_6.SEQ_MODE=4'b0000;
    defparam reset_ibuf_gb_io_RNI79U7_LC_12_17_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 reset_ibuf_gb_io_RNI79U7_LC_12_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46777),
            .lcout(red_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1C4K_24_LC_12_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1C4K_24_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1C4K_24_LC_12_18_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1C4K_24_LC_12_18_0  (
            .in0(N__31502),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31627),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI1C4K_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIB4C81_25_LC_12_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIB4C81_25_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIB4C81_25_LC_12_18_1 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIB4C81_25_LC_12_18_1  (
            .in0(N__31751),
            .in1(N__31783),
            .in2(N__31871),
            .in3(N__31823),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIB4C81_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4G5K_25_LC_12_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4G5K_25_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4G5K_25_LC_12_18_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4G5K_25_LC_12_18_2  (
            .in0(N__31782),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31750),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI4G5K_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7OAK_29_LC_12_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7OAK_29_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7OAK_29_LC_12_18_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7OAK_29_LC_12_18_3  (
            .in0(_gnd_net_),
            .in1(N__31712),
            .in2(_gnd_net_),
            .in3(N__31675),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI7OAK_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVJ781_23_LC_12_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVJ781_23_LC_12_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVJ781_23_LC_12_18_5 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVJ781_23_LC_12_18_5  (
            .in0(N__31626),
            .in1(N__31587),
            .in2(N__31556),
            .in3(N__31503),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIVJ781_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.S3_sync0_LC_12_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.S3_sync0_LC_12_18_6 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.S3_sync0_LC_12_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.S3_sync0_LC_12_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31903),
            .lcout(\current_shift_inst.S3_syncZ0Z0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47212),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_LC_12_19_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_LC_12_19_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_LC_12_19_0  (
            .in0(N__47443),
            .in1(N__34223),
            .in2(N__31931),
            .in3(N__47401),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.target_time_2_LC_12_19_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_2_LC_12_19_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_2_LC_12_19_1 .LUT_INIT=16'b1000110000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_2_LC_12_19_1  (
            .in0(N__40217),
            .in1(N__40094),
            .in2(N__31469),
            .in3(N__37465),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47209),
            .ce(N__44449),
            .sr(N__46707));
    defparam \phase_controller_slave.stoper_tr.target_time_3_LC_12_19_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_3_LC_12_19_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_3_LC_12_19_2 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_3_LC_12_19_2  (
            .in0(N__37466),
            .in1(N__40216),
            .in2(_gnd_net_),
            .in3(N__37422),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47209),
            .ce(N__44449),
            .sr(N__46707));
    defparam \phase_controller_slave.stoper_tr.target_time_1_LC_12_19_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_1_LC_12_19_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_1_LC_12_19_3 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_1_LC_12_19_3  (
            .in0(N__37423),
            .in1(N__37046),
            .in2(N__40121),
            .in3(N__37464),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47209),
            .ce(N__44449),
            .sr(N__46707));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1_6_LC_12_19_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1_6_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1_6_LC_12_19_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1_6_LC_12_19_5  (
            .in0(N__37224),
            .in1(N__37326),
            .in2(_gnd_net_),
            .in3(N__40248),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1Z0Z_6 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0_6_LC_12_19_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0_6_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0_6_LC_12_19_6 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0_6_LC_12_19_6  (
            .in0(_gnd_net_),
            .in1(N__47537),
            .in2(N__31922),
            .in3(N__47400),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.target_time_5_LC_12_19_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_5_LC_12_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_5_LC_12_19_7 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_5_LC_12_19_7  (
            .in0(N__40178),
            .in1(N__41490),
            .in2(N__31919),
            .in3(N__37260),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47209),
            .ce(N__44449),
            .sr(N__46707));
    defparam \phase_controller_slave.start_timer_hc_RNO_1_LC_12_21_0 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_hc_RNO_1_LC_12_21_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.start_timer_hc_RNO_1_LC_12_21_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_slave.start_timer_hc_RNO_1_LC_12_21_0  (
            .in0(N__32150),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32166),
            .lcout(),
            .ltout(\phase_controller_slave.start_timer_hc_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.start_timer_hc_LC_12_21_1 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_hc_LC_12_21_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.start_timer_hc_LC_12_21_1 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \phase_controller_slave.start_timer_hc_LC_12_21_1  (
            .in0(N__33288),
            .in1(N__40802),
            .in2(N__31916),
            .in3(N__47615),
            .lcout(\phase_controller_slave.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47200),
            .ce(),
            .sr(N__46716));
    defparam \phase_controller_slave.state_2_LC_12_21_3 .C_ON=1'b0;
    defparam \phase_controller_slave.state_2_LC_12_21_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.state_2_LC_12_21_3 .LUT_INIT=16'b1011101000110000;
    LogicCell40 \phase_controller_slave.state_2_LC_12_21_3  (
            .in0(N__32167),
            .in1(N__47664),
            .in2(N__47641),
            .in3(N__32151),
            .lcout(\phase_controller_slave.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47200),
            .ce(),
            .sr(N__46716));
    defparam \phase_controller_slave.stoper_hc.time_passed_LC_12_21_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.time_passed_LC_12_21_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.time_passed_LC_12_21_6 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_slave.stoper_hc.time_passed_LC_12_21_6  (
            .in0(N__47663),
            .in1(N__37076),
            .in2(N__34187),
            .in3(N__40738),
            .lcout(\phase_controller_slave.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47200),
            .ce(),
            .sr(N__46716));
    defparam \phase_controller_slave.S1_LC_12_22_0 .C_ON=1'b0;
    defparam \phase_controller_slave.S1_LC_12_22_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.S1_LC_12_22_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_slave.S1_LC_12_22_0  (
            .in0(N__32153),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(s3_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47198),
            .ce(),
            .sr(N__46723));
    defparam \phase_controller_slave.state_0_LC_12_22_2 .C_ON=1'b0;
    defparam \phase_controller_slave.state_0_LC_12_22_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.state_0_LC_12_22_2 .LUT_INIT=16'b1100111000001010;
    LogicCell40 \phase_controller_slave.state_0_LC_12_22_2  (
            .in0(N__33304),
            .in1(N__32246),
            .in2(N__33248),
            .in3(N__32219),
            .lcout(\phase_controller_slave.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47198),
            .ce(),
            .sr(N__46723));
    defparam \phase_controller_slave.state_4_LC_12_22_6 .C_ON=1'b0;
    defparam \phase_controller_slave.state_4_LC_12_22_6 .SEQ_MODE=4'b1011;
    defparam \phase_controller_slave.state_4_LC_12_22_6 .LUT_INIT=16'b1000100011111000;
    LogicCell40 \phase_controller_slave.state_4_LC_12_22_6  (
            .in0(N__33305),
            .in1(N__33247),
            .in2(N__33290),
            .in3(N__34453),
            .lcout(\phase_controller_slave.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47198),
            .ce(),
            .sr(N__46723));
    defparam \phase_controller_slave.state_3_LC_12_22_7 .C_ON=1'b0;
    defparam \phase_controller_slave.state_3_LC_12_22_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.state_3_LC_12_22_7 .LUT_INIT=16'b1010101000001100;
    LogicCell40 \phase_controller_slave.state_3_LC_12_22_7  (
            .in0(N__34454),
            .in1(N__32152),
            .in2(N__32171),
            .in3(N__33287),
            .lcout(\phase_controller_slave.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47198),
            .ce(),
            .sr(N__46723));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_16_LC_12_24_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_16_LC_12_24_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_16_LC_12_24_1 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_16_LC_12_24_1  (
            .in0(N__41027),
            .in1(N__40853),
            .in2(N__40691),
            .in3(N__33374),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47194),
            .ce(),
            .sr(N__46730));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_14_LC_12_24_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_14_LC_12_24_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_14_LC_12_24_6 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_14_LC_12_24_6  (
            .in0(N__40683),
            .in1(N__41028),
            .in2(N__40899),
            .in3(N__33386),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47194),
            .ce(),
            .sr(N__46730));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_12_LC_12_24_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_12_LC_12_24_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_12_LC_12_24_7 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_12_LC_12_24_7  (
            .in0(N__41026),
            .in1(N__40852),
            .in2(N__40690),
            .in3(N__33398),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47194),
            .ce(),
            .sr(N__46730));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_19_LC_12_25_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_19_LC_12_25_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_19_LC_12_25_5 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_19_LC_12_25_5  (
            .in0(N__41058),
            .in1(N__40682),
            .in2(N__40918),
            .in3(N__33356),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47191),
            .ce(),
            .sr(N__46734));
    defparam \current_shift_inst.timer_phase.running_RNIL91O_LC_12_26_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.running_RNIL91O_LC_12_26_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.running_RNIL91O_LC_12_26_1 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \current_shift_inst.timer_phase.running_RNIL91O_LC_12_26_1  (
            .in0(N__33491),
            .in1(N__33541),
            .in2(_gnd_net_),
            .in3(N__33514),
            .lcout(\current_shift_inst.timer_phase.N_192_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.running_RNIB31B_LC_12_26_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.running_RNIB31B_LC_12_26_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.running_RNIB31B_LC_12_26_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_phase.running_RNIB31B_LC_12_26_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33513),
            .lcout(\current_shift_inst.timer_phase.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_12_30_6.C_ON=1'b0;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_12_30_6.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_12_30_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_12_30_6 (
            .in0(N__31955),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_clk_12mhz_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_13_5_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_13_5_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_13_5_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_13_5_1  (
            .in0(_gnd_net_),
            .in1(N__33426),
            .in2(_gnd_net_),
            .in3(N__33585),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_321_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_13_LC_13_6_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_13_LC_13_6_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_13_LC_13_6_4 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_13_LC_13_6_4  (
            .in0(N__34960),
            .in1(N__42551),
            .in2(N__44260),
            .in3(N__42461),
            .lcout(measured_delay_hc_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47310),
            .ce(),
            .sr(N__46604));
    defparam \current_shift_inst.meas_state_0_LC_13_7_0 .C_ON=1'b0;
    defparam \current_shift_inst.meas_state_0_LC_13_7_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.meas_state_0_LC_13_7_0 .LUT_INIT=16'b0111111110101010;
    LogicCell40 \current_shift_inst.meas_state_0_LC_13_7_0  (
            .in0(N__32701),
            .in1(N__32385),
            .in2(N__32357),
            .in3(N__32305),
            .lcout(\current_shift_inst.meas_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47298),
            .ce(),
            .sr(N__46609));
    defparam \current_shift_inst.phase_valid_LC_13_7_1 .C_ON=1'b0;
    defparam \current_shift_inst.phase_valid_LC_13_7_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.phase_valid_LC_13_7_1 .LUT_INIT=16'b1010100011111000;
    LogicCell40 \current_shift_inst.phase_valid_LC_13_7_1  (
            .in0(N__32304),
            .in1(N__32843),
            .in2(N__32392),
            .in3(N__32702),
            .lcout(\current_shift_inst.phase_validZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47298),
            .ce(),
            .sr(N__46609));
    defparam \current_shift_inst.timer_s1.running_LC_13_7_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_LC_13_7_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.running_LC_13_7_2 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \current_shift_inst.timer_s1.running_LC_13_7_2  (
            .in0(N__32352),
            .in1(N__32330),
            .in2(_gnd_net_),
            .in3(N__35569),
            .lcout(\current_shift_inst.timer_s1.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47298),
            .ce(),
            .sr(N__46609));
    defparam \delay_measurement_inst.delay_hc_reg_1_LC_13_7_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_1_LC_13_7_4 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_hc_reg_1_LC_13_7_4 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_1_LC_13_7_4  (
            .in0(N__42526),
            .in1(N__34865),
            .in2(N__41252),
            .in3(N__42099),
            .lcout(measured_delay_hc_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47298),
            .ce(),
            .sr(N__46609));
    defparam \delay_measurement_inst.delay_hc_reg_31_LC_13_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_31_LC_13_7_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_31_LC_13_7_5 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_31_LC_13_7_5  (
            .in0(N__42101),
            .in1(N__44017),
            .in2(_gnd_net_),
            .in3(N__42525),
            .lcout(measured_delay_hc_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47298),
            .ce(),
            .sr(N__46609));
    defparam \delay_measurement_inst.delay_hc_reg_2_LC_13_7_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_2_LC_13_7_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_2_LC_13_7_6 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_2_LC_13_7_6  (
            .in0(N__42527),
            .in1(N__34847),
            .in2(N__34106),
            .in3(N__42100),
            .lcout(measured_delay_hc_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47298),
            .ce(),
            .sr(N__46609));
    defparam \current_shift_inst.stop_timer_s1_RNO_0_LC_13_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.stop_timer_s1_RNO_0_LC_13_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.stop_timer_s1_RNO_0_LC_13_8_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.stop_timer_s1_RNO_0_LC_13_8_0  (
            .in0(N__32380),
            .in1(N__32300),
            .in2(N__32356),
            .in3(N__32696),
            .lcout(),
            .ltout(\current_shift_inst.N_199_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.stop_timer_s1_LC_13_8_1 .C_ON=1'b0;
    defparam \current_shift_inst.stop_timer_s1_LC_13_8_1 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.stop_timer_s1_LC_13_8_1 .LUT_INIT=16'b1111110111110000;
    LogicCell40 \current_shift_inst.stop_timer_s1_LC_13_8_1  (
            .in0(N__32700),
            .in1(N__32308),
            .in2(N__32258),
            .in3(N__32329),
            .lcout(\current_shift_inst.stop_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47289),
            .ce(N__40522),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_8_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_8_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_8_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.timer_s1.running_RNII51H_LC_13_8_2  (
            .in0(_gnd_net_),
            .in1(N__35558),
            .in2(_gnd_net_),
            .in3(N__32327),
            .lcout(\current_shift_inst.timer_s1.N_187_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.start_timer_s1_LC_13_8_3 .C_ON=1'b0;
    defparam \current_shift_inst.start_timer_s1_LC_13_8_3 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.start_timer_s1_LC_13_8_3 .LUT_INIT=16'b0111111100001010;
    LogicCell40 \current_shift_inst.start_timer_s1_LC_13_8_3  (
            .in0(N__32698),
            .in1(N__32381),
            .in2(N__32309),
            .in3(N__32351),
            .lcout(\current_shift_inst.start_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47289),
            .ce(N__40522),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_8_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_8_4 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_8_4  (
            .in0(N__32350),
            .in1(N__35559),
            .in2(_gnd_net_),
            .in3(N__32328),
            .lcout(\current_shift_inst.timer_s1.N_191_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.start_timer_phase_LC_13_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.start_timer_phase_LC_13_8_5 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.start_timer_phase_LC_13_8_5 .LUT_INIT=16'b0011111100100010;
    LogicCell40 \current_shift_inst.start_timer_phase_LC_13_8_5  (
            .in0(N__32697),
            .in1(N__32307),
            .in2(N__32842),
            .in3(N__33529),
            .lcout(\current_shift_inst.start_timer_phaseZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47289),
            .ce(N__40522),
            .sr(_gnd_net_));
    defparam \current_shift_inst.stop_timer_phase_LC_13_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.stop_timer_phase_LC_13_8_6 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.stop_timer_phase_LC_13_8_6 .LUT_INIT=16'b1011101010110000;
    LogicCell40 \current_shift_inst.stop_timer_phase_LC_13_8_6  (
            .in0(N__32306),
            .in1(N__32699),
            .in2(N__33482),
            .in3(N__32838),
            .lcout(\current_shift_inst.stop_timer_phaseZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47289),
            .ce(N__40522),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.stop_timer_hc_LC_13_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_hc_LC_13_9_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.stop_timer_hc_LC_13_9_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \delay_measurement_inst.stop_timer_hc_LC_13_9_0  (
            .in0(N__41930),
            .in1(N__35882),
            .in2(N__46781),
            .in3(N__35930),
            .lcout(\delay_measurement_inst.stop_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47282),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_13_LC_13_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_13_LC_13_9_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_13_LC_13_9_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_13_LC_13_9_3  (
            .in0(N__35080),
            .in1(N__35128),
            .in2(N__34961),
            .in3(N__35206),
            .lcout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto5_3_LC_13_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto5_3_LC_13_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto5_3_LC_13_9_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto5_3_LC_13_9_6  (
            .in0(N__34099),
            .in1(N__41248),
            .in2(N__35517),
            .in3(N__42243),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un1_startlto5Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto6_LC_13_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto6_LC_13_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto6_LC_13_9_7 .LUT_INIT=16'b1100110010001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto6_LC_13_9_7  (
            .in0(N__43954),
            .in1(N__34151),
            .in2(N__32276),
            .in3(N__35426),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlt8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto9_0_0_LC_13_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto9_0_0_LC_13_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto9_0_0_LC_13_10_4 .LUT_INIT=16'b1011000000110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto9_0_0_LC_13_10_4  (
            .in0(N__34030),
            .in1(N__33719),
            .in2(N__33876),
            .in3(N__32444),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlt15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_9_LC_13_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_9_LC_13_10_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_9_LC_13_10_5 .LUT_INIT=16'b1011100011111111;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_9_LC_13_10_5  (
            .in0(N__35081),
            .in1(N__42624),
            .in2(N__34046),
            .in3(N__42092),
            .lcout(measured_delay_hc_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47274),
            .ce(),
            .sr(N__46628));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_8_LC_13_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_8_LC_13_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_8_LC_13_11_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_8_LC_13_11_0  (
            .in0(N__44274),
            .in1(N__33901),
            .in2(N__40439),
            .in3(N__33853),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_13_LC_13_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_13_LC_13_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_13_LC_13_11_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_13_LC_13_11_1  (
            .in0(N__35633),
            .in1(N__39302),
            .in2(N__32438),
            .in3(N__32435),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_5_LC_13_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_5_LC_13_11_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_5_LC_13_11_4 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_5_LC_13_11_4  (
            .in0(N__42628),
            .in1(N__34814),
            .in2(N__43958),
            .in3(N__42421),
            .lcout(measured_delay_hc_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47263),
            .ce(),
            .sr(N__46634));
    defparam \delay_measurement_inst.delay_hc_reg_14_LC_13_11_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_14_LC_13_11_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_14_LC_13_11_5 .LUT_INIT=16'b1110111011111010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_14_LC_13_11_5  (
            .in0(N__42418),
            .in1(N__35303),
            .in2(N__33866),
            .in3(N__42625),
            .lcout(measured_delay_hc_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47263),
            .ce(),
            .sr(N__46634));
    defparam \delay_measurement_inst.delay_hc_reg_15_LC_13_11_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_15_LC_13_11_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_15_LC_13_11_6 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_15_LC_13_11_6  (
            .in0(N__42626),
            .in1(N__33902),
            .in2(N__35267),
            .in3(N__42419),
            .lcout(measured_delay_hc_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47263),
            .ce(),
            .sr(N__46634));
    defparam \delay_measurement_inst.delay_hc_reg_16_LC_13_11_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_16_LC_13_11_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_16_LC_13_11_7 .LUT_INIT=16'b1111101111101010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_16_LC_13_11_7  (
            .in0(N__42420),
            .in1(N__42627),
            .in2(N__35210),
            .in3(N__40429),
            .lcout(measured_delay_hc_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47263),
            .ce(),
            .sr(N__46634));
    defparam \phase_controller_inst1.state_RNIR0JF_1_LC_13_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNIR0JF_1_LC_13_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNIR0JF_1_LC_13_12_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.state_RNIR0JF_1_LC_13_12_1  (
            .in0(_gnd_net_),
            .in1(N__43077),
            .in2(_gnd_net_),
            .in3(N__43033),
            .lcout(\phase_controller_inst1.T01_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_RNO_0_3_LC_13_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNO_0_3_LC_13_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNO_0_3_LC_13_12_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.state_RNO_0_3_LC_13_12_2  (
            .in0(N__34545),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43150),
            .lcout(),
            .ltout(\phase_controller_inst1.N_86_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_3_LC_13_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_3_LC_13_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_3_LC_13_12_3 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \phase_controller_inst1.state_3_LC_13_12_3  (
            .in0(N__32507),
            .in1(N__32543),
            .in2(N__32510),
            .in3(N__43175),
            .lcout(\phase_controller_inst1.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47254),
            .ce(),
            .sr(N__46640));
    defparam \phase_controller_inst1.state_4_LC_13_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_4_LC_13_12_5 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst1.state_4_LC_13_12_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \phase_controller_inst1.state_4_LC_13_12_5  (
            .in0(N__43151),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34544),
            .lcout(\phase_controller_inst1.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47254),
            .ce(),
            .sr(N__46640));
    defparam \phase_controller_inst1.S1_LC_13_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.S1_LC_13_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S1_LC_13_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S1_LC_13_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32506),
            .lcout(s1_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47254),
            .ce(),
            .sr(N__46640));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_13_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_13_13_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_13_13_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_13_13_0  (
            .in0(_gnd_net_),
            .in1(N__35797),
            .in2(N__35855),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_3 ),
            .ltout(),
            .carryin(bfn_13_13_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .clk(N__47246),
            .ce(N__32741),
            .sr(N__46647));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_13_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_13_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_13_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_13_13_1  (
            .in0(_gnd_net_),
            .in1(N__35776),
            .in2(N__35828),
            .in3(N__32474),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .clk(N__47246),
            .ce(N__32741),
            .sr(N__46647));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_13_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_13_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_13_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_13_13_2  (
            .in0(_gnd_net_),
            .in1(N__35798),
            .in2(N__35755),
            .in3(N__32465),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .clk(N__47246),
            .ce(N__32741),
            .sr(N__46647));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_13_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_13_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_13_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_13_13_3  (
            .in0(_gnd_net_),
            .in1(N__35777),
            .in2(N__35725),
            .in3(N__32456),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .clk(N__47246),
            .ce(N__32741),
            .sr(N__46647));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_13_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_13_13_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_13_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_13_13_4  (
            .in0(_gnd_net_),
            .in1(N__36130),
            .in2(N__35756),
            .in3(N__32447),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .clk(N__47246),
            .ce(N__32741),
            .sr(N__46647));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_13_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_13_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_13_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_13_13_5  (
            .in0(_gnd_net_),
            .in1(N__36109),
            .in2(N__35726),
            .in3(N__32603),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .clk(N__47246),
            .ce(N__32741),
            .sr(N__46647));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_13_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_13_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_13_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_13_13_6  (
            .in0(_gnd_net_),
            .in1(N__36131),
            .in2(N__36089),
            .in3(N__32600),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .clk(N__47246),
            .ce(N__32741),
            .sr(N__46647));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_13_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_13_13_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_13_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_13_13_7  (
            .in0(_gnd_net_),
            .in1(N__36110),
            .in2(N__36056),
            .in3(N__32588),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .clk(N__47246),
            .ce(N__32741),
            .sr(N__46647));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_13_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_13_14_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_13_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_13_14_0  (
            .in0(_gnd_net_),
            .in1(N__36082),
            .in2(N__36025),
            .in3(N__32579),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_11 ),
            .ltout(),
            .carryin(bfn_13_14_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .clk(N__47238),
            .ce(N__32740),
            .sr(N__46656));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_13_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_13_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_13_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_13_14_1  (
            .in0(_gnd_net_),
            .in1(N__36055),
            .in2(N__35998),
            .in3(N__32570),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .clk(N__47238),
            .ce(N__32740),
            .sr(N__46656));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_13_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_13_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_13_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_13_14_2  (
            .in0(_gnd_net_),
            .in1(N__35971),
            .in2(N__36026),
            .in3(N__32567),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .clk(N__47238),
            .ce(N__32740),
            .sr(N__46656));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_13_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_13_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_13_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_13_14_3  (
            .in0(_gnd_net_),
            .in1(N__35950),
            .in2(N__35999),
            .in3(N__32558),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .clk(N__47238),
            .ce(N__32740),
            .sr(N__46656));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_13_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_13_14_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_13_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_13_14_4  (
            .in0(_gnd_net_),
            .in1(N__35972),
            .in2(N__36364),
            .in3(N__32549),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .clk(N__47238),
            .ce(N__32740),
            .sr(N__46656));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_13_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_13_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_13_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_13_14_5  (
            .in0(_gnd_net_),
            .in1(N__35951),
            .in2(N__36337),
            .in3(N__32546),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .clk(N__47238),
            .ce(N__32740),
            .sr(N__46656));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_13_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_13_14_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_13_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_13_14_6  (
            .in0(_gnd_net_),
            .in1(N__36310),
            .in2(N__36365),
            .in3(N__32672),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .clk(N__47238),
            .ce(N__32740),
            .sr(N__46656));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_13_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_13_14_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_13_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_13_14_7  (
            .in0(_gnd_net_),
            .in1(N__36281),
            .in2(N__36338),
            .in3(N__32663),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .clk(N__47238),
            .ce(N__32740),
            .sr(N__46656));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_13_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_13_15_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_13_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_13_15_0  (
            .in0(_gnd_net_),
            .in1(N__36311),
            .in2(N__36253),
            .in3(N__32654),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_19 ),
            .ltout(),
            .carryin(bfn_13_15_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .clk(N__47230),
            .ce(N__32739),
            .sr(N__46665));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_13_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_13_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_13_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_13_15_1  (
            .in0(_gnd_net_),
            .in1(N__36280),
            .in2(N__36226),
            .in3(N__32645),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .clk(N__47230),
            .ce(N__32739),
            .sr(N__46665));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_13_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_13_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_13_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_13_15_2  (
            .in0(_gnd_net_),
            .in1(N__36199),
            .in2(N__36254),
            .in3(N__32636),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .clk(N__47230),
            .ce(N__32739),
            .sr(N__46665));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_13_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_13_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_13_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_13_15_3  (
            .in0(_gnd_net_),
            .in1(N__36178),
            .in2(N__36227),
            .in3(N__32627),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .clk(N__47230),
            .ce(N__32739),
            .sr(N__46665));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_13_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_13_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_13_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_13_15_4  (
            .in0(_gnd_net_),
            .in1(N__36200),
            .in2(N__36157),
            .in3(N__32624),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .clk(N__47230),
            .ce(N__32739),
            .sr(N__46665));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_13_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_13_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_13_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_13_15_5  (
            .in0(_gnd_net_),
            .in1(N__36179),
            .in2(N__36700),
            .in3(N__32615),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .clk(N__47230),
            .ce(N__32739),
            .sr(N__46665));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_13_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_13_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_13_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_13_15_6  (
            .in0(_gnd_net_),
            .in1(N__36674),
            .in2(N__36158),
            .in3(N__32606),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .clk(N__47230),
            .ce(N__32739),
            .sr(N__46665));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_13_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_13_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_13_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_13_15_7  (
            .in0(_gnd_net_),
            .in1(N__36647),
            .in2(N__36701),
            .in3(N__32780),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .clk(N__47230),
            .ce(N__32739),
            .sr(N__46665));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_13_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_13_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_13_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_13_16_0  (
            .in0(_gnd_net_),
            .in1(N__36673),
            .in2(N__36619),
            .in3(N__32771),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_27 ),
            .ltout(),
            .carryin(bfn_13_16_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .clk(N__47225),
            .ce(N__32737),
            .sr(N__46675));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_13_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_13_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_13_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_13_16_1  (
            .in0(_gnd_net_),
            .in1(N__36646),
            .in2(N__36592),
            .in3(N__32762),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .clk(N__47225),
            .ce(N__32737),
            .sr(N__46675));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_13_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_13_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_13_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_13_16_2  (
            .in0(_gnd_net_),
            .in1(N__36566),
            .in2(N__36620),
            .in3(N__32753),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .clk(N__47225),
            .ce(N__32737),
            .sr(N__46675));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_13_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_13_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_13_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_13_16_3  (
            .in0(_gnd_net_),
            .in1(N__36425),
            .in2(N__36593),
            .in3(N__32744),
            .lcout(\current_shift_inst.timer_s1.elapsed_time_ns_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ),
            .clk(N__47225),
            .ce(N__32737),
            .sr(N__46675));
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_13_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_13_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_13_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_13_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32720),
            .lcout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.S1_rise_LC_13_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.S1_rise_LC_13_17_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.S1_rise_LC_13_17_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \current_shift_inst.S1_rise_LC_13_17_0  (
            .in0(_gnd_net_),
            .in1(N__32807),
            .in2(_gnd_net_),
            .in3(N__32815),
            .lcout(\current_shift_inst.S1_riseZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47222),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.S3_sync_prev_LC_13_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.S3_sync_prev_LC_13_17_1 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.S3_sync_prev_LC_13_17_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.S3_sync_prev_LC_13_17_1  (
            .in0(N__32795),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.S3_sync_prevZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47222),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.S1_sync0_LC_13_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.S1_sync0_LC_13_17_2 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.S1_sync0_LC_13_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.S1_sync0_LC_13_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32875),
            .lcout(\current_shift_inst.S1_syncZ0Z0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47222),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.S1_sync1_LC_13_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.S1_sync1_LC_13_17_3 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.S1_sync1_LC_13_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.S1_sync1_LC_13_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32855),
            .lcout(\current_shift_inst.S1_syncZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47222),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.S3_rise_LC_13_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.S3_rise_LC_13_17_4 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.S3_rise_LC_13_17_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \current_shift_inst.S3_rise_LC_13_17_4  (
            .in0(_gnd_net_),
            .in1(N__32849),
            .in2(_gnd_net_),
            .in3(N__32794),
            .lcout(\current_shift_inst.S3_riseZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47222),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.S1_sync_prev_LC_13_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.S1_sync_prev_LC_13_17_5 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.S1_sync_prev_LC_13_17_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.S1_sync_prev_LC_13_17_5  (
            .in0(N__32816),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.S1_sync_prevZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47222),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.S3_sync1_LC_13_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.S3_sync1_LC_13_17_7 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.S3_sync1_LC_13_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.S3_sync1_LC_13_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32801),
            .lcout(\current_shift_inst.S3_syncZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47222),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.target_time_6_LC_13_18_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_6_LC_13_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_6_LC_13_18_0 .LUT_INIT=16'b0100010001000101;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_6_LC_13_18_0  (
            .in0(N__37350),
            .in1(N__40249),
            .in2(N__41492),
            .in3(N__37256),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47216),
            .ce(N__44444),
            .sr(N__46688));
    defparam \phase_controller_slave.stoper_tr.target_time_4_LC_13_18_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_4_LC_13_18_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_4_LC_13_18_1 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_4_LC_13_18_1  (
            .in0(N__37255),
            .in1(N__41485),
            .in2(N__43501),
            .in3(N__37349),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47216),
            .ce(N__44444),
            .sr(N__46688));
    defparam \phase_controller_slave.stoper_tr.target_time_7_LC_13_18_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_7_LC_13_18_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_7_LC_13_18_2 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_7_LC_13_18_2  (
            .in0(N__41482),
            .in1(N__37328),
            .in2(_gnd_net_),
            .in3(N__37254),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47216),
            .ce(N__44444),
            .sr(N__46688));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_6_LC_13_18_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_6_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_6_LC_13_18_3 .LUT_INIT=16'b0001010100010001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_6_LC_13_18_3  (
            .in0(N__47534),
            .in1(N__47707),
            .in2(N__47442),
            .in3(N__47390),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.target_time_8_LC_13_18_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_8_LC_13_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_8_LC_13_18_4 .LUT_INIT=16'b1111101000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_8_LC_13_18_4  (
            .in0(N__41483),
            .in1(_gnd_net_),
            .in2(N__32978),
            .in3(N__37226),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47216),
            .ce(N__44444),
            .sr(N__46688));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_13_LC_13_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_13_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_13_LC_13_18_5 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_13_LC_13_18_5  (
            .in0(_gnd_net_),
            .in1(N__41481),
            .in2(_gnd_net_),
            .in3(N__47831),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.target_time_9_LC_13_18_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_9_LC_13_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_9_LC_13_18_6 .LUT_INIT=16'b1100111111001101;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_9_LC_13_18_6  (
            .in0(N__47391),
            .in1(N__47435),
            .in2(N__32975),
            .in3(N__47536),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47216),
            .ce(N__44444),
            .sr(N__46688));
    defparam \phase_controller_slave.stoper_tr.target_time_14_LC_13_18_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_14_LC_13_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_14_LC_13_18_7 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_14_LC_13_18_7  (
            .in0(N__47535),
            .in1(N__41484),
            .in2(_gnd_net_),
            .in3(N__47708),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47216),
            .ce(N__44444),
            .sr(N__46688));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_13_19_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_13_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_13_19_0  (
            .in0(_gnd_net_),
            .in1(N__32960),
            .in2(N__32972),
            .in3(N__34365),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_13_19_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_13_19_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_13_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_13_19_1  (
            .in0(_gnd_net_),
            .in1(N__32945),
            .in2(N__32954),
            .in3(N__34345),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_13_19_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_13_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_13_19_2  (
            .in0(_gnd_net_),
            .in1(N__32930),
            .in2(N__32939),
            .in3(N__34309),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_13_19_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_13_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_13_19_3  (
            .in0(_gnd_net_),
            .in1(N__32912),
            .in2(N__32924),
            .in3(N__34279),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_13_19_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_13_19_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_13_19_4  (
            .in0(_gnd_net_),
            .in1(N__32894),
            .in2(N__32906),
            .in3(N__34249),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_13_19_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_13_19_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_13_19_5  (
            .in0(_gnd_net_),
            .in1(N__33128),
            .in2(N__33137),
            .in3(N__34726),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_13_19_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_13_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_13_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_13_19_6  (
            .in0(_gnd_net_),
            .in1(N__33110),
            .in2(N__33122),
            .in3(N__34699),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_13_19_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_13_19_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_13_19_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_13_19_7  (
            .in0(_gnd_net_),
            .in1(N__33095),
            .in2(N__33104),
            .in3(N__34666),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_13_20_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_13_20_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_13_20_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_13_20_0  (
            .in0(_gnd_net_),
            .in1(N__33077),
            .in2(N__33089),
            .in3(N__37517),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_13_20_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_13_20_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_13_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_13_20_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_13_20_1  (
            .in0(N__34636),
            .in1(N__33056),
            .in2(N__33071),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_13_20_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_13_20_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_13_20_2  (
            .in0(_gnd_net_),
            .in1(N__33032),
            .in2(N__33050),
            .in3(N__34607),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_13_20_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_13_20_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_13_20_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_13_20_3  (
            .in0(_gnd_net_),
            .in1(N__33008),
            .in2(N__33026),
            .in3(N__37655),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_13_20_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_13_20_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_13_20_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_13_20_4  (
            .in0(_gnd_net_),
            .in1(N__32984),
            .in2(N__33002),
            .in3(N__37541),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_13_20_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_13_20_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_13_20_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_13_20_5  (
            .in0(_gnd_net_),
            .in1(N__33203),
            .in2(N__33218),
            .in3(N__38324),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_13_20_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_13_20_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_13_20_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_13_20_6  (
            .in0(_gnd_net_),
            .in1(N__33179),
            .in2(N__33197),
            .in3(N__37679),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_13_20_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_13_20_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_13_20_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_13_20_7  (
            .in0(_gnd_net_),
            .in1(N__33173),
            .in2(N__44471),
            .in3(N__37631),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_13_21_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_13_21_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_13_21_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_13_21_0  (
            .in0(_gnd_net_),
            .in1(N__33167),
            .in2(N__33146),
            .in3(N__38222),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_13_21_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_13_21_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_13_21_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_13_21_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_13_21_1  (
            .in0(_gnd_net_),
            .in1(N__33161),
            .in2(N__33323),
            .in3(N__38198),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_13_21_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_13_21_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_13_21_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_13_21_2  (
            .in0(_gnd_net_),
            .in1(N__33155),
            .in2(N__33314),
            .in3(N__37760),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_13_21_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_13_21_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_13_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_13_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33149),
            .lcout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.target_time_17_LC_13_21_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_17_LC_13_21_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_17_LC_13_21_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_17_LC_13_21_4  (
            .in0(N__43297),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47206),
            .ce(N__44445),
            .sr(N__46711));
    defparam \phase_controller_slave.stoper_tr.target_time_18_LC_13_21_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_18_LC_13_21_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_18_LC_13_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_18_LC_13_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43211),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47206),
            .ce(N__44445),
            .sr(N__46711));
    defparam \phase_controller_slave.stoper_tr.target_time_19_LC_13_21_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_19_LC_13_21_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_19_LC_13_21_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_19_LC_13_21_6  (
            .in0(N__41576),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47206),
            .ce(N__44445),
            .sr(N__46711));
    defparam \phase_controller_slave.start_timer_tr_RNO_0_LC_13_22_0 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_tr_RNO_0_LC_13_22_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.start_timer_tr_RNO_0_LC_13_22_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.start_timer_tr_RNO_0_LC_13_22_0  (
            .in0(_gnd_net_),
            .in1(N__33242),
            .in2(_gnd_net_),
            .in3(N__33303),
            .lcout(),
            .ltout(\phase_controller_slave.N_210_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.start_timer_tr_LC_13_22_1 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_tr_LC_13_22_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.start_timer_tr_LC_13_22_1 .LUT_INIT=16'b1100110111001100;
    LogicCell40 \phase_controller_slave.start_timer_tr_LC_13_22_1  (
            .in0(N__33289),
            .in1(N__33266),
            .in2(N__33254),
            .in3(N__37951),
            .lcout(\phase_controller_slave.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47202),
            .ce(),
            .sr(N__46717));
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNI38A6_0_LC_13_22_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNI38A6_0_LC_13_22_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNI38A6_0_LC_13_22_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.stoper_state_RNI38A6_0_LC_13_22_2  (
            .in0(_gnd_net_),
            .in1(N__37859),
            .in2(_gnd_net_),
            .in3(N__38145),
            .lcout(\phase_controller_slave.stoper_tr.time_passed11 ),
            .ltout(\phase_controller_slave.stoper_tr.time_passed11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.time_passed_LC_13_22_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.time_passed_LC_13_22_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.time_passed_LC_13_22_3 .LUT_INIT=16'b1010100010111000;
    LogicCell40 \phase_controller_slave.stoper_tr.time_passed_LC_13_22_3  (
            .in0(N__33243),
            .in1(N__33224),
            .in2(N__33251),
            .in3(N__34410),
            .lcout(\phase_controller_slave.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47202),
            .ce(),
            .sr(N__46717));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_11_LC_13_22_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_11_LC_13_22_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_11_LC_13_22_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_11_LC_13_22_4  (
            .in0(N__37861),
            .in1(N__38147),
            .in2(N__37998),
            .in3(N__34592),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47202),
            .ce(),
            .sr(N__46717));
    defparam \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_13_22_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_13_22_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_13_22_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_13_22_6  (
            .in0(N__37947),
            .in1(N__37860),
            .in2(_gnd_net_),
            .in3(N__38146),
            .lcout(\phase_controller_slave.stoper_tr.time_passed_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_13_23_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_13_23_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_13_23_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_13_23_0  (
            .in0(_gnd_net_),
            .in1(N__34208),
            .in2(N__38291),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_23_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_13_23_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_13_23_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_13_23_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_13_23_1  (
            .in0(_gnd_net_),
            .in1(N__38252),
            .in2(_gnd_net_),
            .in3(N__33350),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_13_23_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_13_23_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_13_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_13_23_2  (
            .in0(_gnd_net_),
            .in1(N__34577),
            .in2(N__36833),
            .in3(N__33347),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_13_23_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_13_23_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_13_23_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_13_23_3  (
            .in0(_gnd_net_),
            .in1(N__37601),
            .in2(_gnd_net_),
            .in3(N__33344),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_13_23_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_13_23_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_13_23_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_13_23_4  (
            .in0(_gnd_net_),
            .in1(N__37568),
            .in2(_gnd_net_),
            .in3(N__33341),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_13_23_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_13_23_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_13_23_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_13_23_5  (
            .in0(_gnd_net_),
            .in1(N__37487),
            .in2(_gnd_net_),
            .in3(N__33338),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_13_23_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_13_23_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_13_23_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_13_23_6  (
            .in0(_gnd_net_),
            .in1(N__36749),
            .in2(_gnd_net_),
            .in3(N__33335),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_13_23_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_13_23_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_13_23_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_13_23_7  (
            .in0(_gnd_net_),
            .in1(N__36725),
            .in2(_gnd_net_),
            .in3(N__33332),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_13_24_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_13_24_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_13_24_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_13_24_0  (
            .in0(_gnd_net_),
            .in1(N__38509),
            .in2(_gnd_net_),
            .in3(N__33329),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9 ),
            .ltout(),
            .carryin(bfn_13_24_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_13_24_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_13_24_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_13_24_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_13_24_1  (
            .in0(_gnd_net_),
            .in1(N__37733),
            .in2(_gnd_net_),
            .in3(N__33326),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_13_24_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_13_24_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_13_24_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_13_24_2  (
            .in0(_gnd_net_),
            .in1(N__37705),
            .in2(_gnd_net_),
            .in3(N__33401),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_13_24_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_13_24_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_13_24_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_13_24_3  (
            .in0(_gnd_net_),
            .in1(N__36961),
            .in2(_gnd_net_),
            .in3(N__33392),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_13_24_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_13_24_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_13_24_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_13_24_4  (
            .in0(_gnd_net_),
            .in1(N__36934),
            .in2(_gnd_net_),
            .in3(N__33389),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_13_24_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_13_24_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_13_24_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_13_24_5  (
            .in0(_gnd_net_),
            .in1(N__36895),
            .in2(_gnd_net_),
            .in3(N__33380),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_13_24_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_13_24_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_13_24_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_13_24_6  (
            .in0(_gnd_net_),
            .in1(N__38476),
            .in2(_gnd_net_),
            .in3(N__33377),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_13_24_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_13_24_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_13_24_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_13_24_7  (
            .in0(_gnd_net_),
            .in1(N__37174),
            .in2(_gnd_net_),
            .in3(N__33368),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_13_25_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_13_25_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_13_25_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_13_25_0  (
            .in0(_gnd_net_),
            .in1(N__37150),
            .in2(_gnd_net_),
            .in3(N__33365),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17 ),
            .ltout(),
            .carryin(bfn_13_25_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_13_25_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_13_25_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_13_25_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_13_25_1  (
            .in0(_gnd_net_),
            .in1(N__37126),
            .in2(_gnd_net_),
            .in3(N__33362),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_13_25_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_13_25_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_13_25_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_13_25_2  (
            .in0(_gnd_net_),
            .in1(N__37099),
            .in2(_gnd_net_),
            .in3(N__33359),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_phase.running_LC_13_26_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.running_LC_13_26_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_phase.running_LC_13_26_2 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \current_shift_inst.timer_phase.running_LC_13_26_2  (
            .in0(N__33542),
            .in1(N__33515),
            .in2(_gnd_net_),
            .in3(N__33489),
            .lcout(\current_shift_inst.timer_phase.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47192),
            .ce(),
            .sr(N__46735));
    defparam \current_shift_inst.timer_phase.running_RNIC90O_LC_13_27_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_phase.running_RNIC90O_LC_13_27_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_phase.running_RNIC90O_LC_13_27_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.timer_phase.running_RNIC90O_LC_13_27_7  (
            .in0(_gnd_net_),
            .in1(N__33512),
            .in2(_gnd_net_),
            .in3(N__33490),
            .lcout(\current_shift_inst.timer_phase.N_188_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.S2_LC_13_28_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.S2_LC_13_28_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S2_LC_13_28_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S2_LC_13_28_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43100),
            .lcout(s2_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47189),
            .ce(),
            .sr(N__46739));
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_14_5_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_14_5_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_14_5_5 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_LC_14_5_5  (
            .in0(N__35903),
            .in1(N__33431),
            .in2(_gnd_net_),
            .in3(N__33591),
            .lcout(\delay_measurement_inst.delay_hc_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47326),
            .ce(),
            .sr(N__46596));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJG9N1_1_LC_14_6_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJG9N1_1_LC_14_6_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJG9N1_1_LC_14_6_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJG9N1_1_LC_14_6_3  (
            .in0(N__35538),
            .in1(N__34839),
            .in2(N__34813),
            .in3(N__34858),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINGQU3_9_LC_14_6_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINGQU3_9_LC_14_6_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINGQU3_9_LC_14_6_4 .LUT_INIT=16'b0011111100101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINGQU3_9_LC_14_6_4  (
            .in0(N__35075),
            .in1(N__34871),
            .in2(N__33434),
            .in3(N__35259),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_2_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_14_7_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_14_7_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_14_7_0 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_14_7_0  (
            .in0(N__33593),
            .in1(N__35899),
            .in2(_gnd_net_),
            .in3(N__33427),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_322_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOHNN2_6_LC_14_7_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOHNN2_6_LC_14_7_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOHNN2_6_LC_14_7_1 .LUT_INIT=16'b0010101000001010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOHNN2_6_LC_14_7_1  (
            .in0(N__33691),
            .in1(N__35117),
            .in2(N__35076),
            .in3(N__33611),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1LC84_14_LC_14_7_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1LC84_14_LC_14_7_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1LC84_14_LC_14_7_2 .LUT_INIT=16'b1100111000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1LC84_14_LC_14_7_2  (
            .in0(N__35302),
            .in1(N__35257),
            .in2(N__33404),
            .in3(N__33554),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt30_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_14_7_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_14_7_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_14_7_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_14_7_3  (
            .in0(_gnd_net_),
            .in1(N__41792),
            .in2(_gnd_net_),
            .in3(N__41697),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_10_LC_14_7_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_10_LC_14_7_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_10_LC_14_7_4 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_10_LC_14_7_4  (
            .in0(N__33620),
            .in1(N__34823),
            .in2(N__33605),
            .in3(N__33560),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOVQ9D_14_LC_14_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOVQ9D_14_LC_14_7_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOVQ9D_14_LC_14_7_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOVQ9D_14_LC_14_7_5  (
            .in0(N__35597),
            .in1(N__33656),
            .in2(N__33602),
            .in3(N__33599),
            .lcout(\delay_measurement_inst.un1_elapsed_time_hc ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_14_7_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_14_7_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_14_7_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_14_7_6  (
            .in0(N__33592),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI93LG1_14_LC_14_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI93LG1_14_LC_14_8_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI93LG1_14_LC_14_8_0 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI93LG1_14_LC_14_8_0  (
            .in0(N__35249),
            .in1(N__35288),
            .in2(_gnd_net_),
            .in3(N__33553),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI537G_17_LC_14_8_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI537G_17_LC_14_8_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI537G_17_LC_14_8_1 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI537G_17_LC_14_8_1  (
            .in0(N__42205),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42481),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4UNN2_4_LC_14_8_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4UNN2_4_LC_14_8_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4UNN2_4_LC_14_8_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4UNN2_4_LC_14_8_2  (
            .in0(N__33569),
            .in1(N__35449),
            .in2(N__33563),
            .in3(N__34803),
            .lcout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_14_8_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_14_8_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_14_8_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_14_8_3  (
            .in0(N__35002),
            .in1(N__34947),
            .in2(N__34983),
            .in3(N__35031),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_14_8_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_14_8_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_14_8_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_14_8_5  (
            .in0(N__42204),
            .in1(N__42480),
            .in2(N__42129),
            .in3(N__35194),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ0JH1_6_LC_14_8_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ0JH1_6_LC_14_8_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ0JH1_6_LC_14_8_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ0JH1_6_LC_14_8_6  (
            .in0(N__41793),
            .in1(N__41698),
            .in2(N__35124),
            .in3(N__35256),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52G18_14_LC_14_8_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52G18_14_LC_14_8_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52G18_14_LC_14_8_7 .LUT_INIT=16'b0101110100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52G18_14_LC_14_8_7  (
            .in0(N__33692),
            .in1(N__33680),
            .in2(N__33671),
            .in3(N__33668),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP8VO1_20_LC_14_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP8VO1_20_LC_14_9_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP8VO1_20_LC_14_9_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP8VO1_20_LC_14_9_0  (
            .in0(N__35144),
            .in1(N__35156),
            .in2(N__35171),
            .in3(N__33646),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_1 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5483B_31_LC_14_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5483B_31_LC_14_9_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5483B_31_LC_14_9_1 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5483B_31_LC_14_9_1  (
            .in0(N__35593),
            .in1(N__35315),
            .in2(N__33662),
            .in3(N__33629),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto31_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_14_9_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_14_9_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_14_9_4  (
            .in0(_gnd_net_),
            .in1(N__35143),
            .in2(_gnd_net_),
            .in3(N__35155),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINN412_20_LC_14_9_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINN412_20_LC_14_9_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINN412_20_LC_14_9_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINN412_20_LC_14_9_5  (
            .in0(N__33647),
            .in1(N__35313),
            .in2(N__33659),
            .in3(N__35170),
            .lcout(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_14_9_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_14_9_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_14_9_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_14_9_6  (
            .in0(N__35351),
            .in1(N__35360),
            .in2(N__35342),
            .in3(N__35369),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5483B_0_31_LC_14_9_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5483B_0_31_LC_14_9_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5483B_0_31_LC_14_9_7 .LUT_INIT=16'b0011001100010011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5483B_0_31_LC_14_9_7  (
            .in0(N__35592),
            .in1(N__35314),
            .in2(N__33638),
            .in3(N__33628),
            .lcout(\delay_measurement_inst.delay_hc_reg3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOJD01_11_LC_14_10_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOJD01_11_LC_14_10_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOJD01_11_LC_14_10_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOJD01_11_LC_14_10_1  (
            .in0(N__35260),
            .in1(N__34984),
            .in2(N__35012),
            .in3(N__35298),
            .lcout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_10_LC_14_10_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_10_LC_14_10_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_10_LC_14_10_2 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_10_LC_14_10_2  (
            .in0(N__42621),
            .in1(N__35039),
            .in2(N__35677),
            .in3(N__42378),
            .lcout(measured_delay_hc_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47283),
            .ce(),
            .sr(N__46618));
    defparam \delay_measurement_inst.delay_hc_reg_11_LC_14_10_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_11_LC_14_10_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_11_LC_14_10_4 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_11_LC_14_10_4  (
            .in0(N__42622),
            .in1(N__35011),
            .in2(N__39350),
            .in3(N__42379),
            .lcout(measured_delay_hc_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47283),
            .ce(),
            .sr(N__46618));
    defparam \delay_measurement_inst.delay_hc_reg_12_LC_14_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_12_LC_14_10_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_12_LC_14_10_5 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_12_LC_14_10_5  (
            .in0(N__42380),
            .in1(N__34985),
            .in2(N__39405),
            .in3(N__42623),
            .lcout(measured_delay_hc_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47283),
            .ce(),
            .sr(N__46618));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto13_3_1_LC_14_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto13_3_1_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto13_3_1_LC_14_10_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto13_3_1_LC_14_10_6  (
            .in0(N__39379),
            .in1(N__39331),
            .in2(N__44273),
            .in3(N__35657),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un1_startlto13_3Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto13_3_LC_14_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto13_3_LC_14_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto13_3_LC_14_10_7 .LUT_INIT=16'b0101000001110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto13_3_LC_14_10_7  (
            .in0(N__34029),
            .in1(N__41756),
            .in2(N__33722),
            .in3(N__41671),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_1_LC_14_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_1_LC_14_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_1_LC_14_11_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_26_1_LC_14_11_4  (
            .in0(N__42019),
            .in1(N__33711),
            .in2(N__42682),
            .in3(N__42049),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_20_LC_14_11_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_20_LC_14_11_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_20_LC_14_11_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_20_LC_14_11_5  (
            .in0(N__33713),
            .in1(N__42620),
            .in2(_gnd_net_),
            .in3(N__42417),
            .lcout(measured_delay_hc_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47275),
            .ce(),
            .sr(N__46629));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_2_0_LC_14_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_2_0_LC_14_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_2_0_LC_14_11_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto30_2_0_LC_14_11_6  (
            .in0(N__42020),
            .in1(N__33712),
            .in2(N__42683),
            .in3(N__41876),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un1_startlto30_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_3_LC_14_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_3_LC_14_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto30_3_LC_14_11_7 .LUT_INIT=16'b0011000001110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto30_3_LC_14_11_7  (
            .in0(N__33903),
            .in1(N__35576),
            .in2(N__33701),
            .in3(N__33698),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlt31_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNII60D_0_LC_14_12_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNII60D_0_LC_14_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.stoper_state_RNII60D_0_LC_14_12_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \phase_controller_slave.stoper_tr.stoper_state_RNII60D_0_LC_14_12_5  (
            .in0(N__38045),
            .in1(N__37826),
            .in2(_gnd_net_),
            .in3(N__38117),
            .lcout(\phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.start_timer_tr_LC_14_13_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_tr_LC_14_13_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.start_timer_tr_LC_14_13_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \delay_measurement_inst.start_timer_tr_LC_14_13_0  (
            .in0(N__34905),
            .in1(N__33833),
            .in2(_gnd_net_),
            .in3(N__33805),
            .lcout(\delay_measurement_inst.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47255),
            .ce(),
            .sr(N__46641));
    defparam \delay_measurement_inst.prev_tr_sig_LC_14_13_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.prev_tr_sig_LC_14_13_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.prev_tr_sig_LC_14_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.prev_tr_sig_LC_14_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34906),
            .lcout(\delay_measurement_inst.prev_tr_sigZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47255),
            .ce(),
            .sr(N__46641));
    defparam \delay_measurement_inst.tr_state_RNIMR6L_0_LC_14_13_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.tr_state_RNIMR6L_0_LC_14_13_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.tr_state_RNIMR6L_0_LC_14_13_2 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \delay_measurement_inst.tr_state_RNIMR6L_0_LC_14_13_2  (
            .in0(N__34904),
            .in1(N__33832),
            .in2(_gnd_net_),
            .in3(N__33804),
            .lcout(\delay_measurement_inst.tr_state_RNIMR6LZ0Z_0 ),
            .ltout(\delay_measurement_inst.tr_state_RNIMR6LZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.stop_timer_tr_LC_14_13_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_tr_LC_14_13_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.stop_timer_tr_LC_14_13_3 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \delay_measurement_inst.stop_timer_tr_LC_14_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33791),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.stop_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47255),
            .ce(),
            .sr(N__46641));
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_14_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_14_13_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_14_13_4 .LUT_INIT=16'b0101111100001010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_LC_14_13_4  (
            .in0(N__39255),
            .in1(_gnd_net_),
            .in2(N__37405),
            .in3(N__37378),
            .lcout(\delay_measurement_inst.delay_tr_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47255),
            .ce(),
            .sr(N__46641));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_14_13_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_14_13_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_14_13_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_14_13_5  (
            .in0(_gnd_net_),
            .in1(N__37398),
            .in2(_gnd_net_),
            .in3(N__39254),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_323_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.T01_LC_14_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.T01_LC_14_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.T01_LC_14_13_7 .LUT_INIT=16'b1010101010111010;
    LogicCell40 \phase_controller_inst1.T01_LC_14_13_7  (
            .in0(N__33788),
            .in1(N__43117),
            .in2(N__34474),
            .in3(N__43152),
            .lcout(shift_flag_start),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47255),
            .ce(),
            .sr(N__46641));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_14_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_14_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_14_14_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_14_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33755),
            .lcout(\current_shift_inst.un4_control_input_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_14_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_14_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_14_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_14_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33740),
            .lcout(\current_shift_inst.un4_control_input_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_14_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_14_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_14_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_14_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33986),
            .lcout(\current_shift_inst.un4_control_input_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_14_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_14_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_14_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_14_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33968),
            .lcout(\current_shift_inst.un4_control_input_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_14_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_14_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_14_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_14_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33950),
            .lcout(\current_shift_inst.un4_control_input_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_14_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_14_15_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_14_15_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_10_LC_14_15_0  (
            .in0(N__47605),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39469),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47239),
            .ce(N__46858),
            .sr(N__46657));
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_14_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_14_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_14_15_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_12_LC_14_15_2  (
            .in0(N__47606),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39496),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47239),
            .ce(N__46858),
            .sr(N__46657));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_14_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_14_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_14_15_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_14_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33932),
            .lcout(\current_shift_inst.un4_control_input_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.target_time_0_LC_14_16_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_0_LC_14_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_0_LC_14_16_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_0_LC_14_16_0  (
            .in0(N__44164),
            .in1(N__43853),
            .in2(N__42259),
            .in3(N__40336),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47231),
            .ce(N__43700),
            .sr(N__46666));
    defparam \phase_controller_slave.stoper_hc.target_time_15_LC_14_16_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_15_LC_14_16_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_15_LC_14_16_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_15_LC_14_16_1  (
            .in0(N__43855),
            .in1(N__44166),
            .in2(_gnd_net_),
            .in3(N__33917),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47231),
            .ce(N__43700),
            .sr(N__46666));
    defparam \phase_controller_slave.stoper_hc.target_time_14_LC_14_16_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_14_LC_14_16_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_14_LC_14_16_3 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_14_LC_14_16_3  (
            .in0(N__43854),
            .in1(N__44165),
            .in2(_gnd_net_),
            .in3(N__33877),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47231),
            .ce(N__43700),
            .sr(N__46666));
    defparam \phase_controller_slave.stoper_hc.target_timeZ0Z_6_LC_14_16_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_timeZ0Z_6_LC_14_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_timeZ0Z_6_LC_14_16_6 .LUT_INIT=16'b0000001000000011;
    LogicCell40 \phase_controller_slave.stoper_hc.target_timeZ0Z_6_LC_14_16_6  (
            .in0(N__34165),
            .in1(N__40335),
            .in2(N__44198),
            .in3(N__43852),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ1Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47231),
            .ce(N__43700),
            .sr(N__46666));
    defparam \phase_controller_slave.stoper_hc.target_time_10_LC_14_17_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_10_LC_14_17_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_10_LC_14_17_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_10_LC_14_17_0  (
            .in0(N__44167),
            .in1(N__35670),
            .in2(_gnd_net_),
            .in3(N__43856),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47226),
            .ce(N__43687),
            .sr(N__46676));
    defparam \phase_controller_slave.stoper_hc.target_time_3_LC_14_17_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_3_LC_14_17_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_3_LC_14_17_1 .LUT_INIT=16'b1111111110101000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_3_LC_14_17_1  (
            .in0(N__43860),
            .in1(N__40318),
            .in2(N__35518),
            .in3(N__44173),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47226),
            .ce(N__43687),
            .sr(N__46676));
    defparam \phase_controller_slave.stoper_hc.target_time_12_LC_14_17_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_12_LC_14_17_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_12_LC_14_17_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_12_LC_14_17_2  (
            .in0(N__44169),
            .in1(N__39406),
            .in2(_gnd_net_),
            .in3(N__43858),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47226),
            .ce(N__43687),
            .sr(N__46676));
    defparam \phase_controller_slave.stoper_hc.target_time_11_LC_14_17_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_11_LC_14_17_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_11_LC_14_17_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_11_LC_14_17_3  (
            .in0(N__43857),
            .in1(N__44168),
            .in2(_gnd_net_),
            .in3(N__39353),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47226),
            .ce(N__43687),
            .sr(N__46676));
    defparam \phase_controller_slave.stoper_hc.target_time_2_LC_14_17_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_2_LC_14_17_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_2_LC_14_17_4 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_2_LC_14_17_4  (
            .in0(N__40316),
            .in1(N__34115),
            .in2(N__44199),
            .in3(N__43859),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47226),
            .ce(N__43687),
            .sr(N__46676));
    defparam \phase_controller_slave.stoper_hc.target_time_9_LC_14_17_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_9_LC_14_17_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_9_LC_14_17_5 .LUT_INIT=16'b0000000000110001;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_9_LC_14_17_5  (
            .in0(N__43863),
            .in1(N__44178),
            .in2(N__34055),
            .in3(N__40319),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47226),
            .ce(N__43687),
            .sr(N__46676));
    defparam \phase_controller_slave.stoper_hc.target_time_4_LC_14_17_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_4_LC_14_17_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_4_LC_14_17_6 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_4_LC_14_17_6  (
            .in0(N__40317),
            .in1(N__35427),
            .in2(N__44200),
            .in3(N__43861),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47226),
            .ce(N__43687),
            .sr(N__46676));
    defparam \phase_controller_slave.stoper_hc.target_time_7_LC_14_17_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_7_LC_14_17_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_7_LC_14_17_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_7_LC_14_17_7  (
            .in0(N__43862),
            .in1(N__44177),
            .in2(_gnd_net_),
            .in3(N__41675),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47226),
            .ce(N__43687),
            .sr(N__46676));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_7_LC_14_18_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_7_LC_14_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_7_LC_14_18_0 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_7_LC_14_18_0  (
            .in0(N__40663),
            .in1(N__40860),
            .in2(N__41029),
            .in3(N__33998),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47223),
            .ce(),
            .sr(N__46681));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_8_LC_14_18_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_8_LC_14_18_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_8_LC_14_18_1 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_8_LC_14_18_1  (
            .in0(N__40859),
            .in1(N__41000),
            .in2(N__40667),
            .in3(N__34199),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47223),
            .ce(),
            .sr(N__46681));
    defparam \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_14_18_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_14_18_3 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_14_18_3  (
            .in0(N__40858),
            .in1(_gnd_net_),
            .in2(N__40666),
            .in3(N__40999),
            .lcout(\phase_controller_slave.stoper_hc.time_passed_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_14_18_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_14_18_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_14_18_4  (
            .in0(N__34439),
            .in1(N__34369),
            .in2(_gnd_net_),
            .in3(N__34411),
            .lcout(),
            .ltout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_1_LC_14_18_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_1_LC_14_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_1_LC_14_18_5 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_1_LC_14_18_5  (
            .in0(N__38024),
            .in1(N__37892),
            .in2(N__34172),
            .in3(N__38143),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47223),
            .ce(),
            .sr(N__46681));
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_0_LC_14_18_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_0_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_0_LC_14_18_6 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_0_LC_14_18_6  (
            .in0(N__40998),
            .in1(N__40640),
            .in2(_gnd_net_),
            .in3(N__40857),
            .lcout(\phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_10_LC_14_18_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_10_LC_14_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_10_LC_14_18_7 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_10_LC_14_18_7  (
            .in0(N__37858),
            .in1(N__38142),
            .in2(N__38047),
            .in3(N__34619),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47223),
            .ce(),
            .sr(N__46681));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_2_LC_14_19_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_2_LC_14_19_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_2_LC_14_19_0 .LUT_INIT=16'b1010101010000010;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_2_LC_14_19_0  (
            .in0(N__34334),
            .in1(N__37875),
            .in2(N__38046),
            .in3(N__38173),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47217),
            .ce(),
            .sr(N__46689));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_3_LC_14_19_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_3_LC_14_19_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_3_LC_14_19_1 .LUT_INIT=16'b1100100011000100;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_3_LC_14_19_1  (
            .in0(N__37873),
            .in1(N__34298),
            .in2(N__38179),
            .in3(N__38022),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47217),
            .ce(),
            .sr(N__46689));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_4_LC_14_19_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_4_LC_14_19_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_4_LC_14_19_2 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_4_LC_14_19_2  (
            .in0(N__38015),
            .in1(N__37876),
            .in2(N__34268),
            .in3(N__38165),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47217),
            .ce(),
            .sr(N__46689));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_5_LC_14_19_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_5_LC_14_19_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_5_LC_14_19_3 .LUT_INIT=16'b1100100011000100;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_5_LC_14_19_3  (
            .in0(N__37874),
            .in1(N__34745),
            .in2(N__38180),
            .in3(N__38023),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47217),
            .ce(),
            .sr(N__46689));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_3_LC_14_19_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_3_LC_14_19_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_3_LC_14_19_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_3_LC_14_19_4  (
            .in0(N__41053),
            .in1(N__40664),
            .in2(N__40914),
            .in3(N__34238),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47217),
            .ce(),
            .sr(N__46689));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_7_LC_14_19_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_7_LC_14_19_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_7_LC_14_19_5 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_7_LC_14_19_5  (
            .in0(N__38164),
            .in1(N__38018),
            .in2(N__37899),
            .in3(N__34688),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47217),
            .ce(),
            .sr(N__46689));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_8_LC_14_19_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_8_LC_14_19_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_8_LC_14_19_6 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_8_LC_14_19_6  (
            .in0(N__38016),
            .in1(N__37877),
            .in2(N__34655),
            .in3(N__38166),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47217),
            .ce(),
            .sr(N__46689));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_6_LC_14_19_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_6_LC_14_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_6_LC_14_19_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_6_LC_14_19_7  (
            .in0(N__38163),
            .in1(N__38017),
            .in2(N__37898),
            .in3(N__34715),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47217),
            .ce(),
            .sr(N__46689));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_3_LC_14_20_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_3_LC_14_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_3_LC_14_20_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_3_LC_14_20_1  (
            .in0(N__43205),
            .in1(N__41568),
            .in2(N__43296),
            .in3(N__44386),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_5_3_LC_14_20_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_5_3_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_5_3_LC_14_20_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_5_3_LC_14_20_2  (
            .in0(N__40164),
            .in1(N__43497),
            .in2(N__34226),
            .in3(N__47824),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_5Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_15_LC_14_20_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_15_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_15_LC_14_20_4 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_15_LC_14_20_4  (
            .in0(N__44387),
            .in1(N__43206),
            .in2(N__41575),
            .in3(N__43289),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNIDEUE_0_LC_14_20_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNIDEUE_0_LC_14_20_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.stoper_state_RNIDEUE_0_LC_14_20_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.stoper_state_RNIDEUE_0_LC_14_20_5  (
            .in0(_gnd_net_),
            .in1(N__41022),
            .in2(_gnd_net_),
            .in3(N__40628),
            .lcout(\phase_controller_slave.stoper_hc.time_passed11 ),
            .ltout(\phase_controller_slave.stoper_hc.time_passed11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_20_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_20_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_20_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34211),
            .in3(N__40716),
            .lcout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSR_LC_14_20_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSR_LC_14_20_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSR_LC_14_20_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSR_LC_14_20_7  (
            .in0(N__40717),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37062),
            .lcout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1B6_LC_14_21_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1B6_LC_14_21_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1B6_LC_14_21_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1B6_LC_14_21_1  (
            .in0(_gnd_net_),
            .in1(N__34432),
            .in2(_gnd_net_),
            .in3(N__34403),
            .lcout(\phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.un1_start_LC_14_21_3 .C_ON=1'b0;
    defparam \phase_controller_slave.un1_start_LC_14_21_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.un1_start_LC_14_21_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_slave.un1_start_LC_14_21_3  (
            .in0(N__34557),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34475),
            .lcout(\phase_controller_slave.un1_startZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_21_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_21_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_21_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_21_7  (
            .in0(_gnd_net_),
            .in1(N__34431),
            .in2(_gnd_net_),
            .in3(N__34402),
            .lcout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_14_22_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_14_22_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_14_22_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_14_22_0  (
            .in0(_gnd_net_),
            .in1(N__34379),
            .in2(N__34373),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_22_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_14_22_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_14_22_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_14_22_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_14_22_1  (
            .in0(_gnd_net_),
            .in1(N__34349),
            .in2(_gnd_net_),
            .in3(N__34325),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_14_22_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_14_22_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_14_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_14_22_2  (
            .in0(_gnd_net_),
            .in1(N__34322),
            .in2(N__34316),
            .in3(N__34286),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_14_22_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_14_22_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_14_22_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_14_22_3  (
            .in0(_gnd_net_),
            .in1(N__34283),
            .in2(_gnd_net_),
            .in3(N__34256),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_14_22_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_14_22_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_14_22_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_14_22_4  (
            .in0(_gnd_net_),
            .in1(N__34253),
            .in2(_gnd_net_),
            .in3(N__34733),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_14_22_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_14_22_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_14_22_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_14_22_5  (
            .in0(_gnd_net_),
            .in1(N__34730),
            .in2(_gnd_net_),
            .in3(N__34706),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_14_22_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_14_22_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_14_22_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_14_22_6  (
            .in0(_gnd_net_),
            .in1(N__34703),
            .in2(_gnd_net_),
            .in3(N__34673),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_14_22_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_14_22_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_14_22_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_14_22_7  (
            .in0(_gnd_net_),
            .in1(N__34670),
            .in2(_gnd_net_),
            .in3(N__34643),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_14_23_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_14_23_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_14_23_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_14_23_0  (
            .in0(_gnd_net_),
            .in1(N__37513),
            .in2(_gnd_net_),
            .in3(N__34640),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9 ),
            .ltout(),
            .carryin(bfn_14_23_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_14_23_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_14_23_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_14_23_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_14_23_1  (
            .in0(_gnd_net_),
            .in1(N__34637),
            .in2(_gnd_net_),
            .in3(N__34610),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_14_23_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_14_23_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_14_23_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_14_23_2  (
            .in0(_gnd_net_),
            .in1(N__34606),
            .in2(_gnd_net_),
            .in3(N__34586),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_14_23_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_14_23_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_14_23_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_14_23_3  (
            .in0(_gnd_net_),
            .in1(N__37651),
            .in2(_gnd_net_),
            .in3(N__34583),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_14_23_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_14_23_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_14_23_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_14_23_4  (
            .in0(_gnd_net_),
            .in1(N__37537),
            .in2(_gnd_net_),
            .in3(N__34580),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_14_23_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_14_23_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_14_23_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_14_23_5  (
            .in0(_gnd_net_),
            .in1(N__38320),
            .in2(_gnd_net_),
            .in3(N__34781),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_14_23_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_14_23_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_14_23_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_14_23_6  (
            .in0(_gnd_net_),
            .in1(N__37675),
            .in2(_gnd_net_),
            .in3(N__34778),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_14_23_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_14_23_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_14_23_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_14_23_7  (
            .in0(_gnd_net_),
            .in1(N__37627),
            .in2(_gnd_net_),
            .in3(N__34775),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_14_24_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_14_24_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_14_24_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_14_24_0  (
            .in0(_gnd_net_),
            .in1(N__38218),
            .in2(_gnd_net_),
            .in3(N__34772),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17 ),
            .ltout(),
            .carryin(bfn_14_24_0_),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_14_24_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_14_24_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_14_24_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_14_24_1  (
            .in0(_gnd_net_),
            .in1(N__38194),
            .in2(_gnd_net_),
            .in3(N__34769),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_14_24_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_14_24_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_14_24_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_14_24_2  (
            .in0(_gnd_net_),
            .in1(N__37756),
            .in2(_gnd_net_),
            .in3(N__34766),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_13_LC_14_25_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_13_LC_14_25_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_13_LC_14_25_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_13_LC_14_25_0  (
            .in0(N__41066),
            .in1(N__40680),
            .in2(N__40909),
            .in3(N__34763),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47196),
            .ce(),
            .sr(N__46726));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_17_LC_14_25_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_17_LC_14_25_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_17_LC_14_25_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_17_LC_14_25_4  (
            .in0(N__41067),
            .in1(N__40681),
            .in2(N__40910),
            .in3(N__34757),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47196),
            .ce(),
            .sr(N__46726));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_18_LC_14_25_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_18_LC_14_25_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_18_LC_14_25_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_18_LC_14_25_7  (
            .in0(N__40679),
            .in1(N__41068),
            .in2(N__40917),
            .in3(N__34751),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47196),
            .ce(),
            .sr(N__46726));
    defparam SB_DFF_inst_DELAY_TR1_LC_15_5_1.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_TR1_LC_15_5_1.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_TR1_LC_15_5_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_DELAY_TR1_LC_15_5_1 (
            .in0(N__34925),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(delay_tr_d1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47334),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_DELAY_TR2_LC_15_5_4.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_TR2_LC_15_5_4.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_TR2_LC_15_5_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_DELAY_TR2_LC_15_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34916),
            .lcout(delay_tr_d2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47334),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHUIH1_4_LC_15_6_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHUIH1_4_LC_15_6_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHUIH1_4_LC_15_6_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHUIH1_4_LC_15_6_2  (
            .in0(N__41696),
            .in1(N__35448),
            .in2(N__41797),
            .in3(N__35258),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_15_6_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_15_6_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_15_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_15_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38456),
            .lcout(\delay_measurement_inst.elapsed_time_hc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47327),
            .ce(N__35695),
            .sr(N__46597));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_15_6_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_15_6_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_15_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_15_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38435),
            .lcout(\delay_measurement_inst.elapsed_time_hc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47327),
            .ce(N__35695),
            .sr(N__46597));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOKRB1_10_LC_15_6_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOKRB1_10_LC_15_6_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOKRB1_10_LC_15_6_7 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOKRB1_10_LC_15_6_7  (
            .in0(N__35539),
            .in1(N__42130),
            .in2(N__35038),
            .in3(N__34840),
            .lcout(\delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_15_7_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_15_7_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_15_7_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_15_7_0  (
            .in0(_gnd_net_),
            .in1(N__38455),
            .in2(N__38413),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.elapsed_time_hc_3 ),
            .ltout(),
            .carryin(bfn_15_7_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__47319),
            .ce(N__35696),
            .sr(N__46600));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_15_7_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_15_7_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_15_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_15_7_1  (
            .in0(_gnd_net_),
            .in1(N__38434),
            .in2(N__38389),
            .in3(N__34817),
            .lcout(\delay_measurement_inst.elapsed_time_hc_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__47319),
            .ce(N__35696),
            .sr(N__46600));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_15_7_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_15_7_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_15_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_15_7_2  (
            .in0(_gnd_net_),
            .in1(N__38364),
            .in2(N__38414),
            .in3(N__34784),
            .lcout(\delay_measurement_inst.elapsed_time_hc_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__47319),
            .ce(N__35696),
            .sr(N__46600));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_15_7_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_15_7_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_15_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_15_7_3  (
            .in0(_gnd_net_),
            .in1(N__38346),
            .in2(N__38390),
            .in3(N__35090),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__47319),
            .ce(N__35696),
            .sr(N__46600));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_15_7_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_15_7_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_15_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_15_7_4  (
            .in0(_gnd_net_),
            .in1(N__38365),
            .in2(N__38698),
            .in3(N__35087),
            .lcout(\delay_measurement_inst.elapsed_time_hc_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__47319),
            .ce(N__35696),
            .sr(N__46600));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_15_7_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_15_7_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_15_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_15_7_5  (
            .in0(_gnd_net_),
            .in1(N__38347),
            .in2(N__38674),
            .in3(N__35084),
            .lcout(\delay_measurement_inst.elapsed_time_hc_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__47319),
            .ce(N__35696),
            .sr(N__46600));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_15_7_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_15_7_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_15_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_15_7_6  (
            .in0(_gnd_net_),
            .in1(N__38651),
            .in2(N__38699),
            .in3(N__35042),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__47319),
            .ce(N__35696),
            .sr(N__46600));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_15_7_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_15_7_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_15_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_15_7_7  (
            .in0(_gnd_net_),
            .in1(N__38627),
            .in2(N__38675),
            .in3(N__35015),
            .lcout(\delay_measurement_inst.elapsed_time_hc_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__47319),
            .ce(N__35696),
            .sr(N__46600));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_15_8_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_15_8_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_15_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_15_8_0  (
            .in0(_gnd_net_),
            .in1(N__38650),
            .in2(N__38602),
            .in3(N__34988),
            .lcout(\delay_measurement_inst.elapsed_time_hc_11 ),
            .ltout(),
            .carryin(bfn_15_8_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__47311),
            .ce(N__35697),
            .sr(N__46605));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_15_8_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_15_8_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_15_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_15_8_1  (
            .in0(_gnd_net_),
            .in1(N__38626),
            .in2(N__38578),
            .in3(N__34964),
            .lcout(\delay_measurement_inst.elapsed_time_hc_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__47311),
            .ce(N__35697),
            .sr(N__46605));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_15_8_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_15_8_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_15_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_15_8_2  (
            .in0(_gnd_net_),
            .in1(N__38553),
            .in2(N__38603),
            .in3(N__34928),
            .lcout(\delay_measurement_inst.elapsed_time_hc_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__47311),
            .ce(N__35697),
            .sr(N__46605));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_15_8_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_15_8_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_15_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_15_8_3  (
            .in0(_gnd_net_),
            .in1(N__38535),
            .in2(N__38579),
            .in3(N__35270),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__47311),
            .ce(N__35697),
            .sr(N__46605));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_15_8_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_15_8_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_15_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_15_8_4  (
            .in0(_gnd_net_),
            .in1(N__38554),
            .in2(N__38878),
            .in3(N__35213),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__47311),
            .ce(N__35697),
            .sr(N__46605));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_15_8_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_15_8_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_15_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_15_8_5  (
            .in0(_gnd_net_),
            .in1(N__38536),
            .in2(N__38854),
            .in3(N__35183),
            .lcout(\delay_measurement_inst.elapsed_time_hc_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__47311),
            .ce(N__35697),
            .sr(N__46605));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_15_8_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_15_8_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_15_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_15_8_6  (
            .in0(_gnd_net_),
            .in1(N__38831),
            .in2(N__38879),
            .in3(N__35180),
            .lcout(\delay_measurement_inst.elapsed_time_hc_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__47311),
            .ce(N__35697),
            .sr(N__46605));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_15_8_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_15_8_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_15_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_15_8_7  (
            .in0(_gnd_net_),
            .in1(N__38807),
            .in2(N__38855),
            .in3(N__35177),
            .lcout(\delay_measurement_inst.elapsed_time_hc_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__47311),
            .ce(N__35697),
            .sr(N__46605));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_15_9_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_15_9_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_15_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_15_9_0  (
            .in0(_gnd_net_),
            .in1(N__38830),
            .in2(N__38782),
            .in3(N__35174),
            .lcout(\delay_measurement_inst.elapsed_time_hc_19 ),
            .ltout(),
            .carryin(bfn_15_9_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__47299),
            .ce(N__35698),
            .sr(N__46610));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_15_9_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_15_9_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_15_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_15_9_1  (
            .in0(_gnd_net_),
            .in1(N__38806),
            .in2(N__38758),
            .in3(N__35159),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__47299),
            .ce(N__35698),
            .sr(N__46610));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_15_9_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_15_9_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_15_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_15_9_2  (
            .in0(_gnd_net_),
            .in1(N__38733),
            .in2(N__38783),
            .in3(N__35147),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__47299),
            .ce(N__35698),
            .sr(N__46610));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_15_9_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_15_9_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_15_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_15_9_3  (
            .in0(_gnd_net_),
            .in1(N__38715),
            .in2(N__38759),
            .in3(N__35132),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__47299),
            .ce(N__35698),
            .sr(N__46610));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_15_9_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_15_9_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_15_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_15_9_4  (
            .in0(_gnd_net_),
            .in1(N__38734),
            .in2(N__39232),
            .in3(N__35363),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__47299),
            .ce(N__35698),
            .sr(N__46610));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_15_9_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_15_9_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_15_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_15_9_5  (
            .in0(_gnd_net_),
            .in1(N__38716),
            .in2(N__39208),
            .in3(N__35354),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__47299),
            .ce(N__35698),
            .sr(N__46610));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_15_9_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_15_9_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_15_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_15_9_6  (
            .in0(_gnd_net_),
            .in1(N__39185),
            .in2(N__39233),
            .in3(N__35345),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__47299),
            .ce(N__35698),
            .sr(N__46610));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_15_9_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_15_9_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_15_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_15_9_7  (
            .in0(_gnd_net_),
            .in1(N__39161),
            .in2(N__39209),
            .in3(N__35333),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__47299),
            .ce(N__35698),
            .sr(N__46610));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_15_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_15_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_15_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_15_10_0  (
            .in0(_gnd_net_),
            .in1(N__39184),
            .in2(N__39136),
            .in3(N__35330),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ),
            .ltout(),
            .carryin(bfn_15_10_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__47290),
            .ce(N__35699),
            .sr(N__46614));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_15_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_15_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_15_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_15_10_1  (
            .in0(_gnd_net_),
            .in1(N__39160),
            .in2(N__39112),
            .in3(N__35327),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__47290),
            .ce(N__35699),
            .sr(N__46614));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_15_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_15_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_15_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_15_10_2  (
            .in0(_gnd_net_),
            .in1(N__39088),
            .in2(N__39137),
            .in3(N__35324),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__47290),
            .ce(N__35699),
            .sr(N__46614));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_15_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_15_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_15_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_15_10_3  (
            .in0(_gnd_net_),
            .in1(N__38935),
            .in2(N__39113),
            .in3(N__35321),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__47290),
            .ce(N__35699),
            .sr(N__46614));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_15_10_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_15_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_15_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_15_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35318),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47290),
            .ce(N__35699),
            .sr(N__46614));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_15_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_15_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_15_11_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_15_11_2  (
            .in0(N__41660),
            .in1(N__43955),
            .in2(N__41763),
            .in3(N__35656),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_15_11_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_15_11_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_15_11_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_15_11_5  (
            .in0(N__35624),
            .in1(N__35618),
            .in2(N__35612),
            .in3(N__35603),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_15_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_15_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_15_11_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_15_11_6  (
            .in0(N__40440),
            .in1(N__42183),
            .in2(N__42053),
            .in3(N__42339),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_15_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_15_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_15_11_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIUKI8_LC_15_11_7  (
            .in0(N__35570),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.timer_s1.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_3_LC_15_12_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_3_LC_15_12_0 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_hc_reg_3_LC_15_12_0 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_3_LC_15_12_0  (
            .in0(N__42649),
            .in1(N__35543),
            .in2(N__35500),
            .in3(N__42442),
            .lcout(measured_delay_hc_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47276),
            .ce(),
            .sr(N__46630));
    defparam \delay_measurement_inst.delay_hc_reg_4_LC_15_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_4_LC_15_12_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_4_LC_15_12_1 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_4_LC_15_12_1  (
            .in0(N__42443),
            .in1(N__42650),
            .in2(N__35422),
            .in3(N__35453),
            .lcout(measured_delay_hc_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47276),
            .ce(),
            .sr(N__46630));
    defparam \delay_measurement_inst.delay_tr_reg_15_LC_15_12_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_15_LC_15_12_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_15_LC_15_12_3 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_15_LC_15_12_3  (
            .in0(N__45159),
            .in1(N__47487),
            .in2(N__47806),
            .in3(N__47723),
            .lcout(measured_delay_tr_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47276),
            .ce(),
            .sr(N__46630));
    defparam \delay_measurement_inst.delay_tr_reg_7_LC_15_12_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_7_LC_15_12_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_7_LC_15_12_4 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_7_LC_15_12_4  (
            .in0(N__47724),
            .in1(N__43594),
            .in2(N__37313),
            .in3(N__44717),
            .lcout(measured_delay_tr_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47276),
            .ce(),
            .sr(N__46630));
    defparam \delay_measurement_inst.delay_tr_reg_8_LC_15_12_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_8_LC_15_12_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_8_LC_15_12_5 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_8_LC_15_12_5  (
            .in0(N__44663),
            .in1(N__37202),
            .in2(N__43603),
            .in3(N__47725),
            .lcout(measured_delay_tr_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47276),
            .ce(),
            .sr(N__46630));
    defparam \delay_measurement_inst.start_timer_hc_LC_15_12_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_hc_LC_15_12_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.start_timer_hc_LC_15_12_6 .LUT_INIT=16'b1001100110101010;
    LogicCell40 \delay_measurement_inst.start_timer_hc_LC_15_12_6  (
            .in0(N__35929),
            .in1(N__35868),
            .in2(_gnd_net_),
            .in3(N__41931),
            .lcout(\delay_measurement_inst.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47276),
            .ce(),
            .sr(N__46630));
    defparam \delay_measurement_inst.prev_hc_sig_LC_15_12_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.prev_hc_sig_LC_15_12_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.prev_hc_sig_LC_15_12_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \delay_measurement_inst.prev_hc_sig_LC_15_12_7  (
            .in0(N__41932),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.prev_hc_sigZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47276),
            .ce(),
            .sr(N__46630));
    defparam \current_shift_inst.timer_s1.counter_0_LC_15_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_0_LC_15_13_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_0_LC_15_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_0_LC_15_13_0  (
            .in0(N__36533),
            .in1(N__35850),
            .in2(_gnd_net_),
            .in3(N__35831),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_15_13_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_0 ),
            .clk(N__47264),
            .ce(N__36409),
            .sr(N__46635));
    defparam \current_shift_inst.timer_s1.counter_1_LC_15_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_1_LC_15_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_1_LC_15_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_1_LC_15_13_1  (
            .in0(N__36541),
            .in1(N__35820),
            .in2(_gnd_net_),
            .in3(N__35801),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_0 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_1 ),
            .clk(N__47264),
            .ce(N__36409),
            .sr(N__46635));
    defparam \current_shift_inst.timer_s1.counter_2_LC_15_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_2_LC_15_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_2_LC_15_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_2_LC_15_13_2  (
            .in0(N__36534),
            .in1(N__35796),
            .in2(_gnd_net_),
            .in3(N__35780),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_1 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_2 ),
            .clk(N__47264),
            .ce(N__36409),
            .sr(N__46635));
    defparam \current_shift_inst.timer_s1.counter_3_LC_15_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_3_LC_15_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_3_LC_15_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_3_LC_15_13_3  (
            .in0(N__36542),
            .in1(N__35775),
            .in2(_gnd_net_),
            .in3(N__35759),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_3 ),
            .clk(N__47264),
            .ce(N__36409),
            .sr(N__46635));
    defparam \current_shift_inst.timer_s1.counter_4_LC_15_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_4_LC_15_13_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_4_LC_15_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_4_LC_15_13_4  (
            .in0(N__36535),
            .in1(N__35743),
            .in2(_gnd_net_),
            .in3(N__35729),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_4 ),
            .clk(N__47264),
            .ce(N__36409),
            .sr(N__46635));
    defparam \current_shift_inst.timer_s1.counter_5_LC_15_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_5_LC_15_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_5_LC_15_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_5_LC_15_13_5  (
            .in0(N__36543),
            .in1(N__35718),
            .in2(_gnd_net_),
            .in3(N__35702),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_5 ),
            .clk(N__47264),
            .ce(N__36409),
            .sr(N__46635));
    defparam \current_shift_inst.timer_s1.counter_6_LC_15_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_6_LC_15_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_6_LC_15_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_6_LC_15_13_6  (
            .in0(N__36536),
            .in1(N__36129),
            .in2(_gnd_net_),
            .in3(N__36113),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_6 ),
            .clk(N__47264),
            .ce(N__36409),
            .sr(N__46635));
    defparam \current_shift_inst.timer_s1.counter_7_LC_15_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_7_LC_15_13_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_7_LC_15_13_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_7_LC_15_13_7  (
            .in0(N__36544),
            .in1(N__36108),
            .in2(_gnd_net_),
            .in3(N__36092),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_7 ),
            .clk(N__47264),
            .ce(N__36409),
            .sr(N__46635));
    defparam \current_shift_inst.timer_s1.counter_8_LC_15_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_8_LC_15_14_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_8_LC_15_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_8_LC_15_14_0  (
            .in0(N__36548),
            .in1(N__36078),
            .in2(_gnd_net_),
            .in3(N__36059),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_15_14_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_8 ),
            .clk(N__47256),
            .ce(N__36407),
            .sr(N__46642));
    defparam \current_shift_inst.timer_s1.counter_9_LC_15_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_9_LC_15_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_9_LC_15_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_9_LC_15_14_1  (
            .in0(N__36540),
            .in1(N__36045),
            .in2(_gnd_net_),
            .in3(N__36029),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_9 ),
            .clk(N__47256),
            .ce(N__36407),
            .sr(N__46642));
    defparam \current_shift_inst.timer_s1.counter_10_LC_15_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_10_LC_15_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_10_LC_15_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_10_LC_15_14_2  (
            .in0(N__36545),
            .in1(N__36018),
            .in2(_gnd_net_),
            .in3(N__36002),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_9 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_10 ),
            .clk(N__47256),
            .ce(N__36407),
            .sr(N__46642));
    defparam \current_shift_inst.timer_s1.counter_11_LC_15_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_11_LC_15_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_11_LC_15_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_11_LC_15_14_3  (
            .in0(N__36537),
            .in1(N__35991),
            .in2(_gnd_net_),
            .in3(N__35975),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_11 ),
            .clk(N__47256),
            .ce(N__36407),
            .sr(N__46642));
    defparam \current_shift_inst.timer_s1.counter_12_LC_15_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_12_LC_15_14_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_12_LC_15_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_12_LC_15_14_4  (
            .in0(N__36546),
            .in1(N__35970),
            .in2(_gnd_net_),
            .in3(N__35954),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_12 ),
            .clk(N__47256),
            .ce(N__36407),
            .sr(N__46642));
    defparam \current_shift_inst.timer_s1.counter_13_LC_15_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_13_LC_15_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_13_LC_15_14_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_13_LC_15_14_5  (
            .in0(N__36538),
            .in1(N__35949),
            .in2(_gnd_net_),
            .in3(N__35933),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_13 ),
            .clk(N__47256),
            .ce(N__36407),
            .sr(N__46642));
    defparam \current_shift_inst.timer_s1.counter_14_LC_15_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_14_LC_15_14_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_14_LC_15_14_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_14_LC_15_14_6  (
            .in0(N__36547),
            .in1(N__36357),
            .in2(_gnd_net_),
            .in3(N__36341),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_14 ),
            .clk(N__47256),
            .ce(N__36407),
            .sr(N__46642));
    defparam \current_shift_inst.timer_s1.counter_15_LC_15_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_15_LC_15_14_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_15_LC_15_14_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_15_LC_15_14_7  (
            .in0(N__36539),
            .in1(N__36330),
            .in2(_gnd_net_),
            .in3(N__36314),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_15 ),
            .clk(N__47256),
            .ce(N__36407),
            .sr(N__46642));
    defparam \current_shift_inst.timer_s1.counter_16_LC_15_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_16_LC_15_15_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_16_LC_15_15_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_16_LC_15_15_0  (
            .in0(N__36519),
            .in1(N__36303),
            .in2(_gnd_net_),
            .in3(N__36284),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_15_15_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_16 ),
            .clk(N__47247),
            .ce(N__36410),
            .sr(N__46648));
    defparam \current_shift_inst.timer_s1.counter_17_LC_15_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_17_LC_15_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_17_LC_15_15_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_17_LC_15_15_1  (
            .in0(N__36523),
            .in1(N__36276),
            .in2(_gnd_net_),
            .in3(N__36257),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_17 ),
            .clk(N__47247),
            .ce(N__36410),
            .sr(N__46648));
    defparam \current_shift_inst.timer_s1.counter_18_LC_15_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_18_LC_15_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_18_LC_15_15_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_18_LC_15_15_2  (
            .in0(N__36520),
            .in1(N__36246),
            .in2(_gnd_net_),
            .in3(N__36230),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_17 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_18 ),
            .clk(N__47247),
            .ce(N__36410),
            .sr(N__46648));
    defparam \current_shift_inst.timer_s1.counter_19_LC_15_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_19_LC_15_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_19_LC_15_15_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_19_LC_15_15_3  (
            .in0(N__36524),
            .in1(N__36219),
            .in2(_gnd_net_),
            .in3(N__36203),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_19 ),
            .clk(N__47247),
            .ce(N__36410),
            .sr(N__46648));
    defparam \current_shift_inst.timer_s1.counter_20_LC_15_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_20_LC_15_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_20_LC_15_15_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_20_LC_15_15_4  (
            .in0(N__36521),
            .in1(N__36198),
            .in2(_gnd_net_),
            .in3(N__36182),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_20 ),
            .clk(N__47247),
            .ce(N__36410),
            .sr(N__46648));
    defparam \current_shift_inst.timer_s1.counter_21_LC_15_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_21_LC_15_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_21_LC_15_15_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_21_LC_15_15_5  (
            .in0(N__36525),
            .in1(N__36177),
            .in2(_gnd_net_),
            .in3(N__36161),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_21 ),
            .clk(N__47247),
            .ce(N__36410),
            .sr(N__46648));
    defparam \current_shift_inst.timer_s1.counter_22_LC_15_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_22_LC_15_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_22_LC_15_15_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_22_LC_15_15_6  (
            .in0(N__36522),
            .in1(N__36150),
            .in2(_gnd_net_),
            .in3(N__36134),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_22 ),
            .clk(N__47247),
            .ce(N__36410),
            .sr(N__46648));
    defparam \current_shift_inst.timer_s1.counter_23_LC_15_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_23_LC_15_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_23_LC_15_15_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_23_LC_15_15_7  (
            .in0(N__36526),
            .in1(N__36693),
            .in2(_gnd_net_),
            .in3(N__36677),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_23 ),
            .clk(N__47247),
            .ce(N__36410),
            .sr(N__46648));
    defparam \current_shift_inst.timer_s1.counter_24_LC_15_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_24_LC_15_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_24_LC_15_16_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_24_LC_15_16_0  (
            .in0(N__36527),
            .in1(N__36669),
            .in2(_gnd_net_),
            .in3(N__36650),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_15_16_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_24 ),
            .clk(N__47240),
            .ce(N__36408),
            .sr(N__46658));
    defparam \current_shift_inst.timer_s1.counter_25_LC_15_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_25_LC_15_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_25_LC_15_16_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_25_LC_15_16_1  (
            .in0(N__36531),
            .in1(N__36642),
            .in2(_gnd_net_),
            .in3(N__36623),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_25 ),
            .clk(N__47240),
            .ce(N__36408),
            .sr(N__46658));
    defparam \current_shift_inst.timer_s1.counter_26_LC_15_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_26_LC_15_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_26_LC_15_16_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_26_LC_15_16_2  (
            .in0(N__36528),
            .in1(N__36612),
            .in2(_gnd_net_),
            .in3(N__36596),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_25 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_26 ),
            .clk(N__47240),
            .ce(N__36408),
            .sr(N__46658));
    defparam \current_shift_inst.timer_s1.counter_27_LC_15_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_27_LC_15_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_27_LC_15_16_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_27_LC_15_16_3  (
            .in0(N__36532),
            .in1(N__36585),
            .in2(_gnd_net_),
            .in3(N__36569),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_27 ),
            .clk(N__47240),
            .ce(N__36408),
            .sr(N__46658));
    defparam \current_shift_inst.timer_s1.counter_28_LC_15_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_28_LC_15_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_28_LC_15_16_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_28_LC_15_16_4  (
            .in0(N__36529),
            .in1(N__36565),
            .in2(_gnd_net_),
            .in3(N__36551),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_28 ),
            .clk(N__47240),
            .ce(N__36408),
            .sr(N__46658));
    defparam \current_shift_inst.timer_s1.counter_29_LC_15_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.counter_29_LC_15_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_29_LC_15_16_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \current_shift_inst.timer_s1.counter_29_LC_15_16_5  (
            .in0(N__36424),
            .in1(N__36530),
            .in2(_gnd_net_),
            .in3(N__36428),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47240),
            .ce(N__36408),
            .sr(N__46658));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0_c_LC_15_17_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0_c_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0_c_LC_15_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0_c_LC_15_17_0  (
            .in0(_gnd_net_),
            .in1(N__36371),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_17_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_15_17_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_15_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_15_17_1  (
            .in0(_gnd_net_),
            .in1(N__36854),
            .in2(N__41210),
            .in3(N__38286),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_15_17_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_15_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_15_17_2  (
            .in0(_gnd_net_),
            .in1(N__36839),
            .in2(N__36848),
            .in3(N__38251),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_15_17_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_15_17_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_15_17_3  (
            .in0(N__36826),
            .in1(N__36800),
            .in2(N__36809),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_15_17_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_15_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_15_17_4  (
            .in0(_gnd_net_),
            .in1(N__36785),
            .in2(N__36794),
            .in3(N__37597),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_15_17_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_15_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_15_17_5  (
            .in0(_gnd_net_),
            .in1(N__36779),
            .in2(N__43730),
            .in3(N__37564),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_15_17_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_15_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_15_17_6  (
            .in0(_gnd_net_),
            .in1(N__36764),
            .in2(N__36773),
            .in3(N__37486),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_15_17_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_15_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_15_17_7  (
            .in0(_gnd_net_),
            .in1(N__36731),
            .in2(N__36758),
            .in3(N__36742),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_15_18_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_15_18_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_15_18_0  (
            .in0(N__36718),
            .in1(N__36707),
            .in2(N__40466),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(bfn_15_18_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_15_18_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_15_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_15_18_1  (
            .in0(_gnd_net_),
            .in1(N__37034),
            .in2(N__37028),
            .in3(N__38510),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_15_18_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_15_18_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_15_18_2  (
            .in0(N__37732),
            .in1(N__37004),
            .in2(N__37019),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_15_18_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_15_18_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_15_18_3  (
            .in0(_gnd_net_),
            .in1(N__36986),
            .in2(N__36998),
            .in3(N__37706),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_15_18_4 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_15_18_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_15_18_4  (
            .in0(_gnd_net_),
            .in1(N__36947),
            .in2(N__36980),
            .in3(N__36968),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_15_18_5 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_15_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_15_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_15_18_5  (
            .in0(_gnd_net_),
            .in1(N__36920),
            .in2(N__44225),
            .in3(N__36941),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_15_18_6 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_15_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_15_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_15_18_6  (
            .in0(_gnd_net_),
            .in1(N__36881),
            .in2(N__36914),
            .in3(N__36899),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_15_18_7 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_15_18_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_15_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_15_18_7  (
            .in0(_gnd_net_),
            .in1(N__36860),
            .in2(N__36875),
            .in3(N__38477),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_15_19_0 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_15_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_15_19_0  (
            .in0(_gnd_net_),
            .in1(N__37160),
            .in2(N__40409),
            .in3(N__37181),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_16 ),
            .ltout(),
            .carryin(bfn_15_19_0_),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_15_19_1 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_15_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_15_19_1  (
            .in0(_gnd_net_),
            .in1(N__37136),
            .in2(N__40475),
            .in3(N__37154),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_17 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_15_19_2 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_15_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_15_19_2  (
            .in0(_gnd_net_),
            .in1(N__40400),
            .in2(N__37112),
            .in3(N__37130),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_15_19_3 .C_ON=1'b1;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_15_19_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_15_19_3  (
            .in0(N__37103),
            .in1(N__37085),
            .in2(N__40355),
            .in3(_gnd_net_),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_15_19_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_15_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_15_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_15_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37079),
            .lcout(\phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_2_LC_15_19_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_2_LC_15_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_2_LC_15_19_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_2_LC_15_19_6  (
            .in0(N__41437),
            .in1(N__37275),
            .in2(_gnd_net_),
            .in3(N__37361),
            .lcout(\phase_controller_inst1.stoper_tr.N_20_li ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_15_19_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_15_19_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_15_19_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_15_19_7  (
            .in0(N__37075),
            .in1(N__38287),
            .in2(_gnd_net_),
            .in3(N__40718),
            .lcout(\phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_15_20_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_15_20_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_15_20_0 .LUT_INIT=16'b1010001000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_2_LC_15_20_0  (
            .in0(N__40093),
            .in1(N__37437),
            .in2(N__40215),
            .in3(N__37455),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47218),
            .ce(N__46827),
            .sr(N__46690));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2_1_LC_15_20_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2_1_LC_15_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2_1_LC_15_20_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2_1_LC_15_20_1  (
            .in0(_gnd_net_),
            .in1(N__40205),
            .in2(_gnd_net_),
            .in3(N__40092),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_15_20_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_15_20_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_15_20_2 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_1_LC_15_20_2  (
            .in0(N__40117),
            .in1(N__37438),
            .in2(N__37469),
            .in3(N__37454),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47218),
            .ce(N__46827),
            .sr(N__46690));
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_15_20_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_15_20_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_15_20_3 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_3_LC_15_20_3  (
            .in0(N__37456),
            .in1(N__40206),
            .in2(_gnd_net_),
            .in3(N__37439),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47218),
            .ce(N__46827),
            .sr(N__46690));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_15_20_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_15_20_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_15_20_7 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_15_20_7  (
            .in0(N__37409),
            .in1(N__37385),
            .in2(_gnd_net_),
            .in3(N__39266),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_324_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_15_21_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_15_21_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_15_21_0 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_5_LC_15_21_0  (
            .in0(N__37279),
            .in1(N__41452),
            .in2(N__40177),
            .in3(N__37363),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47213),
            .ce(N__46857),
            .sr(N__46701));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_15_21_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_15_21_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_15_21_1 .LUT_INIT=16'b0100010001000101;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_LC_15_21_1  (
            .in0(N__37364),
            .in1(N__40250),
            .in2(N__41480),
            .in3(N__37280),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47213),
            .ce(N__46857),
            .sr(N__46701));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_15_21_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_15_21_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_15_21_2 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_LC_15_21_2  (
            .in0(N__37278),
            .in1(N__43502),
            .in2(N__41479),
            .in3(N__37362),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47213),
            .ce(N__46857),
            .sr(N__46701));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_15_21_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_15_21_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_15_21_3 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_LC_15_21_3  (
            .in0(N__41451),
            .in1(N__37327),
            .in2(_gnd_net_),
            .in3(N__37276),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47213),
            .ce(N__46857),
            .sr(N__46701));
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_15_21_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_15_21_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_15_21_4 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_8_LC_15_21_4  (
            .in0(N__37277),
            .in1(N__41453),
            .in2(_gnd_net_),
            .in3(N__37225),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47213),
            .ce(N__46857),
            .sr(N__46701));
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_15_21_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_15_21_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_15_21_6 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_14_LC_15_21_6  (
            .in0(N__41447),
            .in1(N__47539),
            .in2(_gnd_net_),
            .in3(N__47706),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47213),
            .ce(N__46857),
            .sr(N__46701));
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_15_21_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_15_21_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_15_21_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_17_LC_15_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43298),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47213),
            .ce(N__46857),
            .sr(N__46701));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_15_LC_15_22_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_15_LC_15_22_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_15_LC_15_22_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_15_LC_15_22_0  (
            .in0(N__37885),
            .in1(N__38162),
            .in2(N__38044),
            .in3(N__37685),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47210),
            .ce(),
            .sr(N__46708));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_12_LC_15_22_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_12_LC_15_22_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_12_LC_15_22_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_12_LC_15_22_2  (
            .in0(N__37884),
            .in1(N__38161),
            .in2(N__38043),
            .in3(N__37661),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47210),
            .ce(),
            .sr(N__46708));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_16_LC_15_22_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_16_LC_15_22_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_16_LC_15_22_3 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_16_LC_15_22_3  (
            .in0(N__38160),
            .in1(N__38005),
            .in2(N__37901),
            .in3(N__37637),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47210),
            .ce(),
            .sr(N__46708));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_4_LC_15_22_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_4_LC_15_22_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_4_LC_15_22_5 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_4_LC_15_22_5  (
            .in0(N__41054),
            .in1(N__40630),
            .in2(N__40902),
            .in3(N__37613),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47210),
            .ce(),
            .sr(N__46708));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_5_LC_15_22_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_5_LC_15_22_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_5_LC_15_22_6 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_5_LC_15_22_6  (
            .in0(N__40629),
            .in1(N__40872),
            .in2(N__41069),
            .in3(N__37580),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47210),
            .ce(),
            .sr(N__46708));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_13_LC_15_22_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_13_LC_15_22_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_13_LC_15_22_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_13_LC_15_22_7  (
            .in0(N__38159),
            .in1(N__38004),
            .in2(N__37900),
            .in3(N__37547),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47210),
            .ce(),
            .sr(N__46708));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_9_LC_15_23_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_9_LC_15_23_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_9_LC_15_23_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_9_LC_15_23_0  (
            .in0(N__37895),
            .in1(N__38178),
            .in2(N__38050),
            .in3(N__37523),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47207),
            .ce(),
            .sr(N__46712));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_6_LC_15_23_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_6_LC_15_23_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_6_LC_15_23_1 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_6_LC_15_23_1  (
            .in0(N__40632),
            .in1(N__40895),
            .in2(N__37499),
            .in3(N__41061),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47207),
            .ce(),
            .sr(N__46712));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_14_LC_15_23_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_14_LC_15_23_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_14_LC_15_23_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_14_LC_15_23_2  (
            .in0(N__37893),
            .in1(N__38176),
            .in2(N__38048),
            .in3(N__38330),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47207),
            .ce(),
            .sr(N__46712));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_1_LC_15_23_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_1_LC_15_23_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_1_LC_15_23_3 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_1_LC_15_23_3  (
            .in0(N__40631),
            .in1(N__40894),
            .in2(N__38306),
            .in3(N__41060),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47207),
            .ce(),
            .sr(N__46712));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_2_LC_15_23_4 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_2_LC_15_23_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_2_LC_15_23_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_2_LC_15_23_4  (
            .in0(N__41059),
            .in1(N__40633),
            .in2(N__40915),
            .in3(N__38264),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47207),
            .ce(),
            .sr(N__46712));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_17_LC_15_23_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_17_LC_15_23_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_17_LC_15_23_5 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_17_LC_15_23_5  (
            .in0(N__38174),
            .in1(N__38037),
            .in2(N__38234),
            .in3(N__37896),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47207),
            .ce(),
            .sr(N__46712));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_18_LC_15_23_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_18_LC_15_23_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_18_LC_15_23_6 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_18_LC_15_23_6  (
            .in0(N__37894),
            .in1(N__38177),
            .in2(N__38049),
            .in3(N__38204),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47207),
            .ce(),
            .sr(N__46712));
    defparam \phase_controller_slave.stoper_tr.accumulated_time_19_LC_15_23_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_19_LC_15_23_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.accumulated_time_19_LC_15_23_7 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_tr.accumulated_time_19_LC_15_23_7  (
            .in0(N__38175),
            .in1(N__38038),
            .in2(N__37910),
            .in3(N__37897),
            .lcout(\phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47207),
            .ce(),
            .sr(N__46712));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_10_LC_15_24_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_10_LC_15_24_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_10_LC_15_24_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_10_LC_15_24_2  (
            .in0(N__41062),
            .in1(N__40635),
            .in2(N__40900),
            .in3(N__37742),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47203),
            .ce(),
            .sr(N__46718));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_11_LC_15_24_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_11_LC_15_24_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_11_LC_15_24_3 .LUT_INIT=16'b1010100010100010;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_11_LC_15_24_3  (
            .in0(N__37715),
            .in1(N__40861),
            .in2(N__40665),
            .in3(N__41065),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47203),
            .ce(),
            .sr(N__46718));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_9_LC_15_24_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_9_LC_15_24_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_9_LC_15_24_6 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_9_LC_15_24_6  (
            .in0(N__41063),
            .in1(N__40636),
            .in2(N__40901),
            .in3(N__38519),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47203),
            .ce(),
            .sr(N__46718));
    defparam \phase_controller_slave.stoper_hc.accumulated_time_15_LC_15_24_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_15_LC_15_24_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.accumulated_time_15_LC_15_24_7 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_slave.stoper_hc.accumulated_time_15_LC_15_24_7  (
            .in0(N__40634),
            .in1(N__40862),
            .in2(N__38489),
            .in3(N__41064),
            .lcout(\phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47203),
            .ce(),
            .sr(N__46718));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_3_LC_16_6_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_3_LC_16_6_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_3_LC_16_6_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_3_LC_16_6_5  (
            .in0(_gnd_net_),
            .in1(N__41824),
            .in2(_gnd_net_),
            .in3(N__41836),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_16_7_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_16_7_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_16_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_0_LC_16_7_0  (
            .in0(N__39031),
            .in1(N__38454),
            .in2(_gnd_net_),
            .in3(N__38438),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_16_7_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .clk(N__47328),
            .ce(N__38909),
            .sr(N__46598));
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_16_7_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_16_7_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_16_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_1_LC_16_7_1  (
            .in0(N__39049),
            .in1(N__38433),
            .in2(_gnd_net_),
            .in3(N__38417),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .clk(N__47328),
            .ce(N__38909),
            .sr(N__46598));
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_16_7_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_16_7_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_16_7_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_2_LC_16_7_2  (
            .in0(N__39032),
            .in1(N__38412),
            .in2(_gnd_net_),
            .in3(N__38393),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .clk(N__47328),
            .ce(N__38909),
            .sr(N__46598));
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_16_7_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_16_7_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_16_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_3_LC_16_7_3  (
            .in0(N__39050),
            .in1(N__38388),
            .in2(_gnd_net_),
            .in3(N__38369),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .clk(N__47328),
            .ce(N__38909),
            .sr(N__46598));
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_16_7_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_16_7_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_16_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_4_LC_16_7_4  (
            .in0(N__39033),
            .in1(N__38366),
            .in2(_gnd_net_),
            .in3(N__38351),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .clk(N__47328),
            .ce(N__38909),
            .sr(N__46598));
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_16_7_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_16_7_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_16_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_5_LC_16_7_5  (
            .in0(N__39051),
            .in1(N__38348),
            .in2(_gnd_net_),
            .in3(N__38333),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .clk(N__47328),
            .ce(N__38909),
            .sr(N__46598));
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_16_7_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_16_7_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_16_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_6_LC_16_7_6  (
            .in0(N__39034),
            .in1(N__38697),
            .in2(_gnd_net_),
            .in3(N__38678),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .clk(N__47328),
            .ce(N__38909),
            .sr(N__46598));
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_16_7_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_16_7_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_16_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_7_LC_16_7_7  (
            .in0(N__39052),
            .in1(N__38673),
            .in2(_gnd_net_),
            .in3(N__38654),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .clk(N__47328),
            .ce(N__38909),
            .sr(N__46598));
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_16_8_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_16_8_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_16_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_8_LC_16_8_0  (
            .in0(N__39056),
            .in1(N__38649),
            .in2(_gnd_net_),
            .in3(N__38630),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_16_8_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .clk(N__47320),
            .ce(N__38916),
            .sr(N__46601));
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_16_8_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_16_8_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_16_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_9_LC_16_8_1  (
            .in0(N__39070),
            .in1(N__38625),
            .in2(_gnd_net_),
            .in3(N__38606),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .clk(N__47320),
            .ce(N__38916),
            .sr(N__46601));
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_16_8_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_16_8_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_16_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_10_LC_16_8_2  (
            .in0(N__39053),
            .in1(N__38601),
            .in2(_gnd_net_),
            .in3(N__38582),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .clk(N__47320),
            .ce(N__38916),
            .sr(N__46601));
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_16_8_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_16_8_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_16_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_11_LC_16_8_3  (
            .in0(N__39071),
            .in1(N__38577),
            .in2(_gnd_net_),
            .in3(N__38558),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .clk(N__47320),
            .ce(N__38916),
            .sr(N__46601));
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_16_8_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_16_8_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_16_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_12_LC_16_8_4  (
            .in0(N__39054),
            .in1(N__38555),
            .in2(_gnd_net_),
            .in3(N__38540),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .clk(N__47320),
            .ce(N__38916),
            .sr(N__46601));
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_16_8_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_16_8_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_16_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_13_LC_16_8_5  (
            .in0(N__39072),
            .in1(N__38537),
            .in2(_gnd_net_),
            .in3(N__38522),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .clk(N__47320),
            .ce(N__38916),
            .sr(N__46601));
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_16_8_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_16_8_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_16_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_14_LC_16_8_6  (
            .in0(N__39055),
            .in1(N__38877),
            .in2(_gnd_net_),
            .in3(N__38858),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .clk(N__47320),
            .ce(N__38916),
            .sr(N__46601));
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_16_8_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_16_8_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_16_8_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_15_LC_16_8_7  (
            .in0(N__39069),
            .in1(N__38853),
            .in2(_gnd_net_),
            .in3(N__38834),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .clk(N__47320),
            .ce(N__38916),
            .sr(N__46601));
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_16_9_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_16_9_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_16_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_16_LC_16_9_0  (
            .in0(N__39057),
            .in1(N__38829),
            .in2(_gnd_net_),
            .in3(N__38810),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_16_9_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .clk(N__47312),
            .ce(N__38917),
            .sr(N__46606));
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_16_9_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_16_9_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_16_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_17_LC_16_9_1  (
            .in0(N__39061),
            .in1(N__38805),
            .in2(_gnd_net_),
            .in3(N__38786),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .clk(N__47312),
            .ce(N__38917),
            .sr(N__46606));
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_16_9_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_16_9_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_16_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_18_LC_16_9_2  (
            .in0(N__39058),
            .in1(N__38781),
            .in2(_gnd_net_),
            .in3(N__38762),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .clk(N__47312),
            .ce(N__38917),
            .sr(N__46606));
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_16_9_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_16_9_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_16_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_19_LC_16_9_3  (
            .in0(N__39062),
            .in1(N__38757),
            .in2(_gnd_net_),
            .in3(N__38738),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .clk(N__47312),
            .ce(N__38917),
            .sr(N__46606));
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_16_9_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_16_9_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_16_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_20_LC_16_9_4  (
            .in0(N__39059),
            .in1(N__38735),
            .in2(_gnd_net_),
            .in3(N__38720),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .clk(N__47312),
            .ce(N__38917),
            .sr(N__46606));
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_16_9_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_16_9_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_16_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_21_LC_16_9_5  (
            .in0(N__39063),
            .in1(N__38717),
            .in2(_gnd_net_),
            .in3(N__38702),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .clk(N__47312),
            .ce(N__38917),
            .sr(N__46606));
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_16_9_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_16_9_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_16_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_22_LC_16_9_6  (
            .in0(N__39060),
            .in1(N__39231),
            .in2(_gnd_net_),
            .in3(N__39212),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .clk(N__47312),
            .ce(N__38917),
            .sr(N__46606));
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_16_9_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_16_9_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_16_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_23_LC_16_9_7  (
            .in0(N__39064),
            .in1(N__39207),
            .in2(_gnd_net_),
            .in3(N__39188),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .clk(N__47312),
            .ce(N__38917),
            .sr(N__46606));
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_16_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_16_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_16_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_24_LC_16_10_0  (
            .in0(N__39065),
            .in1(N__39183),
            .in2(_gnd_net_),
            .in3(N__39164),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_16_10_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .clk(N__47300),
            .ce(N__38924),
            .sr(N__46611));
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_16_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_16_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_16_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_25_LC_16_10_1  (
            .in0(N__39073),
            .in1(N__39159),
            .in2(_gnd_net_),
            .in3(N__39140),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .clk(N__47300),
            .ce(N__38924),
            .sr(N__46611));
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_16_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_16_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_16_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_26_LC_16_10_2  (
            .in0(N__39066),
            .in1(N__39135),
            .in2(_gnd_net_),
            .in3(N__39116),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .clk(N__47300),
            .ce(N__38924),
            .sr(N__46611));
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_16_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_16_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_16_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_27_LC_16_10_3  (
            .in0(N__39074),
            .in1(N__39111),
            .in2(_gnd_net_),
            .in3(N__39092),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .clk(N__47300),
            .ce(N__38924),
            .sr(N__46611));
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_16_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_16_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_16_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_28_LC_16_10_4  (
            .in0(N__39067),
            .in1(N__39089),
            .in2(_gnd_net_),
            .in3(N__39077),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ),
            .clk(N__47300),
            .ce(N__38924),
            .sr(N__46611));
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_16_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_16_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_16_10_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_29_LC_16_10_5  (
            .in0(N__38936),
            .in1(N__39068),
            .in2(_gnd_net_),
            .in3(N__38939),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47300),
            .ce(N__38924),
            .sr(N__46611));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_16_11_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_16_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_16_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_16_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43423),
            .lcout(\delay_measurement_inst.elapsed_time_tr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47291),
            .ce(N__45718),
            .sr(N__46615));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_9_LC_16_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_9_LC_16_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_9_LC_16_11_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_9_LC_16_11_7  (
            .in0(N__42319),
            .in1(N__39401),
            .in2(N__42182),
            .in3(N__39351),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5PP_2_LC_16_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5PP_2_LC_16_12_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5PP_2_LC_16_12_1 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5PP_2_LC_16_12_1  (
            .in0(N__42796),
            .in1(N__47781),
            .in2(N__43402),
            .in3(N__44870),
            .lcout(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI200N_7_LC_16_12_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI200N_7_LC_16_12_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI200N_7_LC_16_12_2 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI200N_7_LC_16_12_2  (
            .in0(N__44662),
            .in1(N__44716),
            .in2(_gnd_net_),
            .in3(N__39446),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC3FA_2_LC_16_12_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC3FA_2_LC_16_12_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC3FA_2_LC_16_12_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC3FA_2_LC_16_12_3  (
            .in0(N__39293),
            .in1(N__42770),
            .in2(N__39287),
            .in3(N__43523),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_375_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5KUTL_31_LC_16_12_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5KUTL_31_LC_16_12_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5KUTL_31_LC_16_12_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5KUTL_31_LC_16_12_4  (
            .in0(N__45802),
            .in1(N__39284),
            .in2(N__39272),
            .in3(N__39437),
            .lcout(\delay_measurement_inst.N_265_i ),
            .ltout(\delay_measurement_inst.N_265_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICTS5M_31_LC_16_12_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICTS5M_31_LC_16_12_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICTS5M_31_LC_16_12_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICTS5M_31_LC_16_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39269),
            .in3(N__46773),
            .lcout(\delay_measurement_inst.N_265_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_13_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_13_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39259),
            .lcout(\delay_measurement_inst.delay_tr_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4T357_15_LC_16_13_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4T357_15_LC_16_13_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4T357_15_LC_16_13_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4T357_15_LC_16_13_1  (
            .in0(N__45153),
            .in1(N__39536),
            .in2(_gnd_net_),
            .in3(N__43239),
            .lcout(\delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI43GB_6_LC_16_13_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI43GB_6_LC_16_13_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI43GB_6_LC_16_13_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI43GB_6_LC_16_13_2  (
            .in0(N__44761),
            .in1(N__44655),
            .in2(_gnd_net_),
            .in3(N__44715),
            .lcout(\delay_measurement_inst.N_410 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI9IAF_1_LC_16_13_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI9IAF_1_LC_16_13_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI9IAF_1_LC_16_13_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI9IAF_1_LC_16_13_3  (
            .in0(N__40138),
            .in1(N__44812),
            .in2(N__44601),
            .in3(N__44760),
            .lcout(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ5M42_2_LC_16_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ5M42_2_LC_16_13_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ5M42_2_LC_16_13_4 .LUT_INIT=16'b0001001100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ5M42_2_LC_16_13_4  (
            .in0(N__42797),
            .in1(N__44594),
            .in2(N__43403),
            .in3(N__42806),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_2_LC_16_13_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_2_LC_16_13_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_2_LC_16_13_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_2_LC_16_13_5  (
            .in0(N__39431),
            .in1(N__43619),
            .in2(N__39440),
            .in3(N__39413),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_364 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI86841_4_LC_16_13_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI86841_4_LC_16_13_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI86841_4_LC_16_13_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI86841_4_LC_16_13_7  (
            .in0(N__47780),
            .in1(N__44811),
            .in2(N__45160),
            .in3(N__44866),
            .lcout(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL5GJ7_15_LC_16_14_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL5GJ7_15_LC_16_14_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL5GJ7_15_LC_16_14_0 .LUT_INIT=16'b0000111100000010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL5GJ7_15_LC_16_14_0  (
            .in0(N__45155),
            .in1(N__42768),
            .in2(N__45801),
            .in3(N__43240),
            .lcout(\delay_measurement_inst.N_271_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO4MS_29_LC_16_14_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO4MS_29_LC_16_14_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO4MS_29_LC_16_14_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO4MS_29_LC_16_14_1  (
            .in0(_gnd_net_),
            .in1(N__45821),
            .in2(_gnd_net_),
            .in3(N__45875),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_16_14_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_16_14_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_16_14_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_16_14_2  (
            .in0(N__45317),
            .in1(N__45356),
            .in2(N__45935),
            .in3(N__45392),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_6_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_16_14_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_16_14_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_16_14_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_16_14_3  (
            .in0(N__45563),
            .in1(N__42812),
            .in2(N__39425),
            .in3(N__39422),
            .lcout(\delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20 ),
            .ltout(\delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI9DQM6_10_LC_16_14_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI9DQM6_10_LC_16_14_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI9DQM6_10_LC_16_14_4 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI9DQM6_10_LC_16_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39416),
            .in3(N__39535),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_409 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_16_14_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_16_14_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_16_14_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_16_14_5  (
            .in0(N__45277),
            .in1(N__44488),
            .in2(N__45235),
            .in3(N__44542),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_16_14_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_16_14_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_16_14_6 .LUT_INIT=16'b0001000101010001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_16_14_6  (
            .in0(N__45154),
            .in1(N__47782),
            .in2(N__39524),
            .in3(N__44602),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_400_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_16_14_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_16_14_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_16_14_7 .LUT_INIT=16'b1101110111011100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_16_14_7  (
            .in0(N__43241),
            .in1(N__45790),
            .in2(N__39521),
            .in3(N__42764),
            .lcout(\delay_measurement_inst.N_358 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_esr_9_LC_16_15_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_9_LC_16_15_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_9_LC_16_15_0 .LUT_INIT=16'b1100110011001101;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_9_LC_16_15_0  (
            .in0(N__39515),
            .in1(N__44603),
            .in2(N__45803),
            .in3(N__43541),
            .lcout(measured_delay_tr_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47257),
            .ce(N__43462),
            .sr(N__46643));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_16_15_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_16_15_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_16_15_1 .LUT_INIT=16'b0000000011110001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_16_15_1  (
            .in0(N__47783),
            .in1(N__45161),
            .in2(N__42769),
            .in3(N__43242),
            .lcout(\delay_measurement_inst.N_394_1 ),
            .ltout(\delay_measurement_inst.N_394_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_esr_10_LC_16_15_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_10_LC_16_15_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_10_LC_16_15_2 .LUT_INIT=16'b1111110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_10_LC_16_15_2  (
            .in0(_gnd_net_),
            .in1(N__45796),
            .in2(N__39518),
            .in3(N__44543),
            .lcout(measured_delay_tr_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47257),
            .ce(N__43462),
            .sr(N__46643));
    defparam \delay_measurement_inst.delay_tr_reg_esr_11_LC_16_15_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_11_LC_16_15_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_11_LC_16_15_3 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_11_LC_16_15_3  (
            .in0(N__45794),
            .in1(N__39512),
            .in2(_gnd_net_),
            .in3(N__44492),
            .lcout(measured_delay_tr_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47257),
            .ce(N__43462),
            .sr(N__46643));
    defparam \delay_measurement_inst.delay_tr_reg_esr_12_LC_16_15_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_12_LC_16_15_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_12_LC_16_15_4 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_12_LC_16_15_4  (
            .in0(N__39513),
            .in1(N__45797),
            .in2(_gnd_net_),
            .in3(N__45281),
            .lcout(measured_delay_tr_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47257),
            .ce(N__43462),
            .sr(N__46643));
    defparam \delay_measurement_inst.delay_tr_reg_esr_13_LC_16_15_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_13_LC_16_15_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_13_LC_16_15_5 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_13_LC_16_15_5  (
            .in0(N__45795),
            .in1(N__39514),
            .in2(_gnd_net_),
            .in3(N__45236),
            .lcout(measured_delay_tr_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47257),
            .ce(N__43462),
            .sr(N__46643));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0_6_LC_16_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0_6_LC_16_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0_6_LC_16_15_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0_6_LC_16_15_6  (
            .in0(N__39489),
            .in1(N__41520),
            .in2(N__41991),
            .in3(N__39462),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_esr_6_LC_16_16_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_6_LC_16_16_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_6_LC_16_16_0 .LUT_INIT=16'b0101111100010011;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_6_LC_16_16_0  (
            .in0(N__43544),
            .in1(N__43592),
            .in2(N__43648),
            .in3(N__44765),
            .lcout(measured_delay_tr_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47248),
            .ce(N__43461),
            .sr(N__46649));
    defparam \delay_measurement_inst.delay_tr_reg_ess_3_LC_16_16_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_ess_3_LC_16_16_1 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_tr_reg_ess_3_LC_16_16_1 .LUT_INIT=16'b1010100010100000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_ess_3_LC_16_16_1  (
            .in0(N__43401),
            .in1(N__43645),
            .in2(N__43602),
            .in3(N__43546),
            .lcout(measured_delay_tr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47248),
            .ce(N__43461),
            .sr(N__46649));
    defparam \delay_measurement_inst.delay_tr_reg_esr_5_LC_16_16_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_5_LC_16_16_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_5_LC_16_16_4 .LUT_INIT=16'b1111000010000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_5_LC_16_16_4  (
            .in0(N__43543),
            .in1(N__43646),
            .in2(N__44819),
            .in3(N__43591),
            .lcout(measured_delay_tr_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47248),
            .ce(N__43461),
            .sr(N__46649));
    defparam \delay_measurement_inst.delay_tr_reg_esr_19_LC_16_16_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_19_LC_16_16_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_19_LC_16_16_5 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_19_LC_16_16_5  (
            .in0(N__45785),
            .in1(N__44930),
            .in2(_gnd_net_),
            .in3(N__43253),
            .lcout(measured_delay_tr_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47248),
            .ce(N__43461),
            .sr(N__46649));
    defparam \delay_measurement_inst.delay_tr_reg_ess_1_LC_16_16_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_ess_1_LC_16_16_6 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_tr_reg_ess_1_LC_16_16_6 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_ess_1_LC_16_16_6  (
            .in0(N__43545),
            .in1(N__43593),
            .in2(N__43649),
            .in3(N__40139),
            .lcout(measured_delay_tr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47248),
            .ce(N__43461),
            .sr(N__46649));
    defparam \delay_measurement_inst.delay_tr_reg_esr_2_LC_16_16_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_2_LC_16_16_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_2_LC_16_16_7 .LUT_INIT=16'b1010100010100000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_2_LC_16_16_7  (
            .in0(N__42789),
            .in1(N__43638),
            .in2(N__43601),
            .in3(N__43542),
            .lcout(measured_delay_tr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47248),
            .ce(N__43461),
            .sr(N__46649));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_0_LC_16_17_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_0_LC_16_17_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_0_LC_16_17_0 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_0_LC_16_17_0  (
            .in0(N__39568),
            .in1(N__39719),
            .in2(N__40019),
            .in3(N__40065),
            .lcout(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47241),
            .ce(N__40518),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_1_LC_16_17_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_1_LC_16_17_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_1_LC_16_17_1 .LUT_INIT=16'b0000110001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_1_LC_16_17_1  (
            .in0(N__40066),
            .in1(N__40011),
            .in2(N__39738),
            .in3(N__39569),
            .lcout(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47241),
            .ce(N__40518),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_0_LC_16_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_0_LC_16_17_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_0_LC_16_17_4 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_0_LC_16_17_4  (
            .in0(N__48028),
            .in1(N__48155),
            .in2(N__43344),
            .in3(N__47894),
            .lcout(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47241),
            .ce(N__40518),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_1_LC_16_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_1_LC_16_17_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_1_LC_16_17_5 .LUT_INIT=16'b0000101000110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_1_LC_16_17_5  (
            .in0(N__48156),
            .in1(N__43334),
            .in2(N__47913),
            .in3(N__48029),
            .lcout(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47241),
            .ce(N__40518),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_16_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_16_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_16_17_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_16_17_6  (
            .in0(N__43333),
            .in1(N__43362),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.stoper_state_0_LC_16_17_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.stoper_state_0_LC_16_17_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_slave.stoper_hc.stoper_state_0_LC_16_17_7 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \phase_controller_slave.stoper_hc.stoper_state_0_LC_16_17_7  (
            .in0(N__41021),
            .in1(N__40579),
            .in2(N__40919),
            .in3(N__40728),
            .lcout(\phase_controller_slave.stoper_hc.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47241),
            .ce(N__40518),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.target_time_17_LC_16_18_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_17_LC_16_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_17_LC_16_18_0 .LUT_INIT=16'b0100010001010101;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_17_LC_16_18_0  (
            .in0(N__44181),
            .in1(N__42347),
            .in2(_gnd_net_),
            .in3(N__43893),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47232),
            .ce(N__43707),
            .sr(N__46667));
    defparam \phase_controller_slave.stoper_hc.target_time_8_LC_16_18_1 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_8_LC_16_18_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_8_LC_16_18_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_8_LC_16_18_1  (
            .in0(N__43896),
            .in1(N__44184),
            .in2(_gnd_net_),
            .in3(N__41767),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47232),
            .ce(N__43707),
            .sr(N__46667));
    defparam \phase_controller_slave.stoper_hc.target_time_16_LC_16_18_2 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_16_LC_16_18_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_16_LC_16_18_2 .LUT_INIT=16'b0100010001010101;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_16_LC_16_18_2  (
            .in0(N__44180),
            .in1(N__40454),
            .in2(_gnd_net_),
            .in3(N__43892),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47232),
            .ce(N__43707),
            .sr(N__46667));
    defparam \phase_controller_slave.stoper_hc.target_time_18_LC_16_18_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_18_LC_16_18_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_18_LC_16_18_3 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_18_LC_16_18_3  (
            .in0(N__43894),
            .in1(N__44182),
            .in2(_gnd_net_),
            .in3(N__42190),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47232),
            .ce(N__43707),
            .sr(N__46667));
    defparam \phase_controller_slave.stoper_hc.target_time_19_LC_16_18_6 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_19_LC_16_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_19_LC_16_18_6 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_19_LC_16_18_6  (
            .in0(N__44179),
            .in1(N__40394),
            .in2(_gnd_net_),
            .in3(N__41888),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47232),
            .ce(N__43707),
            .sr(N__46667));
    defparam \phase_controller_slave.stoper_hc.target_time_1_LC_16_18_7 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_1_LC_16_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_1_LC_16_18_7 .LUT_INIT=16'b1111111110101000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_1_LC_16_18_7  (
            .in0(N__43895),
            .in1(N__40342),
            .in2(N__41275),
            .in3(N__44183),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47232),
            .ce(N__43707),
            .sr(N__46667));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_16_19_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_16_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_16_19_0  (
            .in0(_gnd_net_),
            .in1(N__41192),
            .in2(N__41201),
            .in3(N__45660),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_16_19_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_16_19_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_16_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_16_19_1  (
            .in0(_gnd_net_),
            .in1(N__41186),
            .in2(N__41180),
            .in3(N__45643),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_16_19_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_16_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_16_19_2  (
            .in0(_gnd_net_),
            .in1(N__41156),
            .in2(N__41171),
            .in3(N__45610),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_16_19_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_16_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_16_19_3  (
            .in0(_gnd_net_),
            .in1(N__41138),
            .in2(N__41150),
            .in3(N__46111),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_16_19_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_16_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_16_19_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_16_19_4  (
            .in0(_gnd_net_),
            .in1(N__41117),
            .in2(N__41132),
            .in3(N__46090),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_16_19_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_16_19_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_16_19_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_16_19_5  (
            .in0(_gnd_net_),
            .in1(N__41096),
            .in2(N__41111),
            .in3(N__46069),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_16_19_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_16_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_16_19_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_16_19_6  (
            .in0(N__46048),
            .in1(N__41075),
            .in2(N__41090),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_16_19_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_16_19_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_16_19_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_16_19_7  (
            .in0(N__46027),
            .in1(N__41369),
            .in2(N__41381),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_16_20_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_16_20_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_16_20_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_16_20_0  (
            .in0(_gnd_net_),
            .in1(N__41363),
            .in2(N__47363),
            .in3(N__48214),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_16_20_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_16_20_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_16_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_16_20_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_16_20_1  (
            .in0(N__46003),
            .in1(N__41339),
            .in2(N__41357),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_16_20_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_16_20_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_16_20_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_16_20_2  (
            .in0(_gnd_net_),
            .in1(N__41333),
            .in2(N__41504),
            .in3(N__45982),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_16_20_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_16_20_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_16_20_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_16_20_3  (
            .in0(_gnd_net_),
            .in1(N__41309),
            .in2(N__41327),
            .in3(N__46291),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_16_20_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_16_20_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_16_20_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_16_20_4  (
            .in0(_gnd_net_),
            .in1(N__41303),
            .in2(N__41966),
            .in3(N__46270),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_16_20_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_16_20_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_16_20_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_16_20_5  (
            .in0(_gnd_net_),
            .in1(N__41288),
            .in2(N__41297),
            .in3(N__46249),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_16_20_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_16_20_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_16_20_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_16_20_6  (
            .in0(N__46225),
            .in1(N__41282),
            .in2(N__41393),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_16_20_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_16_20_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_16_20_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_16_20_7  (
            .in0(_gnd_net_),
            .in1(N__41624),
            .in2(N__44357),
            .in3(N__46202),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_16_21_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_16_21_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_16_21_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_16_21_0  (
            .in0(_gnd_net_),
            .in1(N__41606),
            .in2(N__41618),
            .in3(N__46177),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_16_21_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_16_21_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_16_21_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_16_21_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_16_21_1  (
            .in0(_gnd_net_),
            .in1(N__41600),
            .in2(N__41585),
            .in3(N__46156),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_16_21_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_16_21_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_16_21_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_16_21_2  (
            .in0(_gnd_net_),
            .in1(N__41594),
            .in2(N__41540),
            .in3(N__46135),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_16_21_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_16_21_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_16_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_16_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41588),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_16_21_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_16_21_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_16_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_18_LC_16_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43210),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47219),
            .ce(N__46856),
            .sr(N__46691));
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_16_21_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_16_21_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_16_21_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_19_LC_16_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41567),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47219),
            .ce(N__46856),
            .sr(N__46691));
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_16_22_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_16_22_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_16_22_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_11_LC_16_22_0  (
            .in0(N__47593),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41527),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47214),
            .ce(N__46859),
            .sr(N__46702));
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_16_22_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_16_22_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_16_22_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_15_LC_16_22_3  (
            .in0(_gnd_net_),
            .in1(N__41491),
            .in2(_gnd_net_),
            .in3(N__47538),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47214),
            .ce(N__46859),
            .sr(N__46702));
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_16_22_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_16_22_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_16_22_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_13_LC_16_22_4  (
            .in0(N__47594),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41998),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47214),
            .ce(N__46859),
            .sr(N__46702));
    defparam SB_DFF_inst_DELAY_HC1_LC_17_5_2.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_HC1_LC_17_5_2.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_HC1_LC_17_5_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_DELAY_HC1_LC_17_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41954),
            .lcout(delay_hc_d1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47343),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_DELAY_HC2_LC_17_5_6.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_HC2_LC_17_5_6.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_HC2_LC_17_5_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_DELAY_HC2_LC_17_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41945),
            .lcout(delay_hc_d2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47343),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_LC_17_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_LC_17_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_LC_17_7_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_LC_17_7_0  (
            .in0(N__41809),
            .in1(N__44291),
            .in2(N__42275),
            .in3(N__41894),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_25_LC_17_7_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_25_LC_17_7_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_25_LC_17_7_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_25_LC_17_7_2  (
            .in0(N__42466),
            .in1(N__41837),
            .in2(_gnd_net_),
            .in3(N__42559),
            .lcout(measured_delay_hc_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47335),
            .ce(),
            .sr(N__46595));
    defparam \delay_measurement_inst.delay_hc_reg_26_LC_17_7_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_26_LC_17_7_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_26_LC_17_7_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_26_LC_17_7_3  (
            .in0(N__42560),
            .in1(N__41825),
            .in2(_gnd_net_),
            .in3(N__42467),
            .lcout(measured_delay_hc_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47335),
            .ce(),
            .sr(N__46595));
    defparam \delay_measurement_inst.delay_hc_reg_23_LC_17_7_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_23_LC_17_7_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_23_LC_17_7_4 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_23_LC_17_7_4  (
            .in0(N__42465),
            .in1(_gnd_net_),
            .in2(N__41813),
            .in3(N__42558),
            .lcout(measured_delay_hc_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47335),
            .ce(),
            .sr(N__46595));
    defparam \delay_measurement_inst.delay_hc_reg_8_LC_17_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_8_LC_17_8_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_8_LC_17_8_0 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_8_LC_17_8_0  (
            .in0(N__42104),
            .in1(N__41740),
            .in2(N__42651),
            .in3(N__41801),
            .lcout(measured_delay_hc_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47329),
            .ce(),
            .sr(N__46599));
    defparam \delay_measurement_inst.delay_hc_reg_7_LC_17_8_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_7_LC_17_8_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_7_LC_17_8_3 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_7_LC_17_8_3  (
            .in0(N__41648),
            .in1(N__42632),
            .in2(N__41708),
            .in3(N__42103),
            .lcout(measured_delay_hc_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47329),
            .ce(),
            .sr(N__46599));
    defparam \delay_measurement_inst.delay_hc_reg_24_LC_17_8_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_24_LC_17_8_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_24_LC_17_8_5 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_24_LC_17_8_5  (
            .in0(N__42446),
            .in1(N__42274),
            .in2(_gnd_net_),
            .in3(N__42630),
            .lcout(measured_delay_hc_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47329),
            .ce(),
            .sr(N__46599));
    defparam \delay_measurement_inst.delay_hc_reg_0_LC_17_8_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_0_LC_17_8_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_0_LC_17_8_6 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_0_LC_17_8_6  (
            .in0(N__42629),
            .in1(N__42233),
            .in2(_gnd_net_),
            .in3(N__42444),
            .lcout(measured_delay_hc_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47329),
            .ce(),
            .sr(N__46599));
    defparam \delay_measurement_inst.delay_hc_reg_18_LC_17_8_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_18_LC_17_8_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_18_LC_17_8_7 .LUT_INIT=16'b1111111010111010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_18_LC_17_8_7  (
            .in0(N__42445),
            .in1(N__42631),
            .in2(N__42181),
            .in3(N__42209),
            .lcout(measured_delay_hc_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47329),
            .ce(),
            .sr(N__46599));
    defparam \delay_measurement_inst.delay_hc_reg_30_LC_17_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_30_LC_17_9_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_30_LC_17_9_0 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_30_LC_17_9_0  (
            .in0(N__42441),
            .in1(_gnd_net_),
            .in2(N__42653),
            .in3(N__44317),
            .lcout(measured_delay_hc_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47321),
            .ce(),
            .sr(N__46602));
    defparam \delay_measurement_inst.delay_hc_reg_29_LC_17_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_29_LC_17_9_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_29_LC_17_9_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_29_LC_17_9_1  (
            .in0(N__44342),
            .in1(N__42640),
            .in2(_gnd_net_),
            .in3(N__42440),
            .lcout(measured_delay_hc_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47321),
            .ce(),
            .sr(N__46602));
    defparam \delay_measurement_inst.delay_hc_reg_19_LC_17_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_19_LC_17_9_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_19_LC_17_9_3 .LUT_INIT=16'b1110001011111111;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_19_LC_17_9_3  (
            .in0(N__42048),
            .in1(N__42644),
            .in2(N__42134),
            .in3(N__42093),
            .lcout(measured_delay_hc_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47321),
            .ce(),
            .sr(N__46602));
    defparam \delay_measurement_inst.delay_hc_reg_28_LC_17_9_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_28_LC_17_9_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_28_LC_17_9_4 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_28_LC_17_9_4  (
            .in0(N__42439),
            .in1(_gnd_net_),
            .in2(N__42652),
            .in3(N__44330),
            .lcout(measured_delay_hc_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47321),
            .ce(),
            .sr(N__46602));
    defparam \delay_measurement_inst.delay_hc_reg_27_LC_17_9_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_27_LC_17_9_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_27_LC_17_9_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_27_LC_17_9_5  (
            .in0(N__44303),
            .in1(N__42636),
            .in2(_gnd_net_),
            .in3(N__42438),
            .lcout(measured_delay_hc_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47321),
            .ce(),
            .sr(N__46602));
    defparam \delay_measurement_inst.delay_hc_reg_21_LC_17_10_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_21_LC_17_10_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_21_LC_17_10_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_21_LC_17_10_1  (
            .in0(N__42013),
            .in1(N__42645),
            .in2(_gnd_net_),
            .in3(N__42463),
            .lcout(measured_delay_hc_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47313),
            .ce(),
            .sr(N__46607));
    defparam \delay_measurement_inst.delay_hc_reg_22_LC_17_10_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_22_LC_17_10_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_22_LC_17_10_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_22_LC_17_10_3  (
            .in0(N__42667),
            .in1(N__42646),
            .in2(_gnd_net_),
            .in3(N__42464),
            .lcout(measured_delay_hc_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47313),
            .ce(),
            .sr(N__46607));
    defparam \delay_measurement_inst.delay_hc_reg_17_LC_17_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_17_LC_17_10_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_17_LC_17_10_5 .LUT_INIT=16'b1111111111100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_17_LC_17_10_5  (
            .in0(N__42329),
            .in1(N__42647),
            .in2(N__42491),
            .in3(N__42462),
            .lcout(measured_delay_hc_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47313),
            .ce(),
            .sr(N__46607));
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_11_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_11_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_11_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_11_0  (
            .in0(N__42980),
            .in1(N__43419),
            .in2(_gnd_net_),
            .in3(N__42296),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_17_11_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .clk(N__47301),
            .ce(N__42857),
            .sr(N__46612));
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_11_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_11_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_11_1  (
            .in0(N__42961),
            .in1(N__44889),
            .in2(_gnd_net_),
            .in3(N__42293),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .clk(N__47301),
            .ce(N__42857),
            .sr(N__46612));
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_11_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_11_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_11_2  (
            .in0(N__42981),
            .in1(N__44835),
            .in2(_gnd_net_),
            .in3(N__42290),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .clk(N__47301),
            .ce(N__42857),
            .sr(N__46612));
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_11_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_11_3  (
            .in0(N__42962),
            .in1(N__44781),
            .in2(_gnd_net_),
            .in3(N__42287),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .clk(N__47301),
            .ce(N__42857),
            .sr(N__46612));
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_11_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_11_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_11_4  (
            .in0(N__42982),
            .in1(N__44731),
            .in2(_gnd_net_),
            .in3(N__42284),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .clk(N__47301),
            .ce(N__42857),
            .sr(N__46612));
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_11_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_11_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_11_5  (
            .in0(N__42963),
            .in1(N__44677),
            .in2(_gnd_net_),
            .in3(N__42281),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .clk(N__47301),
            .ce(N__42857),
            .sr(N__46612));
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_11_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_11_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_11_6  (
            .in0(N__42983),
            .in1(N__44625),
            .in2(_gnd_net_),
            .in3(N__42278),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .clk(N__47301),
            .ce(N__42857),
            .sr(N__46612));
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_11_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_11_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_11_7  (
            .in0(N__42964),
            .in1(N__44557),
            .in2(_gnd_net_),
            .in3(N__42710),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .clk(N__47301),
            .ce(N__42857),
            .sr(N__46612));
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_12_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_12_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_12_0  (
            .in0(N__42956),
            .in1(N__44511),
            .in2(_gnd_net_),
            .in3(N__42707),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_17_12_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .clk(N__47292),
            .ce(N__42856),
            .sr(N__46616));
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_12_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_12_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_12_1  (
            .in0(N__42968),
            .in1(N__45298),
            .in2(_gnd_net_),
            .in3(N__42704),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .clk(N__47292),
            .ce(N__42856),
            .sr(N__46616));
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_12_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_12_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_12_2  (
            .in0(N__42953),
            .in1(N__45252),
            .in2(_gnd_net_),
            .in3(N__42701),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .clk(N__47292),
            .ce(N__42856),
            .sr(N__46616));
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_12_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_12_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_12_3  (
            .in0(N__42965),
            .in1(N__45201),
            .in2(_gnd_net_),
            .in3(N__42698),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .clk(N__47292),
            .ce(N__42856),
            .sr(N__46616));
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_12_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_12_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_12_4  (
            .in0(N__42954),
            .in1(N__45175),
            .in2(_gnd_net_),
            .in3(N__42695),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .clk(N__47292),
            .ce(N__42856),
            .sr(N__46616));
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_12_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_12_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_12_5  (
            .in0(N__42966),
            .in1(N__45094),
            .in2(_gnd_net_),
            .in3(N__42692),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .clk(N__47292),
            .ce(N__42856),
            .sr(N__46616));
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_12_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_12_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_12_6  (
            .in0(N__42955),
            .in1(N__45051),
            .in2(_gnd_net_),
            .in3(N__42689),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .clk(N__47292),
            .ce(N__42856),
            .sr(N__46616));
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_12_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_12_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_12_7  (
            .in0(N__42967),
            .in1(N__44992),
            .in2(_gnd_net_),
            .in3(N__42686),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .clk(N__47292),
            .ce(N__42856),
            .sr(N__46616));
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_13_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_13_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_13_0  (
            .in0(N__42945),
            .in1(N__44949),
            .in2(_gnd_net_),
            .in3(N__42737),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_17_13_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .clk(N__47284),
            .ce(N__42849),
            .sr(N__46619));
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_13_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_13_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_13_1  (
            .in0(N__42949),
            .in1(N__45583),
            .in2(_gnd_net_),
            .in3(N__42734),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .clk(N__47284),
            .ce(N__42849),
            .sr(N__46619));
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_13_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_13_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_13_2  (
            .in0(N__42946),
            .in1(N__45537),
            .in2(_gnd_net_),
            .in3(N__42731),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .clk(N__47284),
            .ce(N__42849),
            .sr(N__46619));
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_13_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_13_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_13_3  (
            .in0(N__42950),
            .in1(N__45504),
            .in2(_gnd_net_),
            .in3(N__42728),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .clk(N__47284),
            .ce(N__42849),
            .sr(N__46619));
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_13_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_13_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_13_4  (
            .in0(N__42947),
            .in1(N__45471),
            .in2(_gnd_net_),
            .in3(N__42725),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .clk(N__47284),
            .ce(N__42849),
            .sr(N__46619));
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_13_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_13_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_13_5  (
            .in0(N__42951),
            .in1(N__45438),
            .in2(_gnd_net_),
            .in3(N__42722),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .clk(N__47284),
            .ce(N__42849),
            .sr(N__46619));
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_13_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_13_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_13_6  (
            .in0(N__42948),
            .in1(N__45408),
            .in2(_gnd_net_),
            .in3(N__42719),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .clk(N__47284),
            .ce(N__42849),
            .sr(N__46619));
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_13_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_13_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_13_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_13_7  (
            .in0(N__42952),
            .in1(N__45370),
            .in2(_gnd_net_),
            .in3(N__42716),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .clk(N__47284),
            .ce(N__42849),
            .sr(N__46619));
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_14_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_14_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_14_0  (
            .in0(N__42957),
            .in1(N__45336),
            .in2(_gnd_net_),
            .in3(N__42713),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_17_14_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .clk(N__47277),
            .ce(N__42839),
            .sr(N__46631));
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_14_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_14_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_14_1  (
            .in0(N__42969),
            .in1(N__45954),
            .in2(_gnd_net_),
            .in3(N__42995),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .clk(N__47277),
            .ce(N__42839),
            .sr(N__46631));
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_14_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_14_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_14_2  (
            .in0(N__42958),
            .in1(N__45891),
            .in2(_gnd_net_),
            .in3(N__42992),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .clk(N__47277),
            .ce(N__42839),
            .sr(N__46631));
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_14_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_14_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_14_3  (
            .in0(N__42970),
            .in1(N__45837),
            .in2(_gnd_net_),
            .in3(N__42989),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .clk(N__47277),
            .ce(N__42839),
            .sr(N__46631));
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_14_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_14_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_14_4  (
            .in0(N__42959),
            .in1(N__45913),
            .in2(_gnd_net_),
            .in3(N__42986),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ),
            .clk(N__47277),
            .ce(N__42839),
            .sr(N__46631));
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_14_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_14_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_14_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_14_5  (
            .in0(N__45859),
            .in1(N__42960),
            .in2(_gnd_net_),
            .in3(N__42860),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47277),
            .ce(N__42839),
            .sr(N__46631));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_17_15_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_17_15_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_17_15_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_17_15_0  (
            .in0(N__45455),
            .in1(N__45488),
            .in2(N__45422),
            .in3(N__45515),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_7_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_0_16_LC_17_15_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_0_16_LC_17_15_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_0_16_LC_17_15_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_0_16_LC_17_15_3  (
            .in0(N__44973),
            .in1(N__45024),
            .in2(N__44925),
            .in3(N__45075),
            .lcout(\delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_17_15_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_17_15_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_17_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_17_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44897),
            .lcout(\delay_measurement_inst.elapsed_time_tr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47265),
            .ce(N__45725),
            .sr(N__46636));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_17_15_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_17_15_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_17_15_6 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_17_15_6  (
            .in0(N__45076),
            .in1(N__44974),
            .in2(N__44926),
            .in3(N__45025),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_esr_16_LC_17_16_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_16_LC_17_16_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_16_LC_17_16_1 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_16_LC_17_16_1  (
            .in0(N__45080),
            .in1(N__45760),
            .in2(_gnd_net_),
            .in3(N__43254),
            .lcout(measured_delay_tr_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47258),
            .ce(N__43463),
            .sr(N__46644));
    defparam \delay_measurement_inst.delay_tr_reg_esr_17_LC_17_16_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_17_LC_17_16_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_17_LC_17_16_2 .LUT_INIT=16'b1111111100001010;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_17_LC_17_16_2  (
            .in0(N__43255),
            .in1(_gnd_net_),
            .in2(N__45786),
            .in3(N__45029),
            .lcout(measured_delay_tr_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47258),
            .ce(N__43463),
            .sr(N__46644));
    defparam \delay_measurement_inst.delay_tr_reg_esr_18_LC_17_16_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_18_LC_17_16_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_18_LC_17_16_3 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_18_LC_17_16_3  (
            .in0(N__44978),
            .in1(N__45761),
            .in2(_gnd_net_),
            .in3(N__43256),
            .lcout(measured_delay_tr_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47258),
            .ce(N__43463),
            .sr(N__46644));
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_17_17_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_17_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_17_17_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.state_RNI7NN7_0_LC_17_17_0  (
            .in0(_gnd_net_),
            .in1(N__43050),
            .in2(_gnd_net_),
            .in3(N__43003),
            .lcout(\phase_controller_inst1.N_83 ),
            .ltout(\phase_controller_inst1.N_83_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_tr_LC_17_17_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_LC_17_17_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_tr_LC_17_17_1 .LUT_INIT=16'b1111111100000010;
    LogicCell40 \phase_controller_inst1.start_timer_tr_LC_17_17_1  (
            .in0(N__48157),
            .in1(N__43160),
            .in2(N__43127),
            .in3(N__43124),
            .lcout(\phase_controller_inst1.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47249),
            .ce(),
            .sr(N__46650));
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_17_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_17_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_17_17_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_17_17_2  (
            .in0(N__48158),
            .in1(N__47998),
            .in2(_gnd_net_),
            .in3(N__47873),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_17_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_17_17_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_17_17_3 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_LC_17_17_3  (
            .in0(N__43054),
            .in1(N__43366),
            .in2(N__43103),
            .in3(N__43346),
            .lcout(\phase_controller_inst1.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47249),
            .ce(),
            .sr(N__46650));
    defparam \phase_controller_inst1.state_0_LC_17_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_0_LC_17_17_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_0_LC_17_17_5 .LUT_INIT=16'b1100111000001010;
    LogicCell40 \phase_controller_inst1.state_0_LC_17_17_5  (
            .in0(N__43004),
            .in1(N__43096),
            .in2(N__43055),
            .in3(N__43040),
            .lcout(\phase_controller_inst1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47249),
            .ce(),
            .sr(N__46650));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_17_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_17_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_17_17_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_17_17_6  (
            .in0(_gnd_net_),
            .in1(N__47997),
            .in2(_gnd_net_),
            .in3(N__47872),
            .lcout(\phase_controller_inst1.stoper_tr.time_passed11 ),
            .ltout(\phase_controller_inst1.stoper_tr.time_passed11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_17_17_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_17_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_17_17_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_17_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43301),
            .in3(N__43345),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_17_18_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_17_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_17_18_0 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_17_18_0  (
            .in0(N__47889),
            .in1(N__48154),
            .in2(N__48066),
            .in3(N__46016),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47242),
            .ce(),
            .sr(N__46659));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_17_18_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_17_18_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_17_18_1 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_17_18_1  (
            .in0(N__48024),
            .in1(N__47890),
            .in2(N__48179),
            .in3(N__46187),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47242),
            .ce(),
            .sr(N__46659));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_17_18_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_17_18_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_17_18_2 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_17_18_2  (
            .in0(N__47888),
            .in1(N__48153),
            .in2(N__48065),
            .in3(N__46037),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47242),
            .ce(),
            .sr(N__46659));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_17_18_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_17_18_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_17_18_3 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_17_18_3  (
            .in0(N__48025),
            .in1(N__47891),
            .in2(N__48180),
            .in3(N__45632),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47242),
            .ce(),
            .sr(N__46659));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_17_18_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_17_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_17_18_4 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_17_18_4  (
            .in0(N__47886),
            .in1(N__48145),
            .in2(N__48063),
            .in3(N__45599),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47242),
            .ce(),
            .sr(N__46659));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_17_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_17_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_17_18_5 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_17_18_5  (
            .in0(N__48026),
            .in1(N__47892),
            .in2(N__48181),
            .in3(N__46100),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47242),
            .ce(),
            .sr(N__46659));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_17_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_17_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_17_18_6 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_17_18_6  (
            .in0(N__47887),
            .in1(N__48149),
            .in2(N__48064),
            .in3(N__46079),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47242),
            .ce(),
            .sr(N__46659));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_17_18_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_17_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_17_18_7 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_17_18_7  (
            .in0(N__48027),
            .in1(N__47893),
            .in2(N__48182),
            .in3(N__46058),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47242),
            .ce(),
            .sr(N__46659));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_17_19_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_17_19_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_17_19_0 .LUT_INIT=16'b1100100010001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_17_19_0  (
            .in0(N__47910),
            .in1(N__45992),
            .in2(N__48071),
            .in3(N__48173),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47233),
            .ce(),
            .sr(N__46668));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_17_19_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_17_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_17_19_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_17_19_1  (
            .in0(N__43367),
            .in1(N__45664),
            .in2(_gnd_net_),
            .in3(N__43343),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_17_19_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_17_19_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_17_19_2 .LUT_INIT=16'b1110000011010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_17_19_2  (
            .in0(N__48047),
            .in1(N__47933),
            .in2(N__43304),
            .in3(N__48178),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47233),
            .ce(),
            .sr(N__46668));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_17_19_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_17_19_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_17_19_3 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_17_19_3  (
            .in0(N__48174),
            .in1(N__48048),
            .in2(N__47946),
            .in3(N__45971),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47233),
            .ce(),
            .sr(N__46668));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_17_19_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_17_19_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_17_19_4 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_17_19_4  (
            .in0(N__47911),
            .in1(N__48175),
            .in2(N__48072),
            .in3(N__46280),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47233),
            .ce(),
            .sr(N__46668));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_17_19_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_17_19_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_17_19_5 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_17_19_5  (
            .in0(N__48176),
            .in1(N__48049),
            .in2(N__47947),
            .in3(N__46259),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47233),
            .ce(),
            .sr(N__46668));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_17_19_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_17_19_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_17_19_6 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_17_19_6  (
            .in0(N__47912),
            .in1(N__48177),
            .in2(N__48073),
            .in3(N__46238),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47233),
            .ce(),
            .sr(N__46668));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_17_20_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_17_20_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_17_20_0 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_17_20_0  (
            .in0(N__48059),
            .in1(N__48185),
            .in2(N__47948),
            .in3(N__46214),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47227),
            .ce(),
            .sr(N__46677));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_17_20_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_17_20_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_17_20_3 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_17_20_3  (
            .in0(N__47942),
            .in1(N__48061),
            .in2(N__48197),
            .in3(N__46121),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47227),
            .ce(),
            .sr(N__46677));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_17_20_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_17_20_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_17_20_5 .LUT_INIT=16'b1100100010001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_17_20_5  (
            .in0(N__47940),
            .in1(N__46166),
            .in2(N__48195),
            .in3(N__48062),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47227),
            .ce(),
            .sr(N__46677));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_17_20_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_17_20_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_17_20_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_17_20_7  (
            .in0(N__47941),
            .in1(N__48060),
            .in2(N__48196),
            .in3(N__46145),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47227),
            .ce(),
            .sr(N__46677));
    defparam \phase_controller_slave.stoper_tr.target_time_16_LC_17_21_0 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_tr.target_time_16_LC_17_21_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_tr.target_time_16_LC_17_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_slave.stoper_tr.target_time_16_LC_17_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44384),
            .lcout(\phase_controller_slave.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47224),
            .ce(N__44453),
            .sr(N__46682));
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_17_22_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_17_22_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_17_22_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_16_LC_17_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44385),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47220),
            .ce(N__46852),
            .sr(N__46692));
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_4_LC_18_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_4_LC_18_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_4_LC_18_9_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_4_LC_18_9_1  (
            .in0(N__44341),
            .in1(N__44329),
            .in2(N__44318),
            .in3(N__44302),
            .lcout(\phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_slave.stoper_hc.target_time_13_LC_18_10_3 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_13_LC_18_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_13_LC_18_10_3 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_13_LC_18_10_3  (
            .in0(N__44154),
            .in1(N__44282),
            .in2(_gnd_net_),
            .in3(N__43897),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47322),
            .ce(N__43712),
            .sr(N__46603));
    defparam \phase_controller_slave.stoper_hc.target_time_5_LC_18_11_5 .C_ON=1'b0;
    defparam \phase_controller_slave.stoper_hc.target_time_5_LC_18_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_slave.stoper_hc.target_time_5_LC_18_11_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_slave.stoper_hc.target_time_5_LC_18_11_5  (
            .in0(N__44156),
            .in1(N__43957),
            .in2(_gnd_net_),
            .in3(N__43827),
            .lcout(\phase_controller_slave.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47314),
            .ce(N__43711),
            .sr(N__46608));
    defparam \delay_measurement_inst.delay_tr_reg_esr_4_LC_18_12_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_4_LC_18_12_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_4_LC_18_12_6 .LUT_INIT=16'b1010100010100000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_4_LC_18_12_6  (
            .in0(N__44865),
            .in1(N__43647),
            .in2(N__43604),
            .in3(N__43550),
            .lcout(measured_delay_tr_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47302),
            .ce(N__43451),
            .sr(N__46613));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_18_13_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_18_13_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_18_13_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_18_13_0  (
            .in0(_gnd_net_),
            .in1(N__43424),
            .in2(N__44842),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.elapsed_time_tr_3 ),
            .ltout(),
            .carryin(bfn_18_13_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__47293),
            .ce(N__45703),
            .sr(N__46617));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_18_13_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_18_13_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_18_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_18_13_1  (
            .in0(_gnd_net_),
            .in1(N__44893),
            .in2(N__44788),
            .in3(N__44846),
            .lcout(\delay_measurement_inst.elapsed_time_tr_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__47293),
            .ce(N__45703),
            .sr(N__46617));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_18_13_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_18_13_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_18_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_18_13_2  (
            .in0(_gnd_net_),
            .in1(N__44737),
            .in2(N__44843),
            .in3(N__44792),
            .lcout(\delay_measurement_inst.elapsed_time_tr_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__47293),
            .ce(N__45703),
            .sr(N__46617));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_18_13_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_18_13_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_18_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_18_13_3  (
            .in0(_gnd_net_),
            .in1(N__44683),
            .in2(N__44789),
            .in3(N__44741),
            .lcout(\delay_measurement_inst.elapsed_time_tr_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__47293),
            .ce(N__45703),
            .sr(N__46617));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_18_13_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_18_13_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_18_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_18_13_4  (
            .in0(_gnd_net_),
            .in1(N__44738),
            .in2(N__44633),
            .in3(N__44687),
            .lcout(\delay_measurement_inst.elapsed_time_tr_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__47293),
            .ce(N__45703),
            .sr(N__46617));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_18_13_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_18_13_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_18_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_18_13_5  (
            .in0(_gnd_net_),
            .in1(N__44684),
            .in2(N__44569),
            .in3(N__44636),
            .lcout(\delay_measurement_inst.elapsed_time_tr_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__47293),
            .ce(N__45703),
            .sr(N__46617));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_18_13_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_18_13_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_18_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_18_13_6  (
            .in0(_gnd_net_),
            .in1(N__44629),
            .in2(N__44515),
            .in3(N__44573),
            .lcout(\delay_measurement_inst.elapsed_time_tr_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__47293),
            .ce(N__45703),
            .sr(N__46617));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_18_13_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_18_13_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_18_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_18_13_7  (
            .in0(_gnd_net_),
            .in1(N__45297),
            .in2(N__44570),
            .in3(N__44519),
            .lcout(\delay_measurement_inst.elapsed_time_tr_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__47293),
            .ce(N__45703),
            .sr(N__46617));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_18_14_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_18_14_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_18_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_18_14_0  (
            .in0(_gnd_net_),
            .in1(N__44516),
            .in2(N__45259),
            .in3(N__44474),
            .lcout(\delay_measurement_inst.elapsed_time_tr_11 ),
            .ltout(),
            .carryin(bfn_18_14_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__47285),
            .ce(N__45727),
            .sr(N__46620));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_18_14_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_18_14_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_18_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_18_14_1  (
            .in0(_gnd_net_),
            .in1(N__45302),
            .in2(N__45208),
            .in3(N__45263),
            .lcout(\delay_measurement_inst.elapsed_time_tr_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__47285),
            .ce(N__45727),
            .sr(N__46620));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_18_14_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_18_14_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_18_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_18_14_2  (
            .in0(_gnd_net_),
            .in1(N__45181),
            .in2(N__45260),
            .in3(N__45212),
            .lcout(\delay_measurement_inst.elapsed_time_tr_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__47285),
            .ce(N__45727),
            .sr(N__46620));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_18_14_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_18_14_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_18_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_18_14_3  (
            .in0(_gnd_net_),
            .in1(N__45100),
            .in2(N__45209),
            .in3(N__45185),
            .lcout(\delay_measurement_inst.elapsed_time_tr_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__47285),
            .ce(N__45727),
            .sr(N__46620));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_18_14_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_18_14_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_18_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_18_14_4  (
            .in0(_gnd_net_),
            .in1(N__45182),
            .in2(N__45059),
            .in3(N__45104),
            .lcout(\delay_measurement_inst.elapsed_time_tr_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__47285),
            .ce(N__45727),
            .sr(N__46620));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_18_14_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_18_14_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_18_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_18_14_5  (
            .in0(_gnd_net_),
            .in1(N__45101),
            .in2(N__45004),
            .in3(N__45062),
            .lcout(\delay_measurement_inst.elapsed_time_tr_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__47285),
            .ce(N__45727),
            .sr(N__46620));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_18_14_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_18_14_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_18_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_18_14_6  (
            .in0(_gnd_net_),
            .in1(N__45055),
            .in2(N__44953),
            .in3(N__45008),
            .lcout(\delay_measurement_inst.elapsed_time_tr_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__47285),
            .ce(N__45727),
            .sr(N__46620));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_18_14_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_18_14_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_18_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_18_14_7  (
            .in0(_gnd_net_),
            .in1(N__45579),
            .in2(N__45005),
            .in3(N__44960),
            .lcout(\delay_measurement_inst.elapsed_time_tr_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__47285),
            .ce(N__45727),
            .sr(N__46620));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_18_15_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_18_15_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_18_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_18_15_0  (
            .in0(_gnd_net_),
            .in1(N__44957),
            .in2(N__45548),
            .in3(N__44900),
            .lcout(\delay_measurement_inst.elapsed_time_tr_19 ),
            .ltout(),
            .carryin(bfn_18_15_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__47278),
            .ce(N__45726),
            .sr(N__46632));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_18_15_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_18_15_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_18_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_18_15_1  (
            .in0(_gnd_net_),
            .in1(N__45505),
            .in2(N__45590),
            .in3(N__45551),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__47278),
            .ce(N__45726),
            .sr(N__46632));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_18_15_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_18_15_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_18_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_18_15_2  (
            .in0(_gnd_net_),
            .in1(N__45547),
            .in2(N__45478),
            .in3(N__45509),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__47278),
            .ce(N__45726),
            .sr(N__46632));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_18_15_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_18_15_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_18_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_18_15_3  (
            .in0(_gnd_net_),
            .in1(N__45506),
            .in2(N__45445),
            .in3(N__45482),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__47278),
            .ce(N__45726),
            .sr(N__46632));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_18_15_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_18_15_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_18_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_18_15_4  (
            .in0(_gnd_net_),
            .in1(N__45409),
            .in2(N__45479),
            .in3(N__45449),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__47278),
            .ce(N__45726),
            .sr(N__46632));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_18_15_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_18_15_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_18_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_18_15_5  (
            .in0(_gnd_net_),
            .in1(N__45376),
            .in2(N__45446),
            .in3(N__45413),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__47278),
            .ce(N__45726),
            .sr(N__46632));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_18_15_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_18_15_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_18_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_18_15_6  (
            .in0(_gnd_net_),
            .in1(N__45410),
            .in2(N__45340),
            .in3(N__45380),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__47278),
            .ce(N__45726),
            .sr(N__46632));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_18_15_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_18_15_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_18_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_18_15_7  (
            .in0(_gnd_net_),
            .in1(N__45377),
            .in2(N__45958),
            .in3(N__45344),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__47278),
            .ce(N__45726),
            .sr(N__46632));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_18_16_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_18_16_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_18_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_18_16_0  (
            .in0(_gnd_net_),
            .in1(N__45341),
            .in2(N__45898),
            .in3(N__45305),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ),
            .ltout(),
            .carryin(bfn_18_16_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__47266),
            .ce(N__45731),
            .sr(N__46637));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_18_16_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_18_16_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_18_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_18_16_1  (
            .in0(_gnd_net_),
            .in1(N__45962),
            .in2(N__45844),
            .in3(N__45920),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__47266),
            .ce(N__45731),
            .sr(N__46637));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_18_16_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_18_16_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_18_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_18_16_2  (
            .in0(_gnd_net_),
            .in1(N__45917),
            .in2(N__45899),
            .in3(N__45863),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__47266),
            .ce(N__45731),
            .sr(N__46637));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_18_16_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_18_16_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_18_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_18_16_3  (
            .in0(_gnd_net_),
            .in1(N__45860),
            .in2(N__45845),
            .in3(N__45809),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__47266),
            .ce(N__45731),
            .sr(N__46637));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_18_16_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_18_16_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_18_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_18_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45806),
            .lcout(\delay_measurement_inst.elapsed_time_tr_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47266),
            .ce(N__45731),
            .sr(N__46637));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_18_17_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_18_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_18_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_18_17_0  (
            .in0(_gnd_net_),
            .in1(N__45674),
            .in2(N__45668),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_17_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_18_17_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_18_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_18_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_18_17_1  (
            .in0(_gnd_net_),
            .in1(N__45644),
            .in2(_gnd_net_),
            .in3(N__45626),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_18_17_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_18_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_18_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_18_17_2  (
            .in0(_gnd_net_),
            .in1(N__45623),
            .in2(N__45614),
            .in3(N__45593),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_18_17_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_18_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_18_17_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_18_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__46115),
            .in3(N__46094),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_18_17_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_18_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_18_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_18_17_4  (
            .in0(_gnd_net_),
            .in1(N__46091),
            .in2(_gnd_net_),
            .in3(N__46073),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_18_17_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_18_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_18_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_18_17_5  (
            .in0(_gnd_net_),
            .in1(N__46070),
            .in2(_gnd_net_),
            .in3(N__46052),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_18_17_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_18_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_18_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_18_17_6  (
            .in0(_gnd_net_),
            .in1(N__46049),
            .in2(_gnd_net_),
            .in3(N__46031),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_18_17_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_18_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_18_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_18_17_7  (
            .in0(_gnd_net_),
            .in1(N__46028),
            .in2(_gnd_net_),
            .in3(N__46010),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_18_18_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_18_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_18_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_18_18_0  (
            .in0(_gnd_net_),
            .in1(N__48215),
            .in2(_gnd_net_),
            .in3(N__46007),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9 ),
            .ltout(),
            .carryin(bfn_18_18_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_18_18_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_18_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_18_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_18_18_1  (
            .in0(_gnd_net_),
            .in1(N__46004),
            .in2(_gnd_net_),
            .in3(N__45986),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_18_18_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_18_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_18_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_18_18_2  (
            .in0(_gnd_net_),
            .in1(N__45983),
            .in2(_gnd_net_),
            .in3(N__45965),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_18_18_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_18_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_18_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_18_18_3  (
            .in0(_gnd_net_),
            .in1(N__46292),
            .in2(_gnd_net_),
            .in3(N__46274),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_18_18_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_18_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_18_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_18_18_4  (
            .in0(_gnd_net_),
            .in1(N__46271),
            .in2(_gnd_net_),
            .in3(N__46253),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_18_18_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_18_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_18_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_18_18_5  (
            .in0(_gnd_net_),
            .in1(N__46250),
            .in2(_gnd_net_),
            .in3(N__46232),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_18_18_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_18_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_18_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_18_18_6  (
            .in0(_gnd_net_),
            .in1(N__46229),
            .in2(_gnd_net_),
            .in3(N__46205),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_18_18_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_18_18_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_18_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_18_18_7  (
            .in0(_gnd_net_),
            .in1(N__46201),
            .in2(_gnd_net_),
            .in3(N__46181),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_18_19_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_18_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_18_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_18_19_0  (
            .in0(_gnd_net_),
            .in1(N__46178),
            .in2(_gnd_net_),
            .in3(N__46160),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17 ),
            .ltout(),
            .carryin(bfn_18_19_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_18_19_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_18_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_18_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_18_19_1  (
            .in0(_gnd_net_),
            .in1(N__46157),
            .in2(_gnd_net_),
            .in3(N__46139),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_18_19_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_18_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_18_19_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_18_19_2  (
            .in0(_gnd_net_),
            .in1(N__46136),
            .in2(_gnd_net_),
            .in3(N__46124),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_18_20_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_18_20_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_18_20_2 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_18_20_2  (
            .in0(N__47915),
            .in1(N__48184),
            .in2(N__48074),
            .in3(N__48224),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47234),
            .ce(),
            .sr(N__46669));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_18_20_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_18_20_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_18_20_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_18_20_3  (
            .in0(N__48183),
            .in1(N__48067),
            .in2(_gnd_net_),
            .in3(N__47914),
            .lcout(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_0_13_LC_18_20_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_0_13_LC_18_20_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_0_13_LC_18_20_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_0_13_LC_18_20_4  (
            .in0(_gnd_net_),
            .in1(N__47530),
            .in2(_gnd_net_),
            .in3(N__47684),
            .lcout(\phase_controller_inst1.stoper_tr.N_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_14_LC_18_20_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_14_LC_18_20_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_14_LC_18_20_7 .LUT_INIT=16'b1110111011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_14_LC_18_20_7  (
            .in0(N__47810),
            .in1(N__47779),
            .in2(N__47694),
            .in3(N__47735),
            .lcout(measured_delay_tr_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47234),
            .ce(),
            .sr(N__46669));
    defparam \phase_controller_slave.start_timer_hc_RNO_0_LC_18_21_3 .C_ON=1'b0;
    defparam \phase_controller_slave.start_timer_hc_RNO_0_LC_18_21_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_slave.start_timer_hc_RNO_0_LC_18_21_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_slave.start_timer_hc_RNO_0_LC_18_21_3  (
            .in0(_gnd_net_),
            .in1(N__47666),
            .in2(_gnd_net_),
            .in3(N__47642),
            .lcout(\phase_controller_slave.N_211 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_20_20_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_20_20_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_20_20_1 .LUT_INIT=16'b1111010011110101;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_9_LC_20_20_1  (
            .in0(N__47604),
            .in1(N__47540),
            .in2(N__47447),
            .in3(N__47402),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47250),
            .ce(N__46826),
            .sr(N__46670));
endmodule // MAIN
